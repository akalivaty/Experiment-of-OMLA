

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U548 ( .A1(G2105), .A2(G2104), .ZN(n871) );
  INV_X1 U549 ( .A(KEYINPUT105), .ZN(n756) );
  NOR2_X1 U550 ( .A1(n805), .A2(n804), .ZN(n807) );
  AND2_X1 U551 ( .A1(n770), .A2(n769), .ZN(n805) );
  XNOR2_X1 U552 ( .A(n757), .B(n756), .ZN(n758) );
  AND2_X1 U553 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U554 ( .A1(n690), .A2(n689), .ZN(n692) );
  BUF_X1 U555 ( .A(n548), .Z(n533) );
  NOR2_X4 U556 ( .A1(n557), .A2(n556), .ZN(G160) );
  XNOR2_X2 U557 ( .A(KEYINPUT66), .B(n553), .ZN(n557) );
  XNOR2_X1 U558 ( .A(n718), .B(KEYINPUT29), .ZN(n719) );
  XNOR2_X1 U559 ( .A(KEYINPUT31), .B(KEYINPUT103), .ZN(n691) );
  NOR2_X1 U560 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  NOR2_X2 U561 ( .A1(n711), .A2(n710), .ZN(n714) );
  XNOR2_X2 U562 ( .A(n532), .B(KEYINPUT64), .ZN(n548) );
  AND2_X2 U563 ( .A1(G2104), .A2(n531), .ZN(n532) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n527), .Z(n543) );
  INV_X1 U565 ( .A(KEYINPUT102), .ZN(n718) );
  XNOR2_X1 U566 ( .A(n720), .B(n719), .ZN(n723) );
  XNOR2_X1 U567 ( .A(n692), .B(n691), .ZN(n725) );
  INV_X1 U568 ( .A(n707), .ZN(n727) );
  NOR2_X2 U569 ( .A1(G2104), .A2(n524), .ZN(n872) );
  XOR2_X1 U570 ( .A(KEYINPUT77), .B(n591), .Z(n985) );
  NOR2_X1 U571 ( .A1(n523), .A2(n522), .ZN(G171) );
  INV_X1 U572 ( .A(G651), .ZN(n516) );
  NOR2_X1 U573 ( .A1(n516), .A2(G543), .ZN(n512) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n512), .Z(n584) );
  BUF_X1 U575 ( .A(n584), .Z(n642) );
  NAND2_X1 U576 ( .A1(n642), .A2(G64), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT68), .ZN(n515) );
  XOR2_X1 U578 ( .A(G543), .B(KEYINPUT0), .Z(n626) );
  NOR2_X2 U579 ( .A1(G651), .A2(n626), .ZN(n646) );
  NAND2_X1 U580 ( .A1(G52), .A2(n646), .ZN(n514) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n523) );
  NOR2_X2 U582 ( .A1(n626), .A2(n516), .ZN(n640) );
  NAND2_X1 U583 ( .A1(n640), .A2(G77), .ZN(n517) );
  XOR2_X1 U584 ( .A(KEYINPUT69), .B(n517), .Z(n519) );
  NOR2_X2 U585 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U586 ( .A1(n643), .A2(G90), .ZN(n518) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT70), .B(n520), .Z(n521) );
  XNOR2_X1 U589 ( .A(KEYINPUT9), .B(n521), .ZN(n522) );
  AND2_X1 U590 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U591 ( .A(G2105), .ZN(n524) );
  NAND2_X1 U592 ( .A1(G123), .A2(n872), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n525), .B(KEYINPUT18), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n526), .B(KEYINPUT80), .ZN(n529) );
  NAND2_X1 U595 ( .A1(G135), .A2(n543), .ZN(n528) );
  NAND2_X1 U596 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT81), .B(n530), .ZN(n537) );
  INV_X1 U598 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U599 ( .A1(n533), .A2(G99), .ZN(n535) );
  NAND2_X1 U600 ( .A1(G111), .A2(n871), .ZN(n534) );
  AND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U602 ( .A1(n537), .A2(n536), .ZN(n925) );
  XNOR2_X1 U603 ( .A(G2096), .B(n925), .ZN(n538) );
  OR2_X1 U604 ( .A1(G2100), .A2(n538), .ZN(G156) );
  INV_X1 U605 ( .A(G120), .ZN(G236) );
  INV_X1 U606 ( .A(G69), .ZN(G235) );
  INV_X1 U607 ( .A(G108), .ZN(G238) );
  INV_X1 U608 ( .A(G132), .ZN(G219) );
  NAND2_X1 U609 ( .A1(n871), .A2(G114), .ZN(n539) );
  XOR2_X1 U610 ( .A(KEYINPUT93), .B(n539), .Z(n541) );
  NAND2_X1 U611 ( .A1(n872), .A2(G126), .ZN(n540) );
  NAND2_X1 U612 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(n542), .B(KEYINPUT94), .ZN(n547) );
  NAND2_X1 U614 ( .A1(G138), .A2(n543), .ZN(n545) );
  NAND2_X1 U615 ( .A1(G102), .A2(n548), .ZN(n544) );
  NAND2_X1 U616 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U617 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U618 ( .A1(n548), .A2(G101), .ZN(n549) );
  XNOR2_X1 U619 ( .A(n549), .B(KEYINPUT23), .ZN(n550) );
  XNOR2_X1 U620 ( .A(n550), .B(KEYINPUT65), .ZN(n552) );
  NAND2_X1 U621 ( .A1(G125), .A2(n872), .ZN(n551) );
  NAND2_X1 U622 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U623 ( .A1(G113), .A2(n871), .ZN(n555) );
  NAND2_X1 U624 ( .A1(G137), .A2(n543), .ZN(n554) );
  NAND2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U626 ( .A1(G89), .A2(n643), .ZN(n558) );
  XOR2_X1 U627 ( .A(KEYINPUT79), .B(n558), .Z(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G76), .A2(n640), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G63), .A2(n642), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G51), .A2(n646), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U640 ( .A(n569), .B(KEYINPUT10), .Z(n912) );
  NAND2_X1 U641 ( .A1(n912), .A2(G567), .ZN(n570) );
  XOR2_X1 U642 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U643 ( .A1(n642), .A2(G56), .ZN(n571) );
  XOR2_X1 U644 ( .A(KEYINPUT14), .B(n571), .Z(n579) );
  NAND2_X1 U645 ( .A1(G68), .A2(n640), .ZN(n575) );
  XOR2_X1 U646 ( .A(KEYINPUT73), .B(KEYINPUT12), .Z(n573) );
  NAND2_X1 U647 ( .A1(G81), .A2(n643), .ZN(n572) );
  XNOR2_X1 U648 ( .A(n573), .B(n572), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U650 ( .A(n576), .B(KEYINPUT74), .ZN(n577) );
  XOR2_X1 U651 ( .A(KEYINPUT13), .B(n577), .Z(n578) );
  NOR2_X1 U652 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n646), .A2(G43), .ZN(n580) );
  NAND2_X1 U654 ( .A1(n581), .A2(n580), .ZN(n995) );
  INV_X1 U655 ( .A(G860), .ZN(n610) );
  OR2_X1 U656 ( .A1(n995), .A2(n610), .ZN(G153) );
  XNOR2_X1 U657 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U658 ( .A1(G79), .A2(n640), .ZN(n583) );
  NAND2_X1 U659 ( .A1(G92), .A2(n643), .ZN(n582) );
  AND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n584), .A2(G66), .ZN(n585) );
  XOR2_X1 U662 ( .A(KEYINPUT76), .B(n585), .Z(n587) );
  AND2_X1 U663 ( .A1(G54), .A2(n646), .ZN(n586) );
  NOR2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n590), .B(KEYINPUT15), .ZN(n591) );
  INV_X1 U667 ( .A(n985), .ZN(n704) );
  INV_X1 U668 ( .A(G868), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n704), .A2(n601), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT78), .ZN(n594) );
  NAND2_X1 U671 ( .A1(G868), .A2(G301), .ZN(n593) );
  NAND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U673 ( .A1(G65), .A2(n642), .ZN(n596) );
  NAND2_X1 U674 ( .A1(G53), .A2(n646), .ZN(n595) );
  NAND2_X1 U675 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G78), .A2(n640), .ZN(n598) );
  NAND2_X1 U677 ( .A1(G91), .A2(n643), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n989) );
  XNOR2_X1 U680 ( .A(n989), .B(KEYINPUT71), .ZN(G299) );
  NAND2_X1 U681 ( .A1(G286), .A2(G868), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G299), .A2(n601), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U684 ( .A1(n610), .A2(G559), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n604), .A2(n985), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U687 ( .A1(G868), .A2(n995), .ZN(n608) );
  NAND2_X1 U688 ( .A1(G868), .A2(n985), .ZN(n606) );
  NOR2_X1 U689 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U690 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G559), .A2(n985), .ZN(n609) );
  XOR2_X1 U692 ( .A(n995), .B(n609), .Z(n660) );
  NAND2_X1 U693 ( .A1(n610), .A2(n660), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G80), .A2(n640), .ZN(n612) );
  NAND2_X1 U695 ( .A1(G67), .A2(n642), .ZN(n611) );
  NAND2_X1 U696 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U697 ( .A1(G93), .A2(n643), .ZN(n614) );
  NAND2_X1 U698 ( .A1(G55), .A2(n646), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n662) );
  XOR2_X1 U701 ( .A(n617), .B(n662), .Z(G145) );
  NAND2_X1 U702 ( .A1(G75), .A2(n640), .ZN(n619) );
  NAND2_X1 U703 ( .A1(G88), .A2(n643), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U705 ( .A(KEYINPUT84), .B(n620), .ZN(n624) );
  NAND2_X1 U706 ( .A1(G62), .A2(n642), .ZN(n622) );
  NAND2_X1 U707 ( .A1(G50), .A2(n646), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U709 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(n625), .ZN(G303) );
  NAND2_X1 U711 ( .A1(G87), .A2(n626), .ZN(n627) );
  XNOR2_X1 U712 ( .A(n627), .B(KEYINPUT82), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G49), .A2(n646), .ZN(n629) );
  NAND2_X1 U714 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U715 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U716 ( .A1(n642), .A2(n630), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(G288) );
  NAND2_X1 U718 ( .A1(G60), .A2(n642), .ZN(n634) );
  NAND2_X1 U719 ( .A1(G47), .A2(n646), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G72), .A2(n640), .ZN(n635) );
  XNOR2_X1 U722 ( .A(KEYINPUT67), .B(n635), .ZN(n636) );
  NOR2_X1 U723 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n643), .A2(G85), .ZN(n638) );
  NAND2_X1 U725 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U726 ( .A1(G73), .A2(n640), .ZN(n641) );
  XNOR2_X1 U727 ( .A(n641), .B(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G61), .A2(n642), .ZN(n645) );
  NAND2_X1 U729 ( .A1(G86), .A2(n643), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U731 ( .A1(G48), .A2(n646), .ZN(n647) );
  XNOR2_X1 U732 ( .A(KEYINPUT83), .B(n647), .ZN(n648) );
  NOR2_X1 U733 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G305) );
  XNOR2_X1 U735 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n653) );
  XNOR2_X1 U736 ( .A(G288), .B(KEYINPUT19), .ZN(n652) );
  XNOR2_X1 U737 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U738 ( .A(KEYINPUT88), .B(n654), .ZN(n656) );
  XNOR2_X1 U739 ( .A(G290), .B(n662), .ZN(n655) );
  XNOR2_X1 U740 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U741 ( .A(n657), .B(G305), .Z(n658) );
  XNOR2_X1 U742 ( .A(G299), .B(n658), .ZN(n659) );
  XOR2_X1 U743 ( .A(G303), .B(n659), .Z(n891) );
  XNOR2_X1 U744 ( .A(n660), .B(n891), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n661), .A2(G868), .ZN(n664) );
  OR2_X1 U746 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n668), .A2(G2072), .ZN(n669) );
  XOR2_X1 U753 ( .A(KEYINPUT89), .B(n669), .Z(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U755 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U757 ( .A(KEYINPUT90), .B(n670), .Z(n671) );
  XNOR2_X1 U758 ( .A(n671), .B(KEYINPUT22), .ZN(n672) );
  NOR2_X1 U759 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G96), .A2(n673), .ZN(n828) );
  NAND2_X1 U761 ( .A1(n828), .A2(G2106), .ZN(n679) );
  NOR2_X1 U762 ( .A1(G235), .A2(G236), .ZN(n674) );
  XNOR2_X1 U763 ( .A(n674), .B(KEYINPUT91), .ZN(n675) );
  NOR2_X1 U764 ( .A1(G238), .A2(n675), .ZN(n676) );
  NAND2_X1 U765 ( .A1(G57), .A2(n676), .ZN(n827) );
  NAND2_X1 U766 ( .A1(G567), .A2(n827), .ZN(n677) );
  XNOR2_X1 U767 ( .A(KEYINPUT92), .B(n677), .ZN(n678) );
  NAND2_X1 U768 ( .A1(n679), .A2(n678), .ZN(n829) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n680) );
  NOR2_X1 U770 ( .A1(n829), .A2(n680), .ZN(n824) );
  NAND2_X1 U771 ( .A1(n824), .A2(G36), .ZN(G176) );
  NOR2_X1 U772 ( .A1(G164), .A2(G1384), .ZN(n791) );
  AND2_X1 U773 ( .A1(n791), .A2(G40), .ZN(n682) );
  AND2_X2 U774 ( .A1(G160), .A2(n682), .ZN(n707) );
  NAND2_X1 U775 ( .A1(G8), .A2(n727), .ZN(n726) );
  NOR2_X1 U776 ( .A1(G1966), .A2(n726), .ZN(n739) );
  NOR2_X1 U777 ( .A1(G2084), .A2(n727), .ZN(n736) );
  NOR2_X1 U778 ( .A1(n739), .A2(n736), .ZN(n683) );
  NAND2_X1 U779 ( .A1(n683), .A2(G8), .ZN(n684) );
  XNOR2_X1 U780 ( .A(KEYINPUT30), .B(n684), .ZN(n685) );
  NOR2_X1 U781 ( .A1(G168), .A2(n685), .ZN(n690) );
  INV_X1 U782 ( .A(n707), .ZN(n693) );
  NOR2_X1 U783 ( .A1(n709), .A2(G1961), .ZN(n686) );
  XNOR2_X1 U784 ( .A(n686), .B(KEYINPUT101), .ZN(n688) );
  XNOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .ZN(n943) );
  NAND2_X1 U786 ( .A1(n707), .A2(n943), .ZN(n687) );
  NAND2_X1 U787 ( .A1(n688), .A2(n687), .ZN(n721) );
  NOR2_X1 U788 ( .A1(G171), .A2(n721), .ZN(n689) );
  INV_X1 U789 ( .A(n693), .ZN(n709) );
  NAND2_X1 U790 ( .A1(n709), .A2(G2067), .ZN(n695) );
  NAND2_X1 U791 ( .A1(G1348), .A2(n727), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n695), .A2(n694), .ZN(n703) );
  NOR2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n702) );
  AND2_X1 U794 ( .A1(n707), .A2(G1996), .ZN(n696) );
  XNOR2_X1 U795 ( .A(n696), .B(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U796 ( .A1(n727), .A2(G1341), .ZN(n698) );
  INV_X1 U797 ( .A(n995), .ZN(n697) );
  NAND2_X1 U798 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U799 ( .A1(n700), .A2(n699), .ZN(n701) );
  OR2_X1 U800 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n707), .A2(G2072), .ZN(n708) );
  XNOR2_X1 U804 ( .A(n708), .B(KEYINPUT27), .ZN(n711) );
  INV_X1 U805 ( .A(G1956), .ZN(n988) );
  NOR2_X1 U806 ( .A1(n988), .A2(n709), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n714), .A2(n989), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U809 ( .A1(n714), .A2(n989), .ZN(n715) );
  XOR2_X1 U810 ( .A(n715), .B(KEYINPUT28), .Z(n716) );
  NAND2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U812 ( .A1(G171), .A2(n721), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n738) );
  NAND2_X1 U815 ( .A1(n738), .A2(G286), .ZN(n734) );
  INV_X1 U816 ( .A(G8), .ZN(n732) );
  BUF_X1 U817 ( .A(n726), .Z(n766) );
  NOR2_X1 U818 ( .A1(G1971), .A2(n766), .ZN(n729) );
  NOR2_X1 U819 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U820 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U822 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U823 ( .A(n735), .B(KEYINPUT32), .Z(n742) );
  NAND2_X1 U824 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n740) );
  NOR2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U828 ( .A(KEYINPUT104), .B(n743), .Z(n761) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n745) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n1006) );
  INV_X1 U832 ( .A(n766), .ZN(n750) );
  NAND2_X1 U833 ( .A1(n745), .A2(n750), .ZN(n746) );
  NAND2_X1 U834 ( .A1(n746), .A2(KEYINPUT33), .ZN(n748) );
  AND2_X1 U835 ( .A1(n1006), .A2(n748), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n761), .A2(n747), .ZN(n755) );
  INV_X1 U837 ( .A(n748), .ZN(n753) );
  INV_X1 U838 ( .A(KEYINPUT33), .ZN(n749) );
  NAND2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n990) );
  AND2_X1 U840 ( .A1(n749), .A2(n990), .ZN(n751) );
  AND2_X1 U841 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U842 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n757) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n1000) );
  NAND2_X1 U845 ( .A1(n758), .A2(n1000), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT106), .ZN(n770) );
  NOR2_X1 U847 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U848 ( .A1(G8), .A2(n760), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n763) );
  AND2_X1 U850 ( .A1(n763), .A2(n766), .ZN(n768) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U852 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U853 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U855 ( .A1(G131), .A2(n543), .ZN(n772) );
  NAND2_X1 U856 ( .A1(G95), .A2(n533), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n778) );
  NAND2_X1 U858 ( .A1(n872), .A2(G119), .ZN(n773) );
  XNOR2_X1 U859 ( .A(n773), .B(KEYINPUT96), .ZN(n775) );
  NAND2_X1 U860 ( .A1(G107), .A2(n871), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT97), .B(n776), .Z(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U864 ( .A(KEYINPUT98), .B(n779), .Z(n866) );
  NAND2_X1 U865 ( .A1(G1991), .A2(n866), .ZN(n788) );
  NAND2_X1 U866 ( .A1(G117), .A2(n871), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G129), .A2(n872), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n784) );
  NAND2_X1 U869 ( .A1(n533), .A2(G105), .ZN(n782) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n782), .Z(n783) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n543), .A2(G141), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n786), .A2(n785), .ZN(n881) );
  NAND2_X1 U874 ( .A1(G1996), .A2(n881), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U876 ( .A(KEYINPUT99), .B(n789), .ZN(n934) );
  NAND2_X1 U877 ( .A1(G160), .A2(G40), .ZN(n790) );
  NOR2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n818) );
  INV_X1 U879 ( .A(n818), .ZN(n792) );
  NOR2_X1 U880 ( .A1(n934), .A2(n792), .ZN(n811) );
  XOR2_X1 U881 ( .A(KEYINPUT100), .B(n811), .Z(n803) );
  XNOR2_X1 U882 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  NAND2_X1 U883 ( .A1(G104), .A2(n533), .ZN(n793) );
  XOR2_X1 U884 ( .A(KEYINPUT95), .B(n793), .Z(n795) );
  NAND2_X1 U885 ( .A1(n543), .A2(G140), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U887 ( .A(KEYINPUT34), .B(n796), .ZN(n801) );
  NAND2_X1 U888 ( .A1(G116), .A2(n871), .ZN(n798) );
  NAND2_X1 U889 ( .A1(G128), .A2(n872), .ZN(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT35), .B(n799), .Z(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U893 ( .A(KEYINPUT36), .B(n802), .ZN(n888) );
  NOR2_X1 U894 ( .A1(n816), .A2(n888), .ZN(n924) );
  NAND2_X1 U895 ( .A1(n818), .A2(n924), .ZN(n814) );
  NAND2_X1 U896 ( .A1(n803), .A2(n814), .ZN(n804) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n997) );
  NAND2_X1 U898 ( .A1(n997), .A2(n818), .ZN(n806) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n821) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n881), .ZN(n808) );
  XOR2_X1 U901 ( .A(KEYINPUT107), .B(n808), .Z(n920) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n866), .ZN(n928) );
  NOR2_X1 U904 ( .A1(n809), .A2(n928), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n920), .A2(n812), .ZN(n813) );
  XNOR2_X1 U907 ( .A(KEYINPUT39), .B(n813), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n816), .A2(n888), .ZN(n917) );
  NAND2_X1 U910 ( .A1(n817), .A2(n917), .ZN(n819) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U912 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U913 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U914 ( .A1(G2106), .A2(n912), .ZN(G217) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G1), .A2(G3), .ZN(n825) );
  NAND2_X1 U918 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(KEYINPUT108), .ZN(G188) );
  XNOR2_X1 U920 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  NOR2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U923 ( .A(G325), .ZN(G261) );
  INV_X1 U924 ( .A(n829), .ZN(G319) );
  XOR2_X1 U925 ( .A(G2100), .B(G2096), .Z(n831) );
  XNOR2_X1 U926 ( .A(KEYINPUT42), .B(G2678), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n835) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(G2072), .Z(n833) );
  XNOR2_X1 U929 ( .A(G2067), .B(G2090), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U931 ( .A(n835), .B(n834), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2084), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(G227) );
  XNOR2_X1 U934 ( .A(KEYINPUT111), .B(n988), .ZN(n839) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U937 ( .A(n840), .B(KEYINPUT41), .Z(n842) );
  XNOR2_X1 U938 ( .A(G1966), .B(G1961), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U940 ( .A(G1976), .B(G1981), .Z(n844) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1971), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U943 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U944 ( .A(KEYINPUT110), .B(G2474), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(G229) );
  NAND2_X1 U946 ( .A1(n872), .A2(G124), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n849), .B(KEYINPUT44), .ZN(n851) );
  NAND2_X1 U948 ( .A1(G100), .A2(n533), .ZN(n850) );
  NAND2_X1 U949 ( .A1(n851), .A2(n850), .ZN(n855) );
  NAND2_X1 U950 ( .A1(G112), .A2(n871), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G136), .A2(n543), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n854) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(G162) );
  NAND2_X1 U954 ( .A1(n543), .A2(G142), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n856), .B(KEYINPUT114), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G106), .A2(n533), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n859), .B(KEYINPUT45), .ZN(n865) );
  NAND2_X1 U959 ( .A1(n872), .A2(G130), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n860), .B(KEYINPUT112), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G118), .A2(n871), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  XNOR2_X1 U963 ( .A(KEYINPUT113), .B(n863), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n925), .B(n868), .ZN(n880) );
  NAND2_X1 U967 ( .A1(G139), .A2(n543), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G103), .A2(n533), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G115), .A2(n871), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G127), .A2(n872), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U974 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U975 ( .A(KEYINPUT115), .B(n878), .Z(n913) );
  XNOR2_X1 U976 ( .A(G160), .B(n913), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n880), .B(n879), .ZN(n885) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n881), .B(KEYINPUT116), .ZN(n882) );
  XNOR2_X1 U980 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U981 ( .A(n885), .B(n884), .Z(n887) );
  XNOR2_X1 U982 ( .A(G164), .B(G162), .ZN(n886) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n889) );
  XOR2_X1 U984 ( .A(n889), .B(n888), .Z(n890) );
  NOR2_X1 U985 ( .A1(G37), .A2(n890), .ZN(G395) );
  XNOR2_X1 U986 ( .A(n891), .B(n995), .ZN(n892) );
  XOR2_X1 U987 ( .A(n892), .B(n985), .Z(n894) );
  XOR2_X1 U988 ( .A(G286), .B(G171), .Z(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(n896) );
  XOR2_X1 U991 ( .A(KEYINPUT117), .B(n896), .Z(G397) );
  XOR2_X1 U992 ( .A(G2451), .B(G2430), .Z(n898) );
  XNOR2_X1 U993 ( .A(G2438), .B(G2443), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n904) );
  XOR2_X1 U995 ( .A(G2435), .B(G2454), .Z(n900) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n899) );
  XNOR2_X1 U997 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U998 ( .A(G2446), .B(G2427), .Z(n901) );
  XNOR2_X1 U999 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U1000 ( .A(n904), .B(n903), .Z(n905) );
  NAND2_X1 U1001 ( .A1(G14), .A2(n905), .ZN(n911) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n911), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G303), .ZN(G166) );
  INV_X1 U1010 ( .A(G57), .ZN(G237) );
  INV_X1 U1011 ( .A(n911), .ZN(G401) );
  INV_X1 U1012 ( .A(n912), .ZN(G223) );
  INV_X1 U1013 ( .A(KEYINPUT55), .ZN(n959) );
  XOR2_X1 U1014 ( .A(G2072), .B(n913), .Z(n915) );
  XOR2_X1 U1015 ( .A(G164), .B(G2078), .Z(n914) );
  NOR2_X1 U1016 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1017 ( .A(n916), .B(KEYINPUT50), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n932) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n921), .Z(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT118), .B(n922), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n930) );
  XNOR2_X1 U1024 ( .A(G160), .B(G2084), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1030 ( .A(KEYINPUT52), .B(n935), .Z(n936) );
  NAND2_X1 U1031 ( .A1(n959), .A2(n936), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(G29), .ZN(n1020) );
  XOR2_X1 U1033 ( .A(KEYINPUT120), .B(G34), .Z(n939) );
  XNOR2_X1 U1034 ( .A(G2084), .B(KEYINPUT54), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(n939), .B(n938), .ZN(n955) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n953) );
  XNOR2_X1 U1037 ( .A(G2067), .B(G26), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G32), .B(G1996), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n948) );
  XOR2_X1 U1040 ( .A(G2072), .B(G33), .Z(n942) );
  NAND2_X1 U1041 ( .A1(n942), .A2(G28), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G27), .B(n943), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n944), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1046 ( .A(G25), .B(G1991), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n958) );
  NOR2_X1 U1051 ( .A1(G29), .A2(KEYINPUT55), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n956), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n957), .ZN(n1018) );
  OR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n1016) );
  XOR2_X1 U1055 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n982) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G21), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G1961), .B(G5), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n980) );
  XOR2_X1 U1059 ( .A(G1971), .B(G22), .Z(n962) );
  XNOR2_X1 U1060 ( .A(KEYINPUT124), .B(n962), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G1986), .B(G24), .ZN(n964) );
  XNOR2_X1 U1062 ( .A(G23), .B(G1976), .ZN(n963) );
  NOR2_X1 U1063 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1065 ( .A(n967), .B(KEYINPUT58), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(KEYINPUT59), .B(G1348), .ZN(n968) );
  XNOR2_X1 U1067 ( .A(n968), .B(G4), .ZN(n974) );
  XOR2_X1 U1068 ( .A(G1341), .B(G19), .Z(n970) );
  XOR2_X1 U1069 ( .A(G1956), .B(G20), .Z(n969) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1071 ( .A(G6), .B(G1981), .ZN(n971) );
  NOR2_X1 U1072 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1073 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1074 ( .A(n975), .B(KEYINPUT60), .Z(n976) );
  XNOR2_X1 U1075 ( .A(KEYINPUT123), .B(n976), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1077 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1078 ( .A(n982), .B(n981), .ZN(n983) );
  XNOR2_X1 U1079 ( .A(n983), .B(KEYINPUT61), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(G16), .A2(n984), .ZN(n1013) );
  XOR2_X1 U1081 ( .A(G16), .B(KEYINPUT56), .Z(n1011) );
  NAND2_X1 U1082 ( .A1(G1971), .A2(G303), .ZN(n987) );
  XNOR2_X1 U1083 ( .A(G1348), .B(n985), .ZN(n986) );
  NAND2_X1 U1084 ( .A1(n987), .A2(n986), .ZN(n1008) );
  XOR2_X1 U1085 ( .A(n989), .B(n988), .Z(n991) );
  NAND2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(G1961), .B(G171), .ZN(n992) );
  XNOR2_X1 U1088 ( .A(KEYINPUT121), .B(n992), .ZN(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(G1341), .B(n995), .ZN(n996) );
  NOR2_X1 U1091 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G1966), .B(G168), .ZN(n1001) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1095 ( .A(KEYINPUT57), .B(n1002), .Z(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(KEYINPUT122), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT127), .B(n1014), .Z(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1021), .ZN(G150) );
  INV_X1 U1107 ( .A(G150), .ZN(G311) );
endmodule

