//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT75), .B(G902), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n194));
  INV_X1    g008(.A(G107), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n194), .A2(new_n195), .A3(G104), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n192), .A2(G107), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n193), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G101), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT81), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n193), .A2(new_n196), .A3(new_n201), .A4(new_n197), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n202), .A2(KEYINPUT4), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT81), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n198), .A2(new_n204), .A3(G101), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT0), .A2(G128), .ZN(new_n212));
  OR2_X1    g026(.A1(KEYINPUT0), .A2(G128), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n215), .B1(new_n209), .B2(G146), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(KEYINPUT64), .A3(G143), .ZN(new_n217));
  INV_X1    g031(.A(new_n212), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n216), .A2(new_n217), .A3(new_n210), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT4), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n198), .A2(new_n222), .A3(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n206), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(KEYINPUT67), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  OR2_X1    g047(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n228), .B1(new_n234), .B2(new_n229), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n226), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n231), .A2(G137), .ZN(new_n237));
  INV_X1    g051(.A(new_n229), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n226), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n240), .A2(new_n232), .A3(new_n230), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n216), .A2(new_n217), .A3(new_n210), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT1), .B1(new_n209), .B2(G146), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(KEYINPUT1), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n216), .A2(new_n217), .A3(new_n250), .A4(new_n210), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n192), .A2(G107), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n195), .A2(G104), .ZN(new_n254));
  OAI21_X1  g068(.A(G101), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n202), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT10), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n249), .A2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G128), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n263), .A2(new_n246), .B1(new_n208), .B2(new_n210), .ZN(new_n264));
  AND4_X1   g078(.A1(new_n216), .A2(new_n217), .A3(new_n250), .A4(new_n210), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT71), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT69), .B(G128), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(G143), .B2(new_n207), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n211), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n251), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n266), .A2(KEYINPUT10), .A3(new_n272), .A4(new_n256), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n224), .A2(new_n244), .A3(new_n259), .A4(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  INV_X1    g089(.A(G953), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(G227), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n275), .B(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n202), .A2(new_n255), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(new_n251), .A3(new_n270), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n251), .B2(new_n248), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT12), .B(new_n243), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT82), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n243), .B1(new_n284), .B2(new_n285), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n257), .A2(new_n283), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n292), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n243), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n281), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n259), .A2(new_n273), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n244), .B1(new_n296), .B2(new_n224), .ZN(new_n297));
  INV_X1    g111(.A(new_n274), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n278), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI211_X1 g113(.A(G469), .B(new_n191), .C1(new_n295), .C2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n279), .B1(new_n294), .B2(new_n274), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n297), .A2(new_n280), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G469), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT83), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n224), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n243), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n281), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT12), .B1(new_n292), .B2(new_n243), .ZN(new_n312));
  AOI221_X4 g126(.A(new_n290), .B1(new_n242), .B2(new_n236), .C1(new_n257), .C2(new_n283), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n312), .B1(KEYINPUT82), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n298), .B1(new_n314), .B2(new_n288), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(new_n279), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n308), .B1(new_n316), .B2(new_n301), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT83), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n189), .B1(new_n307), .B2(new_n318), .ZN(new_n319));
  AOI211_X1 g133(.A(new_n276), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT21), .B(G898), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G952), .ZN(new_n323));
  AOI211_X1 g137(.A(G953), .B(new_n323), .C1(G234), .C2(G237), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G122), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G119), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G116), .ZN(new_n331));
  INV_X1    g145(.A(G116), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G119), .ZN(new_n333));
  INV_X1    g147(.A(G113), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(KEYINPUT2), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n333), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n333), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT2), .B(G113), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n341), .A2(new_n223), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n206), .A2(new_n342), .A3(KEYINPUT84), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT5), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n344), .B(G113), .C1(KEYINPUT5), .C2(new_n331), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n256), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(KEYINPUT84), .B1(new_n206), .B2(new_n342), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n329), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n206), .A2(new_n342), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT84), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n352), .A2(new_n328), .A3(new_n346), .A4(new_n343), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n353), .A3(KEYINPUT6), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n220), .A2(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n270), .A2(new_n251), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(G125), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G224), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G953), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n357), .B(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n361), .B(new_n329), .C1(new_n347), .C2(new_n348), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT7), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n357), .B1(new_n364), .B2(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n345), .A2(new_n337), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n282), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n367), .A2(new_n346), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n328), .B(KEYINPUT8), .Z(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n357), .A2(new_n364), .A3(new_n359), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(G902), .B1(new_n372), .B2(new_n353), .ZN(new_n373));
  OAI21_X1  g187(.A(G210), .B1(G237), .B2(G902), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n363), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n363), .B2(new_n373), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n326), .B(new_n327), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  OR2_X1    g191(.A1(KEYINPUT73), .A2(G237), .ZN(new_n378));
  NAND2_X1  g192(.A1(KEYINPUT73), .A2(G237), .ZN(new_n379));
  AOI21_X1  g193(.A(G953), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n381));
  INV_X1    g195(.A(new_n379), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT73), .A2(G237), .ZN(new_n383));
  OAI211_X1 g197(.A(G214), .B(new_n276), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n209), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G131), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n385), .A3(new_n225), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G140), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G125), .ZN(new_n391));
  INV_X1    g205(.A(G125), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G140), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT19), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G125), .B(G140), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(KEYINPUT19), .ZN(new_n398));
  AOI21_X1  g212(.A(G146), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n399), .A2(KEYINPUT88), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n391), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n401));
  OR3_X1    g215(.A1(new_n392), .A2(KEYINPUT16), .A3(G140), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G146), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(new_n399), .B2(KEYINPUT88), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n389), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n391), .A2(new_n393), .A3(new_n207), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT86), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT87), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(KEYINPUT86), .A3(KEYINPUT87), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n410), .A2(G146), .A3(new_n394), .A4(new_n411), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n407), .A2(KEYINPUT86), .A3(KEYINPUT87), .ZN(new_n413));
  AOI21_X1  g227(.A(KEYINPUT87), .B1(new_n407), .B2(KEYINPUT86), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n413), .A2(new_n414), .B1(new_n207), .B2(new_n397), .ZN(new_n415));
  NAND2_X1  g229(.A1(KEYINPUT18), .A2(G131), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n386), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n381), .A2(new_n385), .B1(KEYINPUT18), .B2(G131), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n412), .B(new_n415), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G113), .B(G122), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(new_n192), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n406), .A2(new_n419), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(G475), .A2(G902), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n386), .B(new_n416), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n412), .A2(new_n415), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n387), .A2(new_n427), .A3(new_n388), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n401), .A2(new_n402), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n207), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n403), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n225), .B1(new_n381), .B2(new_n385), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n432), .B2(KEYINPUT17), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n425), .A2(new_n426), .B1(new_n428), .B2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n423), .B(new_n424), .C1(new_n434), .C2(new_n422), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT85), .B(KEYINPUT20), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n428), .A2(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n419), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n421), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT89), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n424), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n443), .B2(new_n424), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n423), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n332), .A2(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT91), .B(G122), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(new_n332), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G107), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n195), .B(new_n448), .C1(new_n449), .C2(new_n332), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n267), .A2(G143), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n209), .A2(G128), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT13), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT92), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(new_n209), .A3(KEYINPUT13), .A4(G128), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n454), .A2(new_n457), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G134), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n454), .A2(new_n231), .A3(new_n455), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n449), .B2(new_n332), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n450), .A2(new_n465), .A3(G107), .ZN(new_n466));
  OAI221_X1 g280(.A(new_n448), .B1(KEYINPUT14), .B2(new_n195), .C1(new_n449), .C2(new_n332), .ZN(new_n467));
  INV_X1    g281(.A(new_n463), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n231), .B1(new_n454), .B2(new_n455), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G217), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n187), .A2(new_n472), .A3(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n470), .A3(new_n473), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n190), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n477), .B2(new_n190), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT90), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n440), .B1(new_n484), .B2(new_n421), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n439), .A2(KEYINPUT90), .A3(new_n419), .A4(new_n422), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n301), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G475), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n447), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n377), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g304(.A1(new_n319), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT70), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n240), .A2(new_n225), .A3(new_n232), .A4(new_n230), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n225), .B1(new_n228), .B2(new_n232), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT68), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n264), .A2(new_n265), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT65), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n220), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n214), .A2(KEYINPUT65), .A3(new_n219), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n243), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n228), .A2(new_n232), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT68), .B1(new_n505), .B2(new_n225), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n494), .A2(new_n495), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(KEYINPUT70), .A3(new_n356), .A4(new_n493), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n341), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n266), .A2(new_n508), .A3(new_n272), .A4(new_n493), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n243), .A2(new_n221), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n340), .A3(new_n513), .A4(new_n337), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(KEYINPUT74), .A3(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n380), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n511), .B2(new_n514), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n514), .A2(new_n522), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT74), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n516), .B(new_n521), .C1(new_n523), .C2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n510), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n512), .A2(KEYINPUT30), .A3(new_n513), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT72), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n512), .A2(KEYINPUT72), .A3(new_n513), .A4(KEYINPUT30), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n529), .A2(new_n532), .A3(new_n341), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n520), .A3(new_n514), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT31), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n534), .A2(new_n537), .A3(new_n520), .A4(new_n514), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT32), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n516), .B(new_n520), .C1(new_n523), .C2(new_n526), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n521), .A3(new_n514), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT29), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n524), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n512), .A2(new_n513), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n341), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n514), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n548), .B1(new_n551), .B2(KEYINPUT28), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(KEYINPUT29), .A3(new_n520), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n190), .ZN(new_n554));
  OAI21_X1  g368(.A(G472), .B1(new_n547), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n543), .A2(new_n544), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n249), .A2(G119), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(new_n267), .B2(G119), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT24), .B(G110), .Z(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G110), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT23), .B1(new_n249), .B2(G119), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n558), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n431), .B(new_n561), .C1(new_n562), .C2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n563), .A2(new_n562), .A3(new_n565), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n559), .A2(new_n560), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n403), .B(new_n407), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n276), .A2(G221), .A3(G234), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT77), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n567), .A2(new_n570), .A3(new_n575), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n472), .B1(new_n190), .B2(G234), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT76), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G902), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT79), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n577), .A2(new_n190), .A3(new_n578), .ZN(new_n587));
  XOR2_X1   g401(.A(KEYINPUT78), .B(KEYINPUT25), .Z(new_n588));
  AOI21_X1  g402(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(KEYINPUT25), .A3(new_n190), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n586), .A3(new_n588), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI211_X1 g407(.A(new_n557), .B(new_n585), .C1(new_n593), .C2(new_n582), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n592), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n582), .B1(new_n595), .B2(new_n589), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT80), .B1(new_n596), .B2(new_n584), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n491), .A2(new_n556), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n319), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n539), .A2(KEYINPUT93), .A3(new_n190), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT93), .B1(new_n539), .B2(new_n190), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n541), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n447), .A2(new_n488), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n190), .A2(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n477), .A2(KEYINPUT33), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n475), .B2(new_n476), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n609), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n477), .A2(new_n190), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT94), .B(G478), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n377), .A2(new_n608), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n606), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT95), .ZN(new_n620));
  XOR2_X1   g434(.A(KEYINPUT34), .B(G104), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  INV_X1    g436(.A(new_n483), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n435), .B(new_n437), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(new_n624), .A3(new_n488), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n377), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n606), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  INV_X1    g443(.A(new_n541), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n602), .A2(G472), .ZN(new_n631));
  INV_X1    g445(.A(new_n604), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n576), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(new_n571), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n583), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n596), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n491), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT37), .B(G110), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G12));
  OAI21_X1  g455(.A(new_n327), .B1(new_n375), .B2(new_n376), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n324), .B1(new_n320), .B2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n625), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n556), .A2(new_n643), .A3(new_n319), .A4(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  AOI21_X1  g462(.A(new_n521), .B1(new_n534), .B2(new_n514), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n301), .B1(new_n551), .B2(new_n520), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n543), .A2(new_n544), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n637), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n375), .A2(new_n376), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT38), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n483), .B1(new_n447), .B2(new_n488), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n327), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n645), .B(KEYINPUT39), .Z(new_n659));
  NAND2_X1  g473(.A1(new_n319), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT96), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n653), .B(new_n658), .C1(new_n661), .C2(KEYINPUT40), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n662), .B1(KEYINPUT40), .B2(new_n661), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  NAND2_X1  g478(.A1(new_n613), .A2(new_n616), .ZN(new_n665));
  INV_X1    g479(.A(new_n645), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n607), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n556), .A2(new_n643), .A3(new_n319), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(KEYINPUT97), .B(G146), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G48));
  NOR2_X1   g485(.A1(new_n308), .A2(KEYINPUT98), .ZN(new_n672));
  INV_X1    g486(.A(new_n299), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n280), .B1(new_n314), .B2(new_n288), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n672), .B1(new_n675), .B2(new_n191), .ZN(new_n676));
  OAI221_X1 g490(.A(new_n190), .B1(KEYINPUT98), .B2(new_n308), .C1(new_n673), .C2(new_n674), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n188), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n556), .A2(new_n618), .A3(new_n598), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT41), .B(G113), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT99), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G15));
  NAND4_X1  g497(.A1(new_n556), .A2(new_n598), .A3(new_n626), .A4(new_n679), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G116), .ZN(G18));
  AOI21_X1  g499(.A(new_n678), .B1(new_n325), .B2(new_n322), .ZN(new_n686));
  INV_X1    g500(.A(new_n489), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(new_n556), .A3(new_n687), .A4(new_n643), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  NAND2_X1  g503(.A1(new_n539), .A2(new_n190), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n536), .B(new_n538), .C1(new_n520), .C2(new_n552), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n690), .A2(G472), .B1(new_n540), .B2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n585), .B1(new_n593), .B2(new_n582), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n657), .B(new_n327), .C1(new_n376), .C2(new_n375), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n694), .A2(new_n686), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G122), .ZN(G24));
  NOR2_X1   g512(.A1(new_n678), .A2(new_n642), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n699), .A2(new_n692), .A3(new_n638), .A4(new_n668), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  OR2_X1    g515(.A1(new_n544), .A2(KEYINPUT103), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n544), .A2(KEYINPUT103), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n702), .A2(new_n543), .A3(new_n555), .A4(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n693), .A3(new_n668), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n654), .A2(new_n327), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(KEYINPUT100), .B1(new_n317), .B2(new_n300), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n308), .B(new_n190), .C1(new_n673), .C2(new_n674), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT100), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n305), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n189), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n708), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n305), .A2(new_n711), .A3(new_n710), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n711), .B1(new_n305), .B2(new_n710), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n188), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(KEYINPUT101), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n706), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n707), .B1(new_n718), .B2(KEYINPUT101), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n713), .A2(new_n714), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(KEYINPUT102), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n705), .B1(new_n720), .B2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n556), .A2(new_n598), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n715), .A2(new_n719), .A3(new_n706), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT102), .B1(new_n721), .B2(new_n722), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n225), .ZN(G33));
  OAI211_X1 g548(.A(new_n728), .B(new_n646), .C1(new_n730), .C2(new_n731), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n727), .B1(new_n720), .B2(new_n723), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT104), .A3(new_n646), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G134), .ZN(G36));
  NOR3_X1   g555(.A1(new_n617), .A2(new_n607), .A3(KEYINPUT43), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n617), .B1(new_n607), .B2(KEYINPUT106), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(KEYINPUT106), .B2(new_n607), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n742), .B1(new_n744), .B2(KEYINPUT43), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n605), .A2(new_n638), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(KEYINPUT107), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n316), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(KEYINPUT105), .A3(G469), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n755), .B1(new_n753), .B2(new_n316), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT105), .B1(new_n754), .B2(G469), .ZN(new_n757));
  OAI22_X1  g571(.A1(new_n756), .A2(new_n757), .B1(new_n308), .B2(new_n301), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT46), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n300), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n759), .B2(new_n758), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n188), .A3(new_n659), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n707), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n751), .A2(new_n752), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT108), .B(G137), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G39));
  NOR4_X1   g580(.A1(new_n556), .A2(new_n598), .A3(new_n667), .A4(new_n707), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT47), .B1(new_n761), .B2(new_n188), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  NOR2_X1   g585(.A1(G952), .A2(G953), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n680), .A2(new_n697), .A3(new_n684), .A4(new_n688), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n732), .B(new_n773), .C1(new_n725), .C2(new_n724), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n695), .A2(new_n645), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n652), .A3(new_n713), .A4(new_n637), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n778), .A2(new_n647), .A3(new_n669), .A4(new_n700), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n779), .A2(KEYINPUT52), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n307), .A2(new_n318), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n783), .A2(new_n188), .A3(new_n646), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n189), .B(new_n667), .C1(new_n318), .C2(new_n307), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n556), .B(new_n643), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT110), .A3(new_n700), .A4(new_n778), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n780), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n483), .A2(new_n488), .A3(new_n666), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n638), .A2(new_n791), .A3(new_n624), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n556), .A2(new_n792), .A3(new_n319), .A4(new_n708), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n720), .A2(new_n723), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n692), .A2(new_n638), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n668), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n319), .A2(new_n490), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n319), .A2(new_n490), .A3(new_n638), .ZN(new_n800));
  OAI22_X1  g614(.A1(new_n727), .A2(new_n799), .B1(new_n800), .B2(new_n605), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n617), .A2(new_n607), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n489), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n803), .A2(new_n377), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n601), .A2(new_n605), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n798), .B1(new_n801), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n803), .A2(new_n377), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n633), .A2(new_n598), .A3(new_n319), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n639), .A3(new_n599), .A4(KEYINPUT109), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n797), .A2(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n740), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n776), .A2(new_n790), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  INV_X1    g629(.A(new_n774), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n740), .A3(new_n811), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n788), .A2(new_n789), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n782), .A2(new_n787), .A3(KEYINPUT52), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n815), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n813), .A2(new_n814), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n813), .A2(KEYINPUT114), .A3(new_n821), .A4(new_n814), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n735), .A2(new_n736), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT104), .B1(new_n738), .B2(new_n646), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n797), .A2(new_n810), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n829), .A2(new_n774), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  INV_X1    g646(.A(new_n820), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT53), .A4(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n816), .A2(new_n811), .A3(new_n740), .A4(new_n790), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT111), .B1(new_n835), .B2(new_n815), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n810), .B(new_n797), .C1(new_n827), .C2(new_n828), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n837), .A2(new_n820), .A3(new_n815), .A4(new_n774), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT54), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n826), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n708), .A2(new_n324), .A3(new_n679), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n742), .B(new_n845), .C1(KEYINPUT43), .C2(new_n744), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n704), .A2(new_n693), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(KEYINPUT48), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n845), .A2(new_n652), .A3(new_n597), .A4(new_n594), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n607), .A3(new_n665), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n745), .A2(new_n694), .A3(new_n324), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n699), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n852), .A2(new_n854), .A3(G952), .A4(new_n276), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT118), .Z(new_n856));
  NOR2_X1   g670(.A1(new_n768), .A2(new_n769), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n676), .A2(new_n677), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n188), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n708), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT51), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n656), .A2(new_n327), .A3(new_n678), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n853), .A2(new_n864), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT50), .Z(new_n866));
  NAND3_X1  g680(.A1(new_n851), .A2(new_n608), .A3(new_n617), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT116), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n846), .A2(new_n795), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n850), .B(new_n856), .C1(new_n863), .C2(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n862), .A2(KEYINPUT115), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(KEYINPUT115), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n870), .A2(KEYINPUT117), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n772), .B1(new_n844), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n693), .A2(new_n188), .A3(new_n327), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n858), .B2(KEYINPUT49), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(KEYINPUT49), .B2(new_n858), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n882), .A2(new_n656), .A3(new_n652), .A4(new_n744), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT119), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n824), .A2(new_n825), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT112), .B1(new_n839), .B2(KEYINPUT54), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n839), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n885), .B(new_n878), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n772), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  INV_X1    g705(.A(new_n883), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n884), .A2(new_n893), .ZN(G75));
  NOR2_X1   g708(.A1(new_n276), .A2(G952), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n190), .B1(new_n813), .B2(new_n821), .ZN(new_n897));
  INV_X1    g711(.A(new_n374), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT56), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n354), .A2(new_n362), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n360), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT55), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n896), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n899), .B2(new_n902), .ZN(G51));
  NAND2_X1  g718(.A1(new_n813), .A2(new_n821), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n822), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n308), .A2(new_n301), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n675), .B1(new_n910), .B2(KEYINPUT120), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(KEYINPUT120), .B2(new_n910), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n756), .A2(new_n757), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n897), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n895), .B1(new_n912), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n441), .A2(new_n423), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n895), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n918), .B1(new_n917), .B2(new_n916), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT121), .Z(G60));
  XNOR2_X1  g734(.A(new_n477), .B(KEYINPUT33), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n824), .B(new_n825), .C1(new_n887), .C2(new_n886), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n922), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n925), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n927), .B1(new_n907), .B2(new_n929), .ZN(new_n930));
  AOI211_X1 g744(.A(KEYINPUT122), .B(new_n928), .C1(new_n906), .C2(new_n822), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n896), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT123), .B1(new_n926), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n921), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n844), .B2(new_n924), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT123), .ZN(new_n936));
  INV_X1    g750(.A(new_n822), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n814), .B1(new_n813), .B2(new_n821), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n929), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n907), .A2(new_n927), .A3(new_n929), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n895), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n935), .A2(new_n936), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n933), .A2(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT124), .Z(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n947), .B1(new_n813), .B2(new_n821), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n948), .A2(new_n635), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n949), .B(new_n896), .C1(new_n580), .C2(new_n948), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT61), .B1(new_n949), .B2(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G66));
  OAI21_X1  g766(.A(G953), .B1(new_n321), .B2(new_n358), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT126), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n810), .A2(new_n773), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n900), .B1(G898), .B2(new_n276), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  NAND3_X1  g773(.A1(new_n529), .A2(new_n532), .A3(new_n533), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n396), .A2(new_n398), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(new_n962));
  AND2_X1   g776(.A1(new_n786), .A2(new_n700), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n663), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n967));
  INV_X1    g781(.A(new_n770), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n661), .A2(new_n727), .A3(new_n707), .A4(new_n803), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n967), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n966), .A2(new_n970), .A3(new_n764), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n962), .B1(new_n971), .B2(new_n276), .ZN(new_n972));
  OR3_X1    g786(.A1(new_n762), .A2(new_n695), .A3(new_n847), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n973), .A2(new_n770), .A3(new_n963), .ZN(new_n974));
  INV_X1    g788(.A(new_n733), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n740), .A4(new_n764), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(G953), .ZN(new_n977));
  NAND2_X1  g791(.A1(G900), .A2(G953), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n977), .A2(new_n962), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n276), .B1(G227), .B2(G900), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n971), .B2(new_n955), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n649), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n976), .B2(new_n955), .ZN(new_n987));
  INV_X1    g801(.A(new_n546), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n895), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n984), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n988), .A2(new_n649), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n990), .B1(new_n839), .B2(new_n992), .ZN(G57));
endmodule


