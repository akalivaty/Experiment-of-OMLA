//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n589, new_n590, new_n591, new_n592, new_n593, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G131), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n191), .A3(new_n196), .A4(new_n192), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n200), .A2(new_n202), .A3(KEYINPUT0), .A4(G128), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT0), .B(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n198), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G134), .B2(new_n190), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n193), .A2(new_n209), .B1(new_n192), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n200), .A2(new_n202), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  NOR3_X1   g028(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n199), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT66), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT66), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n221), .B1(G128), .B2(new_n204), .ZN(new_n222));
  OAI22_X1  g036(.A1(new_n211), .A2(KEYINPUT67), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT30), .B(new_n208), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G119), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G116), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT2), .B(G113), .ZN(new_n231));
  OR2_X1    g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n231), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n206), .B1(new_n195), .B2(new_n197), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n193), .A2(new_n209), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n210), .A2(new_n192), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(new_n220), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n204), .A3(G128), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n214), .A2(new_n212), .B1(new_n213), .B2(new_n216), .ZN(new_n242));
  AOI22_X1  g056(.A1(new_n238), .A2(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n235), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n225), .B(new_n234), .C1(new_n245), .C2(KEYINPUT30), .ZN(new_n246));
  INV_X1    g060(.A(new_n234), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(new_n208), .C1(new_n223), .C2(new_n224), .ZN(new_n248));
  INV_X1    g062(.A(G237), .ZN(new_n249));
  INV_X1    g063(.A(G953), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G210), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n246), .A2(new_n248), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n246), .A2(new_n257), .A3(new_n248), .A4(new_n254), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(KEYINPUT31), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT31), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n248), .B1(new_n245), .B2(new_n247), .ZN(new_n263));
  XOR2_X1   g077(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n248), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n254), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(G472), .A2(G902), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(KEYINPUT32), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT72), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT32), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n268), .B1(new_n259), .B2(new_n261), .ZN(new_n275));
  INV_X1    g089(.A(new_n271), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n270), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n271), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n265), .A2(new_n267), .ZN(new_n282));
  INV_X1    g096(.A(new_n254), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n246), .A2(new_n248), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n283), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n267), .B(KEYINPUT71), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n208), .B1(new_n223), .B2(new_n224), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n234), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n248), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT28), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(KEYINPUT70), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n289), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n297));
  OAI221_X1 g111(.A(new_n281), .B1(new_n284), .B2(new_n288), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G472), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n280), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G234), .ZN(new_n301));
  OAI21_X1  g115(.A(G217), .B1(new_n301), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT16), .ZN(new_n303));
  INV_X1    g117(.A(G140), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G125), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(G125), .ZN(new_n306));
  INV_X1    g120(.A(G125), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n305), .B1(new_n309), .B2(new_n303), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(new_n199), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT73), .ZN(new_n312));
  OAI211_X1 g126(.A(G146), .B(new_n305), .C1(new_n309), .C2(new_n303), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n199), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT23), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n316), .B1(G119), .B2(new_n214), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n226), .A2(KEYINPUT23), .A3(G128), .ZN(new_n318));
  OAI22_X1  g132(.A1(new_n317), .A2(new_n318), .B1(G119), .B2(new_n214), .ZN(new_n319));
  XNOR2_X1  g133(.A(G119), .B(G128), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT24), .B(G110), .Z(new_n321));
  AOI22_X1  g135(.A1(new_n319), .A2(G110), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n314), .A2(new_n315), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n319), .A2(G110), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n321), .A2(new_n320), .ZN(new_n325));
  OAI221_X1 g139(.A(new_n313), .B1(G146), .B2(new_n309), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n250), .A2(G221), .A3(G234), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT74), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT22), .B(G137), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n323), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n323), .B2(new_n326), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G902), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n334), .A2(KEYINPUT25), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(KEYINPUT25), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n302), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n333), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n301), .B2(G217), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n300), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT20), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n314), .A2(KEYINPUT85), .A3(new_n315), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n249), .A2(new_n250), .A3(G214), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n346), .B(G143), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(new_n209), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT17), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT85), .B1(new_n314), .B2(new_n315), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n314), .A2(new_n315), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT85), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n355), .A2(KEYINPUT86), .A3(new_n345), .A4(new_n349), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n347), .B(new_n209), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n357), .A2(KEYINPUT17), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(G113), .B(G122), .ZN(new_n360));
  INV_X1    g174(.A(G104), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n360), .B(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n348), .A2(KEYINPUT18), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT18), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n347), .B1(new_n364), .B2(new_n209), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n309), .B(G146), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n359), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n309), .B(KEYINPUT19), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n357), .B(new_n313), .C1(G146), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n367), .ZN(new_n371));
  INV_X1    g185(.A(new_n362), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(G475), .A2(G902), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n343), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n375), .ZN(new_n377));
  AOI211_X1 g191(.A(KEYINPUT20), .B(new_n377), .C1(new_n368), .C2(new_n373), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n359), .A2(new_n367), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n372), .ZN(new_n380));
  AOI21_X1  g194(.A(G902), .B1(new_n380), .B2(new_n368), .ZN(new_n381));
  INV_X1    g195(.A(G475), .ZN(new_n382));
  OAI22_X1  g196(.A1(new_n376), .A2(new_n378), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G128), .B(G143), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(new_n188), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n228), .A2(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n228), .A2(G122), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(KEYINPUT14), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G107), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n386), .B(new_n387), .C1(KEYINPUT14), .C2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n385), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n388), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT87), .B(G107), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n188), .A2(KEYINPUT13), .ZN(new_n396));
  AOI22_X1  g210(.A1(new_n394), .A2(new_n395), .B1(new_n384), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n394), .B2(new_n395), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(G128), .B2(new_n201), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n385), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n393), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT9), .B(G234), .Z(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G217), .A3(new_n250), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(KEYINPUT88), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n404), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n406), .B(new_n393), .C1(new_n400), .C2(new_n398), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(KEYINPUT15), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n408), .B(KEYINPUT89), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(new_n414), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n383), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n242), .A2(new_n307), .A3(new_n241), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n242), .A2(new_n422), .A3(new_n307), .A4(new_n241), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n206), .A2(G125), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G224), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n428), .B2(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n420), .A2(KEYINPUT82), .B1(G125), .B2(new_n206), .ZN(new_n433));
  INV_X1    g247(.A(new_n427), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n433), .A2(KEYINPUT7), .A3(new_n434), .A4(new_n423), .ZN(new_n435));
  INV_X1    g249(.A(G101), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT3), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n391), .A3(G104), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT3), .B1(new_n361), .B2(G107), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n361), .A2(G107), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n436), .B(new_n438), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n391), .A2(G104), .ZN(new_n442));
  OAI21_X1  g256(.A(G101), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT5), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(G113), .C1(KEYINPUT5), .C2(new_n227), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n232), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n232), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n444), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT8), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n432), .A2(new_n435), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n438), .B1(new_n439), .B2(new_n440), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G101), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(KEYINPUT4), .A3(new_n441), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n441), .A2(KEYINPUT4), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n437), .B1(new_n391), .B2(G104), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n391), .A2(G104), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n436), .B1(new_n462), .B2(new_n438), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n458), .A2(new_n464), .A3(new_n234), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n465), .A2(new_n448), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n455), .A2(KEYINPUT84), .B1(new_n452), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT84), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n432), .A2(new_n435), .A3(new_n454), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n425), .B(new_n427), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n452), .B1(new_n465), .B2(new_n448), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT6), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n466), .A2(new_n452), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n472), .A2(new_n473), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT81), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(KEYINPUT81), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n471), .B(new_n476), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n470), .A2(new_n281), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n467), .B2(new_n469), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n483), .A3(new_n481), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(G214), .B1(G237), .B2(G902), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G952), .ZN(new_n492));
  AOI211_X1 g306(.A(G953), .B(new_n492), .C1(G234), .C2(G237), .ZN(new_n493));
  XOR2_X1   g307(.A(KEYINPUT21), .B(G898), .Z(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  AOI211_X1 g309(.A(new_n281), .B(new_n250), .C1(G234), .C2(G237), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n419), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  XOR2_X1   g314(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n501));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n241), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n240), .A2(new_n204), .A3(KEYINPUT76), .A4(G128), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n212), .A2(new_n214), .B1(KEYINPUT1), .B2(new_n216), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT77), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n506), .A2(new_n507), .A3(new_n445), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n506), .B2(new_n445), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n198), .ZN(new_n511));
  OAI21_X1  g325(.A(KEYINPUT10), .B1(new_n215), .B2(new_n222), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT79), .B1(new_n512), .B2(new_n444), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n242), .A2(new_n241), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT79), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n514), .A2(new_n445), .A3(new_n515), .A4(KEYINPUT10), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n459), .A2(new_n463), .ZN(new_n517));
  AOI211_X1 g331(.A(KEYINPUT4), .B(new_n436), .C1(new_n462), .C2(new_n438), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n513), .A2(new_n516), .B1(new_n519), .B2(new_n207), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n510), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n250), .A2(G227), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n522), .B(KEYINPUT75), .ZN(new_n523));
  XNOR2_X1  g337(.A(G110), .B(G140), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n508), .A2(new_n509), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n514), .A2(new_n445), .ZN(new_n528));
  OAI211_X1 g342(.A(KEYINPUT12), .B(new_n198), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT12), .ZN(new_n530));
  INV_X1    g344(.A(new_n509), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n506), .A2(new_n507), .A3(new_n445), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n530), .B1(new_n533), .B2(new_n511), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n526), .B1(new_n529), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n511), .B1(new_n510), .B2(new_n520), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n525), .B1(new_n537), .B2(new_n521), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n500), .B(new_n281), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n525), .A3(new_n521), .ZN(new_n540));
  INV_X1    g354(.A(new_n521), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n541), .B1(new_n529), .B2(new_n534), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n540), .B(G469), .C1(new_n542), .C2(new_n525), .ZN(new_n543));
  NAND2_X1  g357(.A1(G469), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n539), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G221), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n402), .B2(new_n281), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT80), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT80), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n545), .A2(new_n551), .A3(new_n548), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n342), .A2(new_n499), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT91), .B(G101), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(G3));
  NAND2_X1  g371(.A1(new_n270), .A2(new_n271), .ZN(new_n558));
  OAI21_X1  g372(.A(G472), .B1(new_n275), .B2(G902), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n553), .A2(new_n341), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT92), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n485), .A2(new_n562), .A3(new_n487), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n483), .B1(new_n486), .B2(new_n481), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n490), .B1(new_n564), .B2(KEYINPUT92), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n405), .A2(new_n407), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n570), .A2(KEYINPUT93), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(KEYINPUT93), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n405), .B2(KEYINPUT94), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n571), .A2(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(G478), .A3(new_n281), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n416), .A2(new_n410), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n580), .B1(new_n416), .B2(new_n410), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n577), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n383), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(new_n497), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n567), .A2(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(KEYINPUT96), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT34), .B(G104), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G6));
  NOR2_X1   g402(.A1(new_n383), .A2(new_n417), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n497), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n567), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(KEYINPUT35), .B(G107), .Z(new_n593));
  XNOR2_X1  g407(.A(new_n592), .B(new_n593), .ZN(G9));
  NAND2_X1  g408(.A1(new_n323), .A2(new_n326), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n330), .A2(KEYINPUT36), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(new_n339), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n337), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n499), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n553), .A3(new_n560), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT37), .B(G110), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G12));
  AOI21_X1  g417(.A(new_n599), .B1(new_n550), .B2(new_n552), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n376), .A2(new_n378), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n381), .A2(new_n382), .ZN(new_n606));
  INV_X1    g420(.A(G900), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n496), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n493), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n605), .A2(new_n606), .A3(new_n418), .A4(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT97), .B1(new_n611), .B2(new_n566), .ZN(new_n612));
  INV_X1    g426(.A(new_n566), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n589), .A3(new_n614), .A4(new_n610), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n300), .A2(new_n604), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(G128), .ZN(G30));
  XOR2_X1   g431(.A(new_n610), .B(KEYINPUT39), .Z(new_n618));
  OR3_X1    g432(.A1(new_n554), .A2(KEYINPUT40), .A3(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n256), .A2(new_n258), .B1(new_n292), .B2(new_n283), .ZN(new_n620));
  OAI21_X1  g434(.A(G472), .B1(new_n620), .B2(G902), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n280), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT40), .B1(new_n554), .B2(new_n618), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n488), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n383), .A2(new_n418), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n599), .A2(new_n489), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n619), .A2(new_n622), .A3(new_n623), .A4(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G143), .ZN(G45));
  NAND3_X1  g444(.A1(new_n582), .A2(new_n383), .A3(new_n610), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n566), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n300), .A2(new_n604), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G146), .ZN(G48));
  OAI21_X1  g448(.A(new_n281), .B1(new_n535), .B2(new_n538), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G469), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n548), .A3(new_n539), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n566), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g452(.A1(new_n300), .A2(new_n341), .A3(new_n584), .A4(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT41), .B(G113), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G15));
  NAND4_X1  g455(.A1(new_n300), .A2(new_n591), .A3(new_n341), .A4(new_n638), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT99), .B(G116), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G18));
  NOR4_X1   g458(.A1(new_n383), .A2(new_n599), .A3(new_n497), .A4(new_n418), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n300), .A2(new_n638), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G119), .ZN(G21));
  NOR4_X1   g461(.A1(new_n626), .A2(new_n566), .A3(new_n637), .A4(new_n497), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n296), .A2(new_n283), .B1(new_n261), .B2(new_n259), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n276), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n559), .ZN(new_n652));
  INV_X1    g466(.A(new_n341), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n650), .A2(new_n649), .A3(new_n276), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT101), .B(G122), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G24));
  NOR3_X1   g472(.A1(new_n652), .A2(new_n599), .A3(new_n654), .ZN(new_n659));
  INV_X1    g473(.A(new_n631), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n659), .A2(new_n660), .A3(new_n638), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G125), .ZN(G27));
  NAND2_X1  g476(.A1(new_n488), .A2(new_n489), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n549), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n300), .A2(new_n341), .A3(new_n660), .A4(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(KEYINPUT102), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n665), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n277), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(KEYINPUT103), .B2(new_n272), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n299), .B1(new_n674), .B2(new_n277), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n341), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(KEYINPUT42), .A3(new_n660), .A4(new_n664), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G131), .ZN(G33));
  NOR3_X1   g494(.A1(new_n342), .A2(new_n549), .A3(new_n663), .ZN(new_n681));
  INV_X1    g495(.A(new_n611), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G134), .ZN(G36));
  INV_X1    g498(.A(new_n383), .ZN(new_n685));
  AOI21_X1  g499(.A(KEYINPUT43), .B1(new_n685), .B2(new_n582), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n383), .A2(KEYINPUT105), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n383), .A2(KEYINPUT105), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(KEYINPUT43), .A3(new_n582), .A4(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n688), .A2(new_n582), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n692), .A2(KEYINPUT106), .A3(KEYINPUT43), .A4(new_n687), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n686), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n694), .A2(new_n560), .A3(new_n599), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n540), .B1(new_n542), .B2(new_n525), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT45), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n500), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n698), .B2(new_n697), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(KEYINPUT46), .A3(new_n544), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n539), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT46), .B1(new_n700), .B2(new_n544), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n548), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n704), .A2(new_n618), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n705), .A2(new_n706), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n663), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n696), .B(new_n709), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G137), .ZN(G39));
  AND2_X1   g528(.A1(new_n704), .A2(KEYINPUT47), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n704), .A2(KEYINPUT47), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n663), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n660), .A2(new_n653), .A3(new_n718), .ZN(new_n719));
  OR4_X1    g533(.A1(new_n300), .A2(new_n715), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G140), .ZN(G42));
  NAND3_X1  g535(.A1(new_n341), .A2(new_n489), .A3(new_n548), .ZN(new_n722));
  INV_X1    g536(.A(new_n625), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n636), .A2(new_n539), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT108), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n722), .B(new_n723), .C1(KEYINPUT49), .C2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n622), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n692), .A2(new_n687), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n725), .A2(KEYINPUT49), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(new_n727), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  AOI22_X1  g544(.A1(new_n671), .A2(new_n678), .B1(new_n682), .B2(new_n681), .ZN(new_n731));
  INV_X1    g545(.A(new_n583), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n491), .B(new_n498), .C1(new_n732), .C2(new_n589), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n601), .B1(new_n561), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n604), .A2(new_n419), .A3(new_n610), .A4(new_n718), .ZN(new_n736));
  INV_X1    g550(.A(new_n300), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n734), .A2(new_n738), .A3(new_n555), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n642), .A2(new_n639), .A3(new_n646), .A4(new_n656), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n731), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n545), .A2(new_n599), .A3(new_n548), .A4(new_n610), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n626), .A3(new_n566), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n622), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n616), .A2(new_n633), .A3(new_n661), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(KEYINPUT111), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT111), .B1(new_n747), .B2(new_n748), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n616), .A2(new_n633), .A3(new_n661), .A4(new_n746), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT110), .B1(new_n747), .B2(new_n748), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n751), .A2(KEYINPUT112), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT112), .B1(new_n751), .B2(new_n756), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n743), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n752), .A2(KEYINPUT52), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n747), .A2(new_n748), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n740), .B(KEYINPUT109), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n731), .A2(new_n763), .A3(new_n764), .A4(new_n739), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n741), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n759), .A2(new_n760), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT113), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n759), .A2(new_n769), .A3(new_n760), .A4(new_n766), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n741), .A2(new_n731), .A3(new_n764), .A4(new_n739), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n758), .B2(new_n757), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n765), .A2(KEYINPUT53), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(KEYINPUT54), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n694), .A2(new_n609), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(new_n638), .A3(new_n655), .ZN(new_n776));
  INV_X1    g590(.A(new_n637), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n718), .A2(new_n777), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n622), .A2(new_n778), .A3(new_n653), .A4(new_n609), .ZN(new_n779));
  AOI211_X1 g593(.A(new_n492), .B(G953), .C1(new_n779), .C2(new_n732), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n776), .A2(new_n780), .A3(KEYINPUT117), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT117), .B1(new_n776), .B2(new_n780), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT48), .ZN(new_n784));
  NOR4_X1   g598(.A1(new_n694), .A2(new_n676), .A3(new_n609), .A4(new_n778), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n784), .B1(new_n785), .B2(KEYINPUT118), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(KEYINPUT118), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n785), .A2(KEYINPUT118), .A3(new_n784), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n783), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n777), .A2(new_n490), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n625), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n775), .A2(new_n655), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT50), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n795), .B1(KEYINPUT115), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n775), .A2(new_n655), .A3(new_n798), .A4(new_n794), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  OAI22_X1  g615(.A1(new_n717), .A2(new_n715), .B1(new_n548), .B2(new_n725), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n655), .A3(new_n718), .A4(new_n775), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n582), .A2(new_n383), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n779), .A2(new_n804), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(KEYINPUT116), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n694), .A2(new_n609), .A3(new_n778), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n806), .A2(new_n807), .B1(new_n659), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n801), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT51), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n801), .A2(new_n812), .A3(new_n803), .A4(new_n809), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n790), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n768), .A2(new_n770), .A3(new_n774), .A4(new_n814), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n815), .A2(KEYINPUT119), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n492), .A2(new_n250), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n815), .B2(KEYINPUT119), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n730), .B1(new_n816), .B2(new_n818), .ZN(G75));
  AOI21_X1  g633(.A(new_n281), .B1(new_n759), .B2(new_n766), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(G210), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n476), .B1(new_n479), .B2(new_n480), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(new_n471), .ZN(new_n824));
  XOR2_X1   g638(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n821), .A2(new_n822), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n821), .B2(new_n822), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n250), .A2(G952), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(G51));
  NAND3_X1  g644(.A1(new_n731), .A2(new_n739), .A3(new_n742), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n754), .A2(new_n755), .ZN(new_n833));
  INV_X1    g647(.A(new_n750), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n747), .A2(KEYINPUT111), .A3(new_n748), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n751), .A2(new_n756), .A3(KEYINPUT112), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n831), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n765), .A2(new_n741), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT54), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n767), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n759), .A2(new_n766), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(KEYINPUT121), .A3(KEYINPUT54), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n544), .B(KEYINPUT57), .Z(new_n846));
  NAND3_X1  g660(.A1(new_n843), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n538), .B2(new_n535), .ZN(new_n848));
  INV_X1    g662(.A(new_n820), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(new_n700), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n829), .B1(new_n848), .B2(new_n850), .ZN(G54));
  NAND2_X1  g665(.A1(KEYINPUT58), .A2(G475), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n820), .A2(new_n374), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n374), .B1(new_n820), .B2(new_n853), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n854), .A2(new_n855), .A3(new_n829), .ZN(G60));
  XNOR2_X1  g670(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n410), .A2(new_n281), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n843), .A2(new_n576), .A3(new_n845), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n829), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n768), .A2(new_n770), .A3(new_n774), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n576), .B1(new_n863), .B2(new_n859), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(G63));
  NAND2_X1  g679(.A1(G217), .A2(G902), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT60), .Z(new_n867));
  NAND2_X1  g681(.A1(new_n844), .A2(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n333), .B(KEYINPUT123), .Z(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n844), .A2(new_n597), .A3(new_n867), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n861), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n872), .B(new_n873), .ZN(G66));
  OAI21_X1  g688(.A(G953), .B1(new_n495), .B2(new_n426), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n734), .A2(new_n555), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n764), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n877), .B2(G953), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n823), .B1(G898), .B2(new_n250), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(G69));
  AND3_X1   g694(.A1(new_n616), .A2(new_n633), .A3(new_n661), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n629), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT62), .ZN(new_n883));
  INV_X1    g697(.A(new_n342), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n554), .A2(new_n618), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n663), .B1(new_n590), .B2(new_n583), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n883), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n888), .A2(new_n713), .A3(new_n720), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n225), .B1(new_n245), .B2(KEYINPUT30), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(new_n369), .Z(new_n891));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n250), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n891), .ZN(new_n893));
  OAI21_X1  g707(.A(G900), .B1(new_n893), .B2(G227), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(G953), .ZN(new_n895));
  INV_X1    g709(.A(new_n881), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n707), .A2(new_n708), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n676), .A2(new_n566), .A3(new_n626), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n713), .A2(new_n720), .A3(new_n731), .A4(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n250), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n893), .B1(G227), .B2(new_n250), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n892), .B(new_n895), .C1(new_n901), .C2(new_n902), .ZN(G72));
  NAND2_X1  g717(.A1(G472), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT63), .Z(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT124), .ZN(new_n906));
  INV_X1    g720(.A(new_n877), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n900), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n285), .B(KEYINPUT125), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n283), .A3(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n888), .A2(new_n713), .A3(new_n720), .A4(new_n877), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(new_n906), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n909), .A2(new_n283), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n910), .B(new_n861), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n772), .A2(new_n773), .ZN(new_n915));
  INV_X1    g729(.A(new_n905), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n256), .A2(new_n258), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(new_n286), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT126), .Z(new_n919));
  NOR2_X1   g733(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(KEYINPUT127), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n914), .B1(new_n921), .B2(new_n922), .ZN(G57));
endmodule


