//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(KEYINPUT32), .ZN(new_n188));
  INV_X1    g002(.A(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G146), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n191), .A2(G143), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n193), .A2(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(new_n189), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n195), .A2(new_n199), .A3(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT11), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT11), .A3(G134), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n204), .A2(G137), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n205), .A2(new_n207), .A3(new_n208), .A4(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n209), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n204), .A2(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(G131), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n202), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n209), .A3(new_n207), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT0), .A2(G128), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n200), .A2(new_n196), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n192), .A2(new_n194), .A3(new_n217), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n216), .A2(new_n210), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n214), .B1(new_n222), .B2(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n216), .A2(new_n210), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n221), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n224), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT30), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT30), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n224), .A2(KEYINPUT64), .A3(new_n225), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT64), .B1(new_n224), .B2(new_n225), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n228), .B(new_n214), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G116), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT65), .B(G116), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G119), .ZN(new_n237));
  XOR2_X1   g051(.A(KEYINPUT2), .B(G113), .Z(new_n238));
  XNOR2_X1  g052(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n223), .A2(new_n226), .A3(new_n239), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT67), .A2(G953), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT67), .A2(G953), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G237), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(G210), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT27), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT26), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT27), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n246), .A2(new_n251), .A3(G210), .A4(new_n247), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n249), .B2(new_n252), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n243), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n255), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(G101), .A3(new_n253), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n240), .A2(new_n242), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT31), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n241), .B1(new_n232), .B2(new_n239), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT31), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n214), .B1(new_n229), .B2(new_n230), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n239), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n242), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n224), .A2(new_n225), .ZN(new_n271));
  INV_X1    g085(.A(G116), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT65), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT65), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G116), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n275), .A3(G119), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n238), .A2(new_n276), .A3(new_n234), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n238), .B1(new_n234), .B2(new_n276), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n271), .A2(new_n279), .A3(new_n214), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n267), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(KEYINPUT68), .A3(new_n267), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n259), .B1(new_n270), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT69), .B1(new_n266), .B2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT31), .B1(new_n264), .B2(new_n260), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n279), .B1(new_n227), .B2(new_n231), .ZN(new_n289));
  NOR4_X1   g103(.A1(new_n289), .A2(new_n262), .A3(new_n259), .A4(new_n241), .ZN(new_n290));
  OAI211_X1 g104(.A(KEYINPUT69), .B(new_n286), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n188), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT71), .B1(new_n264), .B2(new_n260), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n283), .A2(new_n284), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n241), .B1(new_n239), .B2(new_n268), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n295), .B(new_n260), .C1(new_n267), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n299), .B(new_n259), .C1(new_n289), .C2(new_n241), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n294), .A2(new_n297), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n223), .ZN(new_n302));
  INV_X1    g116(.A(new_n226), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n279), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT28), .B1(new_n304), .B2(new_n241), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n259), .A2(new_n298), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n295), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n295), .A2(new_n305), .A3(KEYINPUT72), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G902), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n301), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G472), .ZN(new_n314));
  INV_X1    g128(.A(new_n187), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT69), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n315), .B1(new_n318), .B2(new_n291), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n320));
  OAI211_X1 g134(.A(new_n293), .B(new_n314), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G140), .ZN(new_n324));
  INV_X1    g138(.A(G140), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n326), .A3(KEYINPUT74), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n325), .A2(KEYINPUT74), .A3(G125), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n322), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n326), .A2(KEYINPUT16), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n191), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n330), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n325), .A2(KEYINPUT74), .A3(G125), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n334), .B2(KEYINPUT74), .ZN(new_n335));
  OAI211_X1 g149(.A(G146), .B(new_n332), .C1(new_n335), .C2(new_n322), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n233), .A2(G128), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n189), .A2(KEYINPUT23), .A3(G119), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n233), .A2(G128), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n338), .B(new_n339), .C1(new_n340), .C2(KEYINPUT23), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n341), .A2(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(KEYINPUT73), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G110), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n189), .A2(G119), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n338), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT24), .B(G110), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n337), .B(new_n344), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n334), .A2(new_n191), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n347), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n341), .B2(G110), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n336), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n246), .ZN(new_n354));
  NAND2_X1  g168(.A1(G221), .A2(G234), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT22), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OR4_X1    g170(.A1(KEYINPUT22), .A2(new_n244), .A3(new_n245), .A4(new_n355), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(new_n206), .ZN(new_n359));
  AOI21_X1  g173(.A(G137), .B1(new_n356), .B2(new_n357), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n352), .A3(new_n361), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n363), .A2(new_n312), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n366));
  INV_X1    g180(.A(G217), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(G234), .B2(new_n312), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n363), .A2(new_n364), .A3(new_n369), .A4(new_n312), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n366), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n363), .A2(new_n364), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n368), .A2(G902), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT75), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n321), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(G113), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(KEYINPUT67), .A2(G953), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT67), .A2(G953), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(G214), .A3(new_n247), .A4(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT84), .B(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g199(.A1(KEYINPUT84), .A2(G143), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n246), .A2(G214), .A3(new_n247), .A4(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT18), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n385), .B(new_n387), .C1(new_n388), .C2(new_n208), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n327), .A2(new_n328), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n349), .B1(new_n390), .B2(new_n191), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AOI211_X1 g206(.A(new_n388), .B(new_n208), .C1(new_n385), .C2(new_n387), .ZN(new_n393));
  OAI21_X1  g207(.A(KEYINPUT85), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n385), .A2(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(KEYINPUT18), .A3(G131), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n389), .A4(new_n391), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(G131), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n385), .A2(new_n387), .A3(new_n208), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n334), .A2(KEYINPUT19), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n390), .B2(KEYINPUT19), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n402), .B(new_n336), .C1(G146), .C2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n380), .B1(new_n399), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT86), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT17), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n208), .C1(new_n385), .C2(new_n387), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n337), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n400), .A2(new_n408), .A3(new_n401), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n399), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n380), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n407), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n394), .A2(new_n398), .B1(new_n410), .B2(new_n411), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT86), .A3(new_n380), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n406), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(G475), .A2(G902), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT20), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT86), .B1(new_n416), .B2(new_n380), .ZN(new_n422));
  AND4_X1   g236(.A1(KEYINPUT86), .A2(new_n399), .A3(new_n380), .A4(new_n412), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n399), .A2(new_n405), .ZN(new_n424));
  OAI22_X1  g238(.A1(new_n422), .A2(new_n423), .B1(new_n380), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT20), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n425), .A2(new_n426), .A3(new_n419), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n422), .A2(new_n423), .B1(new_n380), .B2(new_n416), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n312), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G475), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n189), .A2(G143), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n193), .A2(G128), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(new_n204), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n236), .A2(G122), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n272), .A2(G122), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT14), .ZN(new_n440));
  OAI21_X1  g254(.A(G107), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  OAI221_X1 g255(.A(new_n435), .B1(G107), .B2(new_n438), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n443));
  INV_X1    g257(.A(new_n432), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT13), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n433), .B1(new_n444), .B2(new_n445), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n432), .A2(KEYINPUT87), .A3(KEYINPUT13), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G134), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n434), .A2(new_n204), .ZN(new_n451));
  INV_X1    g265(.A(G107), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n436), .B2(new_n437), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n438), .A2(G107), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n450), .B(new_n451), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT9), .B(G234), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n456), .A2(new_n367), .A3(G953), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n442), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n442), .B2(new_n455), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n462), .A2(KEYINPUT15), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n312), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n463), .B1(new_n460), .B2(G902), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G952), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(G953), .ZN(new_n469));
  INV_X1    g283(.A(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n247), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n312), .B(new_n246), .C1(G234), .C2(G237), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT21), .B(G898), .Z(new_n474));
  OAI21_X1  g288(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(new_n475), .B(KEYINPUT88), .Z(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n428), .A2(new_n431), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G210), .B1(G237), .B2(G902), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n225), .A2(G125), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n202), .A2(new_n323), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT83), .ZN(new_n485));
  INV_X1    g299(.A(G224), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n486), .A2(G953), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT83), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n482), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n485), .B2(new_n489), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n276), .A2(KEYINPUT5), .A3(new_n234), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n234), .A2(KEYINPUT5), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(G113), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n237), .A2(new_n238), .ZN(new_n496));
  OAI21_X1  g310(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT3), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n452), .A3(G104), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n379), .A2(G107), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n243), .A4(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT76), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n379), .B2(G107), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n452), .A2(KEYINPUT76), .A3(G104), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G101), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n495), .A2(new_n496), .A3(new_n501), .A4(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT4), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(G101), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n277), .B2(new_n278), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n508), .A2(G101), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT4), .A3(new_n501), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n507), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n239), .A2(new_n513), .A3(new_n510), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(KEYINPUT82), .A3(new_n507), .ZN(new_n519));
  XNOR2_X1  g333(.A(G110), .B(G122), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n507), .A3(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n520), .B1(new_n515), .B2(new_n516), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n519), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n492), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n520), .B(KEYINPUT8), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n506), .A2(new_n501), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n496), .B2(new_n495), .ZN(new_n532));
  INV_X1    g346(.A(new_n507), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT7), .B1(new_n486), .B2(G953), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n484), .B(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n523), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n312), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n481), .B1(new_n528), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n492), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n519), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n526), .A2(new_n519), .B1(KEYINPUT6), .B2(new_n523), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n540), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n538), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n480), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n539), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G214), .B1(G237), .B2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G469), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT10), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n195), .A2(KEYINPUT77), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n189), .A2(new_n200), .B1(new_n196), .B2(new_n198), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT77), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(new_n554), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n551), .B1(new_n556), .B2(new_n530), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT78), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n216), .A2(new_n558), .A3(new_n210), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n216), .B2(new_n210), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n513), .A2(new_n225), .A3(new_n510), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n551), .B1(new_n553), .B2(new_n195), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n531), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n557), .A2(new_n561), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT79), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n501), .A3(new_n506), .ZN(new_n568));
  AOI22_X1  g382(.A1(new_n568), .A2(new_n551), .B1(new_n531), .B2(new_n563), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT79), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n562), .A4(new_n561), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n566), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n202), .B1(new_n501), .B2(new_n506), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n531), .B2(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n224), .A2(KEYINPUT80), .ZN(new_n575));
  OAI21_X1  g389(.A(KEYINPUT12), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n568), .B1(new_n202), .B2(new_n531), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n578));
  INV_X1    g392(.A(new_n575), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n246), .A2(G227), .ZN(new_n582));
  XOR2_X1   g396(.A(G110), .B(G140), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n572), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n569), .A2(new_n562), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n224), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n585), .B1(new_n572), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n550), .B(new_n312), .C1(new_n586), .C2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n572), .A2(new_n585), .A3(new_n588), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n576), .A2(new_n580), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n592), .B1(new_n571), .B2(new_n566), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n591), .B(G469), .C1(new_n593), .C2(new_n585), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n550), .A2(new_n312), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n590), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G221), .B1(new_n456), .B2(G902), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n597), .A2(KEYINPUT81), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT81), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n479), .B(new_n549), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n377), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(new_n243), .ZN(G3));
  AND4_X1   g417(.A1(new_n376), .A2(new_n546), .A3(new_n547), .A4(new_n476), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n599), .B2(new_n600), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n187), .B1(new_n287), .B2(new_n292), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n318), .B2(new_n291), .ZN(new_n607));
  INV_X1    g421(.A(G472), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n421), .A2(new_n427), .B1(new_n430), .B2(G475), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n461), .A2(new_n312), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n462), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n460), .B(KEYINPUT33), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n462), .A2(G902), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  OR3_X1    g432(.A1(new_n611), .A2(KEYINPUT89), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT89), .B1(new_n611), .B2(new_n618), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT90), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n622), .B(new_n624), .ZN(G6));
  INV_X1    g439(.A(KEYINPUT91), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n421), .A2(new_n427), .A3(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT91), .B(KEYINPUT20), .C1(new_n418), .C2(new_n420), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n431), .A2(new_n467), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR3_X1   g448(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT36), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n353), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n348), .A3(new_n352), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n374), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT92), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT93), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n641), .A2(new_n642), .A3(new_n371), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n641), .B2(new_n371), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n645), .B(new_n606), .C1(new_n608), .C2(new_n607), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n601), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT37), .B(G110), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G12));
  NAND2_X1  g463(.A1(new_n597), .A2(new_n598), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT81), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n597), .A2(KEYINPUT81), .A3(new_n598), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n548), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n471), .ZN(new_n655));
  INV_X1    g469(.A(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n472), .B2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n629), .A2(new_n630), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n654), .A2(new_n658), .A3(new_n321), .A4(new_n645), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT94), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n643), .A2(new_n644), .ZN(new_n661));
  INV_X1    g475(.A(new_n320), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n606), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n318), .A2(new_n291), .ZN(new_n664));
  AOI22_X1  g478(.A1(new_n664), .A2(new_n188), .B1(new_n313), .B2(G472), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n661), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT94), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n654), .A4(new_n658), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT95), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n189), .ZN(G30));
  NAND2_X1  g485(.A1(new_n652), .A2(new_n653), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n657), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(new_n674), .B(KEYINPUT40), .Z(new_n675));
  OAI21_X1  g489(.A(new_n259), .B1(new_n304), .B2(new_n241), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT96), .Z(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n677), .B2(new_n261), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n293), .B1(new_n608), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n320), .B1(new_n664), .B2(new_n187), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n467), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n611), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n546), .B(KEYINPUT38), .Z(new_n685));
  INV_X1    g499(.A(new_n547), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n641), .A2(new_n371), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n675), .A2(new_n682), .A3(new_n684), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NOR3_X1   g504(.A1(new_n611), .A2(new_n618), .A3(new_n657), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n654), .A2(new_n321), .A3(new_n645), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT97), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n666), .A2(KEYINPUT97), .A3(new_n654), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  INV_X1    g511(.A(new_n376), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n698), .B1(new_n663), .B2(new_n665), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n586), .A2(new_n589), .ZN(new_n700));
  OAI21_X1  g514(.A(G469), .B1(new_n700), .B2(G902), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n701), .A2(new_n598), .A3(new_n590), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n702), .A2(new_n548), .A3(new_n477), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n621), .A2(new_n699), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  NAND3_X1  g520(.A1(new_n699), .A2(new_n631), .A3(new_n703), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G116), .ZN(G18));
  INV_X1    g522(.A(new_n702), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n549), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(new_n321), .A3(new_n479), .A4(new_n645), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  OAI21_X1  g527(.A(new_n312), .B1(new_n287), .B2(new_n292), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n295), .A2(new_n305), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n266), .B1(new_n260), .B2(new_n715), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n714), .A2(G472), .B1(new_n187), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n717), .A2(new_n703), .A3(new_n376), .A4(new_n684), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  INV_X1    g533(.A(new_n691), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n187), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n721), .B(new_n687), .C1(new_n607), .C2(new_n608), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n720), .A2(new_n722), .A3(new_n710), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n323), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT99), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n594), .A2(KEYINPUT98), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n572), .A2(new_n581), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n584), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT98), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(G469), .A4(new_n591), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n726), .A2(new_n590), .A3(new_n596), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(new_n598), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n686), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n539), .A2(new_n545), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n725), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n731), .A2(new_n734), .A3(new_n725), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n699), .A3(new_n691), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n731), .A2(new_n734), .A3(new_n725), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n735), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n691), .A2(KEYINPUT42), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n293), .A2(new_n314), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n319), .A2(KEYINPUT32), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n376), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n739), .A2(new_n740), .B1(new_n744), .B2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT100), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(new_n208), .ZN(G33));
  NAND3_X1  g565(.A1(new_n738), .A2(new_n699), .A3(new_n658), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT101), .B(G134), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G36));
  NAND2_X1  g568(.A1(new_n611), .A2(new_n617), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n755), .B1(KEYINPUT103), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n758));
  NAND3_X1  g572(.A1(new_n611), .A2(new_n617), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT104), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n609), .A2(new_n687), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n728), .A2(new_n591), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n550), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT102), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n768), .B1(new_n774), .B2(new_n595), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n772), .B(KEYINPUT102), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT46), .A3(new_n596), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(new_n590), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n778), .A2(new_n598), .A3(new_n673), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n762), .A2(KEYINPUT44), .A3(new_n763), .A4(new_n764), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n539), .A2(new_n545), .A3(new_n547), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT105), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n767), .A2(new_n780), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n778), .B2(new_n598), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n778), .A2(new_n786), .A3(new_n598), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n720), .A2(new_n321), .A3(new_n376), .A4(new_n782), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT106), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND2_X1  g607(.A1(new_n701), .A2(new_n590), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n376), .B(new_n733), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n755), .ZN(new_n798));
  XOR2_X1   g612(.A(new_n798), .B(KEYINPUT107), .Z(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n796), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(KEYINPUT108), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT108), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n685), .ZN(new_n803));
  OR4_X1    g617(.A1(new_n682), .A2(new_n799), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n539), .A2(new_n545), .A3(new_n547), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n709), .A2(new_n655), .A3(new_n805), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n761), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n722), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n682), .A2(new_n698), .A3(new_n806), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n611), .A2(new_n618), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g625(.A1(new_n788), .A2(new_n789), .B1(new_n732), .B2(new_n795), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n760), .A2(new_n376), .A3(new_n655), .A4(new_n717), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n783), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT114), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n811), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n685), .A2(new_n686), .A3(new_n709), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT115), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(KEYINPUT115), .B(KEYINPUT50), .C1(new_n813), .C2(new_n819), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(KEYINPUT116), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n822), .B2(new_n823), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT51), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n807), .A2(new_n747), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT48), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n809), .A2(new_n621), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n832), .B(new_n469), .C1(new_n710), .C2(new_n813), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n834), .B1(new_n817), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT117), .B1(new_n829), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n838), .ZN(new_n840));
  INV_X1    g654(.A(new_n828), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n835), .B1(new_n841), .B2(new_n817), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n723), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n611), .A2(new_n548), .A3(new_n683), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n687), .A2(new_n732), .A3(new_n657), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n682), .A2(new_n731), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n669), .A2(new_n696), .A3(new_n846), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g664(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n723), .B1(new_n660), .B2(new_n668), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n849), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n704), .A2(new_n707), .A3(new_n712), .A4(new_n718), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n739), .A2(new_n740), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n744), .A2(new_n748), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n859), .A3(KEYINPUT53), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n319), .B1(new_n714), .B2(G472), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n611), .A2(new_n618), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n672), .A2(new_n861), .A3(new_n862), .A4(new_n604), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n377), .B2(new_n601), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n611), .A2(new_n467), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n672), .A2(new_n861), .A3(new_n604), .A4(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n601), .B2(new_n646), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n864), .B1(KEYINPUT109), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT109), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n867), .B(new_n870), .C1(new_n601), .C2(new_n646), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n862), .B1(new_n741), .B2(new_n735), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n645), .B1(new_n745), .B2(new_n680), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n627), .A2(new_n628), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n431), .A2(new_n683), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n782), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n874), .B(new_n876), .C1(new_n599), .C2(new_n600), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n872), .A2(new_n722), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n657), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n377), .A2(new_n742), .ZN(new_n880));
  AOI22_X1  g694(.A1(new_n878), .A2(new_n879), .B1(new_n880), .B2(new_n658), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n869), .A2(new_n871), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n860), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n869), .A2(new_n881), .A3(KEYINPUT112), .A4(new_n871), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n855), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n704), .A2(new_n707), .A3(new_n712), .A4(new_n718), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n749), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n871), .A3(new_n869), .A4(new_n881), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n850), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n854), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n886), .B(new_n887), .C1(new_n893), .C2(KEYINPUT53), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n892), .A2(new_n854), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n605), .A2(new_n865), .A3(new_n609), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT109), .B1(new_n896), .B2(new_n647), .ZN(new_n897));
  INV_X1    g711(.A(new_n601), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n862), .A2(new_n610), .B1(new_n898), .B2(new_n699), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n899), .A3(new_n871), .ZN(new_n900));
  INV_X1    g714(.A(new_n862), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n736), .B2(new_n737), .ZN(new_n902));
  INV_X1    g716(.A(new_n722), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n467), .B1(new_n430), .B2(G475), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n805), .A2(new_n627), .A3(new_n628), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(new_n652), .B2(new_n653), .ZN(new_n906));
  AOI22_X1  g720(.A1(new_n902), .A2(new_n903), .B1(new_n666), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n752), .B1(new_n907), .B2(new_n657), .ZN(new_n908));
  NOR4_X1   g722(.A1(new_n900), .A2(new_n908), .A3(new_n749), .A4(new_n888), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n895), .A2(KEYINPUT53), .A3(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT53), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT110), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n890), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n912), .A2(new_n914), .A3(new_n855), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n910), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n894), .B1(new_n916), .B2(new_n887), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT113), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT113), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n919), .B(new_n894), .C1(new_n916), .C2(new_n887), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n845), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(G952), .A2(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n804), .B1(new_n921), .B2(new_n922), .ZN(G75));
  OAI21_X1  g737(.A(new_n883), .B1(new_n900), .B2(new_n908), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n749), .A2(new_n888), .A3(new_n911), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n924), .A2(new_n885), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n854), .B2(new_n852), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n895), .B2(new_n909), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n312), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(G210), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n541), .A2(new_n542), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n492), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n543), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT119), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n931), .A2(new_n932), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n938), .B1(new_n931), .B2(new_n932), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n246), .A2(G952), .ZN(new_n941));
  NOR3_X1   g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(G51));
  OAI21_X1  g756(.A(new_n886), .B1(new_n893), .B2(KEYINPUT53), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(G902), .A3(new_n774), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n943), .A2(new_n946), .A3(G902), .A4(new_n774), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT54), .B1(new_n927), .B2(new_n928), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n894), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n595), .B(KEYINPUT57), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n700), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n948), .B1(new_n954), .B2(KEYINPUT120), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT120), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n952), .A2(new_n956), .A3(new_n953), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n941), .B1(new_n955), .B2(new_n957), .ZN(G54));
  NAND3_X1  g772(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n418), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n418), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n961), .A3(new_n941), .ZN(G60));
  INV_X1    g776(.A(new_n614), .ZN(new_n963));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n950), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n941), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n918), .A2(new_n920), .A3(new_n965), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n969), .B2(new_n614), .ZN(G63));
  AND2_X1   g784(.A1(new_n637), .A2(new_n638), .ZN(new_n971));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT60), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n971), .B(new_n974), .C1(new_n927), .C2(new_n928), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n967), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n372), .B1(new_n943), .B2(new_n974), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT123), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n372), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n929), .B2(new_n973), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n980), .A2(new_n981), .A3(new_n967), .A4(new_n975), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT61), .B1(new_n975), .B2(KEYINPUT122), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n978), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n978), .B2(new_n982), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G66));
  NOR2_X1   g800(.A1(new_n900), .A2(new_n888), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT124), .Z(new_n988));
  NAND2_X1  g802(.A1(new_n474), .A2(G224), .ZN(new_n989));
  AOI22_X1  g803(.A1(new_n988), .A2(new_n246), .B1(G953), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n933), .B1(G898), .B2(new_n246), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n990), .B(new_n991), .Z(G69));
  AND3_X1   g806(.A1(new_n767), .A2(new_n781), .A3(new_n783), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n748), .A2(new_n847), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n780), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AND2_X1   g809(.A1(new_n853), .A2(new_n696), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n791), .A2(new_n859), .A3(new_n752), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n354), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n232), .B(new_n404), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n656), .B2(new_n246), .ZN(new_n1001));
  OR2_X1    g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n782), .B1(new_n901), .B2(new_n865), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1004), .A2(new_n699), .A3(new_n672), .A4(new_n673), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n784), .A2(new_n791), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n996), .A2(new_n689), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1006), .B1(KEYINPUT62), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1008), .B1(KEYINPUT62), .B2(new_n1007), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n1009), .A2(new_n246), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1000), .B(KEYINPUT125), .Z(new_n1011));
  OAI211_X1 g825(.A(new_n1002), .B(new_n1003), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1003), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1011), .B1(new_n1009), .B2(new_n246), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n999), .A2(new_n1001), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  AND2_X1   g830(.A1(new_n1012), .A2(new_n1016), .ZN(G72));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT126), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n1009), .B2(new_n988), .ZN(new_n1021));
  INV_X1    g835(.A(new_n264), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1021), .A2(new_n260), .A3(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n294), .A2(new_n261), .A3(new_n300), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n1019), .ZN(new_n1025));
  OR2_X1    g839(.A1(new_n916), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1020), .B1(new_n998), .B2(new_n988), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n264), .A2(new_n259), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1028), .B(KEYINPUT127), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n941), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1023), .A2(new_n1026), .A3(new_n1030), .ZN(G57));
endmodule


