//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT1), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n222), .A2(new_n208), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(new_n217), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n217), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT64), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(new_n226), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G226), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT16), .ZN(new_n248));
  INV_X1    g0048(.A(G58), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(new_n242), .ZN(new_n250));
  OAI21_X1  g0050(.A(G20), .B1(new_n250), .B2(new_n201), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G159), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n206), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT7), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n259), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n242), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n255), .B1(new_n264), .B2(KEYINPUT74), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT74), .ZN(new_n266));
  AOI211_X1 g0066(.A(new_n266), .B(new_n242), .C1(new_n262), .C2(new_n263), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n248), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT75), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n270), .B(new_n248), .C1(new_n265), .C2(new_n267), .ZN(new_n271));
  NAND3_X1  g0071(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n214), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n263), .A2(KEYINPUT73), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT73), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(KEYINPUT7), .A4(new_n206), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(new_n280), .A3(new_n262), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n254), .B1(new_n281), .B2(G68), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n274), .B1(new_n282), .B2(KEYINPUT16), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n269), .A2(new_n271), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n205), .B2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n206), .A3(G1), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n273), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n286), .A2(new_n289), .B1(new_n288), .B2(new_n285), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(G1), .A3(G13), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n294), .A3(G274), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G232), .A3(new_n291), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n258), .A2(new_n259), .ZN(new_n298));
  INV_X1    g0098(.A(G1698), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n298), .A2(G223), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(G226), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n301));
  INV_X1    g0101(.A(G87), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n257), .A2(new_n302), .A3(KEYINPUT76), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT76), .B1(new_n257), .B2(new_n302), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(new_n301), .A3(new_n303), .A4(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n294), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n297), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(G200), .B2(new_n307), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT78), .A2(KEYINPUT17), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n284), .A2(new_n290), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n284), .A2(new_n290), .A3(new_n310), .ZN(new_n313));
  XOR2_X1   g0113(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n314));
  OAI21_X1  g0114(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n284), .A2(new_n290), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT77), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n307), .A2(G179), .ZN(new_n318));
  INV_X1    g0118(.A(G169), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n307), .A2(G179), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(KEYINPUT77), .C1(new_n319), .C2(new_n307), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT18), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT18), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n316), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n315), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G226), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n294), .A2(new_n291), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n295), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n299), .B1(new_n258), .B2(new_n259), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n333), .A2(G223), .B1(new_n278), .B2(G77), .ZN(new_n334));
  INV_X1    g0134(.A(G222), .ZN(new_n335));
  AOI21_X1  g0135(.A(G1698), .B1(new_n258), .B2(new_n259), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n332), .B1(new_n338), .B2(new_n306), .ZN(new_n339));
  INV_X1    g0139(.A(G200), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n206), .A2(G33), .ZN(new_n342));
  INV_X1    g0142(.A(G150), .ZN(new_n343));
  INV_X1    g0143(.A(new_n252), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n285), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n206), .B1(new_n201), .B2(new_n240), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n273), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n205), .A2(G20), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G50), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n289), .A2(new_n350), .B1(new_n240), .B2(new_n288), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT9), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n339), .A2(G190), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n341), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT10), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n339), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n352), .B1(new_n339), .B2(G169), .ZN(new_n359));
  OR2_X1    g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n285), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n342), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n273), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n205), .B2(G20), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n289), .A2(new_n368), .B1(new_n367), .B2(new_n288), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G244), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n295), .B1(new_n371), .B2(new_n331), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n333), .A2(G238), .B1(new_n278), .B2(G107), .ZN(new_n373));
  INV_X1    g0173(.A(G232), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n337), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(new_n306), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n370), .B1(new_n376), .B2(new_n340), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n376), .A2(G190), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n366), .A2(new_n369), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n380), .B1(new_n376), .B2(G169), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(KEYINPUT66), .B1(new_n357), .B2(new_n376), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n381), .A2(KEYINPUT66), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n329), .A2(new_n361), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n299), .A2(G226), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT67), .B1(new_n278), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT67), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n298), .A2(new_n391), .A3(G226), .A4(new_n299), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(G232), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n298), .A2(KEYINPUT68), .A3(G232), .A4(G1698), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n393), .A2(KEYINPUT69), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT69), .B1(new_n393), .B2(new_n398), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n399), .A2(new_n400), .A3(new_n294), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT70), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n295), .B(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G238), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT71), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n331), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n405), .B2(new_n331), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT13), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n390), .A2(new_n392), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n398), .A2(new_n410), .A3(new_n387), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT69), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n393), .A2(KEYINPUT69), .A3(new_n398), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n414), .A3(new_n306), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  INV_X1    g0216(.A(new_n408), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n409), .A2(G190), .A3(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n288), .A2(new_n242), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT12), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n242), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n367), .B2(new_n342), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT11), .A3(new_n273), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n289), .A2(G68), .A3(new_n348), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT11), .B1(new_n425), .B2(new_n273), .ZN(new_n429));
  OR2_X1    g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n420), .A2(new_n421), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n294), .B1(new_n411), .B2(new_n412), .ZN(new_n434));
  AOI211_X1 g0234(.A(KEYINPUT13), .B(new_n408), .C1(new_n434), .C2(new_n414), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n433), .B(G169), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT72), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n419), .A2(KEYINPUT72), .A3(new_n433), .A4(G169), .ZN(new_n440));
  OAI21_X1  g0240(.A(G169), .B1(new_n435), .B2(new_n436), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT14), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n409), .A2(G179), .A3(new_n418), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n439), .A2(new_n440), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n432), .B1(new_n444), .B2(new_n430), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n386), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT79), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n386), .A2(KEYINPUT79), .A3(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n206), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n298), .A2(new_n454), .A3(new_n206), .A4(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT24), .ZN(new_n457));
  INV_X1    g0257(.A(G116), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n342), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT84), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n206), .B2(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT23), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT23), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n460), .B(new_n463), .C1(new_n206), .C2(G107), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n459), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n456), .A2(new_n457), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n457), .B1(new_n456), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n273), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT25), .ZN(new_n469));
  INV_X1    g0269(.A(new_n288), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(G107), .ZN(new_n471));
  INV_X1    g0271(.A(G107), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n288), .A2(KEYINPUT25), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n257), .A2(G1), .ZN(new_n474));
  NOR3_X1   g0274(.A1(new_n288), .A2(new_n273), .A3(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n471), .A2(new_n473), .B1(new_n475), .B2(G107), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT87), .ZN(new_n479));
  INV_X1    g0279(.A(G274), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n306), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT5), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G41), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(KEYINPUT81), .A3(new_n205), .A4(G45), .ZN(new_n484));
  INV_X1    g0284(.A(G41), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT5), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n205), .B(G45), .C1(new_n485), .C2(KEYINPUT5), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT81), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n481), .A2(new_n484), .A3(new_n486), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n484), .A3(new_n486), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(G264), .A3(new_n294), .ZN(new_n492));
  OAI211_X1 g0292(.A(G257), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G294), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT85), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n336), .A2(new_n496), .A3(G250), .ZN(new_n497));
  OAI211_X1 g0297(.A(G250), .B(new_n299), .C1(new_n276), .C2(new_n277), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n490), .B(new_n492), .C1(new_n500), .C2(new_n294), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G200), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n493), .A2(new_n494), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n496), .B1(new_n336), .B2(G250), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n498), .A2(KEYINPUT85), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n306), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(G190), .A3(new_n490), .A4(new_n492), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n478), .A2(new_n479), .A3(new_n502), .A4(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n502), .A2(new_n508), .A3(new_n468), .A4(new_n476), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT87), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n501), .A2(G169), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n507), .A2(G179), .A3(new_n490), .A4(new_n492), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT86), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT86), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n516), .A2(new_n477), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n512), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n475), .A2(G97), .ZN(new_n521));
  INV_X1    g0321(.A(G97), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n288), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g0324(.A(G97), .B(G107), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g0327(.A1(new_n526), .A2(new_n522), .A3(G107), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n472), .B1(new_n262), .B2(new_n263), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n524), .B1(new_n534), .B2(new_n273), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(new_n299), .C1(new_n276), .C2(new_n277), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT4), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n298), .A2(KEYINPUT4), .A3(G244), .A4(new_n299), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n298), .A2(G250), .A3(G1698), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n538), .A2(new_n539), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT80), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n333), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT80), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n544), .A2(new_n545), .A3(new_n539), .A4(new_n538), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n306), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n491), .A2(new_n294), .ZN(new_n548));
  INV_X1    g0348(.A(G257), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n490), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n535), .B1(new_n552), .B2(new_n319), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n294), .B1(new_n542), .B2(KEYINPUT80), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n550), .B1(new_n554), .B2(new_n546), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n357), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n528), .B1(new_n526), .B2(new_n525), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n558), .A2(new_n206), .B1(new_n367), .B2(new_n344), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n273), .B1(new_n559), .B2(new_n532), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(new_n523), .A3(new_n521), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n552), .B2(G200), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n555), .A2(G190), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT19), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n206), .B1(new_n387), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n302), .A2(new_n522), .A3(new_n472), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n206), .B(G68), .C1(new_n276), .C2(new_n277), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n565), .B1(new_n342), .B2(new_n522), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n273), .B1(new_n288), .B2(new_n364), .ZN(new_n572));
  INV_X1    g0372(.A(new_n364), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n475), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  INV_X1    g0376(.A(G45), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(G1), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n205), .A2(new_n480), .A3(G45), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n294), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n582));
  OAI211_X1 g0382(.A(G238), .B(new_n299), .C1(new_n276), .C2(new_n277), .ZN(new_n583));
  NAND2_X1  g0383(.A1(G33), .A2(G116), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n581), .B1(new_n585), .B2(new_n306), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(G169), .ZN(new_n587));
  AOI211_X1 g0387(.A(G179), .B(new_n581), .C1(new_n585), .C2(new_n306), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n585), .A2(new_n306), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n340), .B1(new_n590), .B2(new_n580), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n571), .A2(new_n273), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n364), .A2(new_n288), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n475), .A2(G87), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n586), .A2(G190), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n575), .A2(new_n589), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n557), .A2(new_n564), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n540), .B(new_n206), .C1(G33), .C2(new_n522), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n273), .C1(new_n206), .C2(G116), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n601), .B(KEYINPUT20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n475), .A2(G116), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G116), .B2(new_n470), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n491), .A2(G270), .A3(new_n294), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT82), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n491), .A2(KEYINPUT82), .A3(G270), .A4(new_n294), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n609), .A2(new_n490), .A3(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n299), .C1(new_n276), .C2(new_n277), .ZN(new_n613));
  INV_X1    g0413(.A(G303), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n298), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n357), .B1(new_n615), .B2(new_n306), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n606), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n306), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n609), .A2(new_n620), .A3(new_n490), .A4(new_n610), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n610), .A2(new_n490), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n624), .A2(KEYINPUT83), .A3(new_n620), .A4(new_n609), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(G169), .B1(new_n602), .B2(new_n604), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n619), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n626), .A2(new_n619), .A3(new_n628), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n618), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n606), .B1(new_n626), .B2(G200), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n308), .B2(new_n626), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n520), .A2(new_n599), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n451), .A2(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n360), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n318), .A2(new_n320), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n327), .B1(new_n316), .B2(new_n639), .ZN(new_n640));
  AOI211_X1 g0440(.A(KEYINPUT18), .B(new_n638), .C1(new_n284), .C2(new_n290), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n444), .A2(new_n430), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n383), .A2(new_n382), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n432), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n315), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n642), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n637), .B1(new_n648), .B2(new_n356), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n515), .A2(new_n477), .ZN(new_n650));
  AOI211_X1 g0450(.A(KEYINPUT21), .B(new_n627), .C1(new_n623), .C2(new_n625), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n617), .B(new_n650), .C1(new_n629), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n557), .A2(new_n564), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n572), .B(new_n594), .C1(new_n586), .C2(new_n340), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT88), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n655), .A2(new_n656), .B1(G190), .B2(new_n586), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n596), .A2(KEYINPUT88), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n575), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n660), .A2(new_n587), .A3(new_n588), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n509), .B2(new_n511), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n652), .A2(new_n654), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n553), .A2(new_n598), .A3(new_n556), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n661), .B1(new_n666), .B2(KEYINPUT26), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n561), .B1(new_n555), .B2(G169), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n547), .A2(new_n551), .A3(new_n357), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT89), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n552), .A2(new_n319), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT89), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n556), .A3(new_n672), .A4(new_n561), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n661), .B1(new_n657), .B2(new_n658), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n670), .A2(new_n673), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n665), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n649), .B1(new_n451), .B2(new_n678), .ZN(G369));
  INV_X1    g0479(.A(new_n632), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n605), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n632), .A2(new_n634), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n689), .B1(new_n690), .B2(new_n688), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  OAI211_X1 g0492(.A(new_n512), .B(new_n519), .C1(new_n478), .C2(new_n687), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n519), .A2(new_n687), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n693), .A2(KEYINPUT90), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n692), .A2(new_n699), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT91), .Z(new_n701));
  NOR2_X1   g0501(.A1(new_n632), .A2(new_n686), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n650), .A2(new_n686), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n701), .A2(new_n703), .A3(new_n705), .ZN(G399));
  INV_X1    g0506(.A(new_n209), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G41), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n567), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n212), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n492), .B1(new_n500), .B2(new_n294), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n616), .A2(new_n586), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n555), .A3(new_n611), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n716), .A2(new_n555), .A3(KEYINPUT92), .A4(new_n611), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n716), .A2(new_n555), .A3(KEYINPUT30), .A4(new_n611), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n586), .A2(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n626), .A2(new_n501), .A3(new_n552), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n723), .A2(new_n724), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n722), .A2(new_n725), .A3(new_n727), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n686), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n732), .B(new_n733), .C1(new_n635), .C2(new_n686), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT94), .B1(new_n678), .B2(new_n686), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n652), .A2(new_n654), .A3(new_n664), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n667), .A2(new_n676), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n686), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n742));
  NAND3_X1  g0542(.A1(new_n736), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT96), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n519), .B(new_n617), .C1(new_n629), .C2(new_n651), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(new_n654), .A3(new_n664), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n553), .A2(new_n598), .A3(new_n675), .A4(new_n556), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n662), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n748), .B1(KEYINPUT26), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n744), .B1(new_n751), .B2(new_n687), .ZN(new_n752));
  AOI211_X1 g0552(.A(KEYINPUT96), .B(new_n686), .C1(new_n746), .C2(new_n750), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n735), .B1(new_n743), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n713), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n287), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n205), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n708), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n692), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G330), .B2(new_n691), .ZN(new_n762));
  OAI21_X1  g0562(.A(G20), .B1(KEYINPUT98), .B2(G169), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(KEYINPUT98), .B2(G169), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n214), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT99), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(KEYINPUT100), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n707), .A2(new_n298), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n577), .B2(new_n213), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(new_n246), .B2(new_n577), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n209), .A2(new_n298), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT97), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G355), .B1(new_n458), .B2(new_n707), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n775), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n308), .A2(new_n340), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n784), .A2(G20), .A3(new_n357), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT102), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n206), .A2(new_n357), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT101), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(KEYINPUT101), .B1(new_n206), .B2(new_n357), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n308), .A2(G200), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n789), .A2(new_n302), .B1(new_n249), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(G190), .A2(G200), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n792), .A2(new_n793), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(G77), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n206), .A2(G190), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n801), .A2(new_n357), .A3(new_n340), .ZN(new_n802));
  INV_X1    g0602(.A(G159), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT32), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n801), .A2(G179), .A3(G200), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n790), .A2(new_n784), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n298), .B1(new_n806), .B2(new_n242), .C1(new_n240), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n794), .A2(new_n357), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n522), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n801), .A2(new_n357), .A3(G200), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n472), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n808), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n800), .A2(new_n805), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n789), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G303), .B1(G311), .B2(new_n799), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n811), .A2(new_n819), .B1(new_n813), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n802), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(G329), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G326), .ZN(new_n824));
  XOR2_X1   g0624(.A(KEYINPUT33), .B(G317), .Z(new_n825));
  OAI221_X1 g0625(.A(new_n278), .B1(new_n807), .B2(new_n824), .C1(new_n806), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n795), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n826), .B1(G322), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n818), .A2(new_n823), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n769), .B1(new_n816), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n760), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n783), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n691), .B2(new_n773), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n762), .A2(new_n833), .ZN(G396));
  NOR2_X1   g0634(.A1(new_n370), .A2(new_n687), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n384), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n644), .B2(new_n836), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n736), .A2(new_n741), .A3(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n840), .A2(KEYINPUT106), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n838), .B(new_n687), .C1(new_n665), .C2(new_n677), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n840), .A2(KEYINPUT106), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n735), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n760), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n844), .A2(new_n735), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n768), .A2(new_n770), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n760), .B1(new_n850), .B2(G77), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n789), .A2(new_n472), .B1(new_n458), .B2(new_n798), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G294), .B2(new_n827), .ZN(new_n853));
  INV_X1    g0653(.A(G311), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n302), .A2(new_n813), .B1(new_n802), .B2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT103), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n278), .B1(new_n807), .B2(new_n614), .ZN(new_n857));
  INV_X1    g0657(.A(new_n806), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n857), .B(new_n812), .C1(G283), .C2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n853), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n298), .B1(new_n813), .B2(new_n242), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n811), .A2(new_n249), .B1(new_n802), .B2(new_n862), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n817), .C2(G50), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT104), .ZN(new_n865));
  INV_X1    g0665(.A(new_n807), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G137), .A2(new_n866), .B1(new_n858), .B2(G150), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n868), .B2(new_n795), .C1(new_n803), .C2(new_n798), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT34), .Z(new_n870));
  OAI21_X1  g0670(.A(new_n860), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n851), .B1(new_n871), .B2(new_n768), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n838), .B2(new_n771), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT105), .Z(new_n874));
  NOR2_X1   g0674(.A1(new_n848), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(G384));
  OR2_X1    g0676(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n877), .A2(G116), .A3(new_n215), .A4(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  OR3_X1    g0680(.A1(new_n212), .A2(new_n367), .A3(new_n250), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n205), .B(G13), .C1(new_n881), .C2(new_n241), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n684), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n642), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n643), .A2(new_n646), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n430), .A2(new_n686), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT108), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n888), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n445), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n644), .A2(new_n686), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n842), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n842), .A2(KEYINPUT107), .A3(new_n894), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n892), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT7), .B1(new_n278), .B2(new_n206), .ZN(new_n900));
  INV_X1    g0700(.A(new_n263), .ZN(new_n901));
  OAI21_X1  g0701(.A(G68), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n254), .B1(new_n902), .B2(new_n266), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n264), .A2(KEYINPUT74), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT16), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n283), .B1(new_n905), .B2(new_n270), .ZN(new_n906));
  INV_X1    g0706(.A(new_n271), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n290), .B(new_n310), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n282), .A2(KEYINPUT16), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n273), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n282), .A2(KEYINPUT16), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n290), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n639), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT109), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(KEYINPUT109), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n884), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n684), .B1(new_n284), .B2(new_n290), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n313), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT37), .B1(new_n316), .B2(new_n324), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n919), .A2(KEYINPUT37), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n316), .A2(new_n324), .A3(new_n327), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n327), .B1(new_n316), .B2(new_n324), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n918), .B1(new_n927), .B2(new_n315), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n923), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n917), .A2(new_n918), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT109), .B1(new_n908), .B2(new_n913), .ZN(new_n931));
  OAI21_X1  g0731(.A(KEYINPUT37), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n921), .A2(new_n922), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(new_n918), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n329), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT38), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n929), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n885), .B1(new_n899), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n444), .A2(new_n430), .A3(new_n687), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n934), .A2(KEYINPUT38), .A3(new_n936), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT110), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n316), .A2(new_n884), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n642), .B2(new_n315), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n316), .A2(new_n639), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n946), .A3(new_n908), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n949), .A2(KEYINPUT37), .B1(new_n921), .B2(new_n922), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n924), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n943), .A2(new_n945), .A3(new_n951), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(KEYINPUT110), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n924), .B1(new_n923), .B2(new_n928), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n945), .B1(new_n955), .B2(new_n943), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n942), .B(new_n952), .C1(new_n954), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n940), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n450), .A2(new_n754), .A3(new_n743), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n649), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n958), .B(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n889), .A2(new_n734), .A3(new_n838), .A4(new_n891), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n962), .B1(new_n938), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n734), .A2(new_n838), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n445), .B(new_n888), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n943), .A2(new_n951), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(KEYINPUT40), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n450), .A2(new_n734), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(G330), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n961), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n205), .B2(new_n757), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n961), .A2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n883), .B1(new_n975), .B2(new_n976), .ZN(G367));
  OAI21_X1  g0777(.A(new_n654), .B1(new_n535), .B2(new_n687), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n553), .A2(new_n556), .A3(new_n686), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n699), .A2(new_n702), .A3(new_n980), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT42), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n557), .B1(new_n978), .B2(new_n519), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n981), .A2(KEYINPUT42), .B1(new_n687), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n595), .A2(new_n686), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n674), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n662), .B2(new_n985), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n982), .A2(new_n984), .B1(KEYINPUT43), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(KEYINPUT43), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n988), .B(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n701), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n980), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n990), .B(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n708), .B(KEYINPUT41), .Z(new_n994));
  NAND2_X1  g0794(.A1(new_n703), .A2(new_n705), .ZN(new_n995));
  INV_X1    g0795(.A(new_n980), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT111), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT111), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n999), .A3(new_n996), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(KEYINPUT44), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT44), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n999), .B1(new_n995), .B2(new_n996), .ZN(new_n1003));
  AOI211_X1 g0803(.A(KEYINPUT111), .B(new_n980), .C1(new_n703), .C2(new_n705), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n703), .A2(new_n705), .A3(new_n980), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1001), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n991), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n699), .A2(new_n702), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1011), .A2(new_n703), .A3(new_n692), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n692), .B1(new_n1011), .B2(new_n703), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n755), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n701), .A2(new_n1001), .A3(new_n1005), .A4(new_n1008), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1010), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n994), .B1(new_n1019), .B2(new_n755), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n993), .B1(new_n1020), .B2(new_n759), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n777), .A2(new_n235), .B1(new_n209), .B2(new_n364), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n760), .B1(new_n774), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1024));
  AOI21_X1  g0824(.A(KEYINPUT46), .B1(new_n817), .B2(G116), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n811), .A2(new_n472), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(KEYINPUT112), .B(G317), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n522), .A2(new_n813), .B1(new_n802), .B2(new_n1027), .ZN(new_n1028));
  NOR4_X1   g0828(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n298), .B1(new_n866), .B2(G311), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n819), .B2(new_n806), .C1(new_n614), .C2(new_n795), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G283), .B2(new_n799), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n298), .B1(new_n806), .B2(new_n803), .C1(new_n868), .C2(new_n807), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n789), .A2(new_n249), .B1(new_n343), .B2(new_n795), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G50), .C2(new_n799), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n813), .A2(new_n367), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n811), .A2(new_n242), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G137), .C2(new_n822), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1029), .A2(new_n1032), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT47), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n769), .B1(new_n1039), .B2(KEYINPUT47), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1023), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n773), .B2(new_n987), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1021), .A2(new_n1043), .ZN(G387));
  NOR2_X1   g0844(.A1(new_n1017), .A2(new_n709), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G322), .A2(new_n866), .B1(new_n858), .B2(G311), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n614), .B2(new_n798), .C1(new_n795), .C2(new_n1027), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT48), .ZN(new_n1050));
  OR2_X1    g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n817), .A2(G294), .B1(G283), .B2(new_n810), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT49), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n278), .B1(new_n802), .B2(new_n824), .C1(new_n458), .C2(new_n813), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n278), .B1(new_n858), .B2(new_n362), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n242), .B2(new_n798), .C1(new_n803), .C2(new_n807), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n789), .A2(new_n367), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n810), .A2(new_n573), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n522), .B2(new_n813), .C1(new_n343), .C2(new_n802), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n795), .A2(new_n240), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n768), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n775), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n710), .ZN(new_n1067));
  AOI211_X1 g0867(.A(G45), .B(new_n1067), .C1(G68), .C2(G77), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n285), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n777), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n232), .B2(new_n577), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n781), .A2(new_n1067), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G107), .C2(new_n209), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n831), .B1(new_n1066), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1065), .B(new_n1075), .C1(new_n699), .C2(new_n773), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(new_n1014), .B2(new_n759), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1047), .A2(new_n1078), .ZN(G393));
  NAND3_X1  g0879(.A1(new_n1010), .A2(new_n759), .A3(new_n1018), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n777), .A2(new_n239), .B1(new_n522), .B2(new_n209), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n760), .B1(new_n774), .B2(new_n1081), .ZN(new_n1082));
  XNOR2_X1  g0882(.A(new_n1082), .B(KEYINPUT113), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n827), .A2(G311), .B1(G317), .B2(new_n866), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT52), .Z(new_n1085));
  AOI211_X1 g0885(.A(new_n298), .B(new_n814), .C1(G303), .C2(new_n858), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G322), .A2(new_n822), .B1(new_n810), .B2(G116), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n817), .A2(G283), .B1(G294), .B2(new_n799), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n811), .A2(new_n367), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n298), .B1(new_n806), .B2(new_n240), .C1(new_n302), .C2(new_n813), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n1090), .B(new_n1091), .C1(G143), .C2(new_n822), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n795), .A2(new_n803), .B1(new_n343), .B2(new_n807), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n817), .A2(G68), .B1(new_n362), .B2(new_n799), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1092), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1089), .A2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1083), .B1(new_n769), .B2(new_n1097), .C1(new_n980), .C2(new_n773), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1019), .A2(new_n708), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1017), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1080), .B(new_n1098), .C1(new_n1099), .C2(new_n1100), .ZN(G390));
  OAI21_X1  g0901(.A(KEYINPUT39), .B1(new_n929), .B2(new_n937), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(KEYINPUT110), .A3(new_n953), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n896), .B(new_n893), .C1(new_n739), .C2(new_n838), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT107), .B1(new_n842), .B2(new_n894), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n966), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1103), .A2(new_n952), .B1(new_n941), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n735), .A2(new_n966), .A3(new_n838), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n838), .B1(new_n752), .B2(new_n753), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n892), .B1(new_n1109), .B2(new_n894), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n967), .A2(new_n941), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1108), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT114), .B1(new_n1107), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n952), .B1(new_n954), .B2(new_n956), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1106), .A2(new_n941), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n734), .A2(G330), .A3(new_n838), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n892), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n751), .A2(new_n687), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT96), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n751), .A2(new_n744), .A3(new_n687), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n839), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n966), .B1(new_n1122), .B2(new_n893), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1111), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1118), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1116), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1113), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1118), .B1(new_n1107), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n450), .A2(new_n735), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n959), .A2(new_n649), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AND2_X1   g0935(.A1(new_n892), .A2(new_n1117), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1136), .A2(new_n1118), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n892), .A2(new_n1117), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1108), .A2(new_n894), .A3(new_n1138), .A4(new_n1109), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1135), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1132), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1134), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1116), .A2(new_n1126), .A3(new_n1125), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1126), .B1(new_n1116), .B2(new_n1125), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1143), .B(new_n1131), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1142), .A2(new_n708), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT118), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT117), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1114), .A2(new_n770), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1090), .ZN(new_n1151));
  OAI221_X1 g0951(.A(new_n1151), .B1(new_n242), .B2(new_n813), .C1(new_n819), .C2(new_n802), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n298), .B1(new_n866), .B2(G283), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n472), .B2(new_n806), .C1(new_n789), .C2(new_n302), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n522), .A2(new_n798), .B1(new_n795), .B2(new_n458), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1152), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G128), .A2(new_n866), .B1(new_n858), .B2(G137), .ZN(new_n1157));
  INV_X1    g0957(.A(G125), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n802), .C1(new_n803), .C2(new_n811), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n862), .A2(new_n795), .B1(new_n798), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n298), .B1(new_n813), .B2(new_n240), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT115), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1159), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n789), .A2(new_n343), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1156), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n760), .B1(new_n362), .B2(new_n850), .C1(new_n1167), .C2(new_n769), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT116), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n1150), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n758), .B1(new_n1172), .B2(new_n1118), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1149), .B(new_n1171), .C1(new_n1128), .C2(new_n1173), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n759), .B(new_n1131), .C1(new_n1144), .C2(new_n1145), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT117), .B1(new_n1175), .B2(new_n1170), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1148), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1114), .A2(new_n1115), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n759), .B1(new_n1178), .B2(new_n1108), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n1127), .B2(new_n1113), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1149), .B1(new_n1180), .B2(new_n1171), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1175), .A2(KEYINPUT117), .A3(new_n1170), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(KEYINPUT118), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1147), .B1(new_n1177), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(G378));
  INV_X1    g0985(.A(KEYINPUT121), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n964), .A2(new_n1186), .A3(G330), .A4(new_n968), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n958), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n684), .B1(new_n347), .B2(new_n351), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n361), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n361), .A2(new_n1192), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1191), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n1193), .A3(new_n1190), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n964), .A2(G330), .A3(new_n968), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n1200), .B2(KEYINPUT121), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1187), .A2(new_n957), .A3(new_n940), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1189), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1201), .B1(new_n1189), .B2(new_n1202), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1199), .A2(new_n770), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n760), .B1(new_n850), .B2(G50), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n298), .A2(G41), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(G33), .A2(G41), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1208), .A2(G50), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n813), .A2(new_n249), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1037), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n820), .B2(new_n802), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n472), .A2(new_n795), .B1(new_n798), .B2(new_n364), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1208), .B1(new_n522), .B2(new_n806), .C1(new_n458), .C2(new_n807), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1213), .A2(new_n1060), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  XOR2_X1   g1016(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1210), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n807), .A2(new_n1158), .B1(new_n806), .B2(new_n862), .ZN(new_n1220));
  INV_X1    g1020(.A(G128), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n795), .A2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(G150), .C2(new_n810), .ZN(new_n1223));
  INV_X1    g1023(.A(G137), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1223), .B1(new_n1224), .B2(new_n798), .C1(new_n789), .C2(new_n1160), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1209), .B1(new_n813), .B2(new_n803), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G124), .B2(new_n822), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT120), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1219), .B1(new_n1218), .B2(new_n1216), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1207), .B1(new_n1232), .B2(new_n768), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(new_n1205), .A2(new_n759), .B1(new_n1206), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1201), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1202), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1187), .B1(new_n957), .B2(new_n940), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1189), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(KEYINPUT57), .A3(new_n1239), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1113), .A2(new_n1127), .B1(new_n1118), .B2(new_n1172), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1134), .B1(new_n1241), .B2(new_n1140), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n708), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1146), .A2(new_n1135), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT57), .B1(new_n1205), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1234), .B1(new_n1243), .B2(new_n1245), .ZN(G375));
  NAND3_X1  g1046(.A1(new_n1134), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n994), .B(KEYINPUT122), .Z(new_n1248));
  NAND3_X1  g1048(.A1(new_n1141), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1140), .A2(new_n759), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n831), .B1(new_n849), .B2(new_n242), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n866), .A2(G132), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1252), .B1(new_n806), .B2(new_n1160), .C1(new_n1224), .C2(new_n795), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT124), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n789), .A2(new_n803), .B1(new_n343), .B2(new_n798), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n811), .A2(new_n240), .B1(new_n802), .B2(new_n1221), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(new_n1255), .A2(new_n278), .A3(new_n1211), .A4(new_n1256), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n789), .A2(new_n522), .B1(new_n472), .B2(new_n798), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n278), .B1(new_n806), .B2(new_n458), .C1(new_n819), .C2(new_n807), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n802), .A2(new_n614), .ZN(new_n1260));
  NOR4_X1   g1060(.A1(new_n1258), .A2(new_n1036), .A3(new_n1259), .A4(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1061), .B1(new_n820), .B2(new_n795), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT123), .Z(new_n1263));
  AOI22_X1  g1063(.A1(new_n1254), .A2(new_n1257), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1251), .B1(new_n769), .B2(new_n1264), .C1(new_n966), .C2(new_n771), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1249), .A2(new_n1250), .A3(new_n1265), .ZN(G381));
  INV_X1    g1066(.A(G396), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1047), .A2(new_n1267), .A3(new_n1078), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1269), .A2(G387), .ZN(new_n1270));
  INV_X1    g1070(.A(G375), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1142), .A2(new_n708), .A3(new_n1146), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1270), .A2(new_n1271), .A3(new_n1274), .ZN(G407));
  NAND2_X1  g1075(.A1(new_n685), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1271), .A2(new_n1274), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(G213), .A3(new_n1278), .ZN(G409));
  AND3_X1   g1079(.A1(new_n1205), .A2(new_n1244), .A3(new_n1248), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1206), .A2(new_n1233), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n758), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1273), .B(new_n1272), .C1(new_n1280), .C2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1184), .B2(G375), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n708), .B1(new_n1286), .B2(new_n1247), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1247), .B2(new_n1286), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1250), .A2(new_n1265), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n875), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1141), .A2(KEYINPUT60), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1247), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n709), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1286), .A2(new_n1247), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1289), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(G384), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1290), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1285), .A2(new_n1276), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1285), .A2(KEYINPUT63), .A3(new_n1297), .A4(new_n1276), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1268), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1267), .B1(new_n1047), .B2(new_n1078), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1021), .A2(new_n1043), .A3(G390), .ZN(new_n1307));
  AOI21_X1  g1107(.A(G390), .B1(new_n1021), .B2(new_n1043), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1306), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G390), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(G387), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1305), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1312), .A2(KEYINPUT125), .A3(new_n1268), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1306), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1021), .A2(new_n1043), .A3(G390), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n1314), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1302), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1277), .A2(G2897), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1290), .B2(new_n1296), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1290), .A2(new_n1296), .A3(new_n1319), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1320), .B(new_n1321), .C1(new_n1285), .C2(new_n1276), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT126), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1309), .A2(new_n1316), .A3(new_n1323), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1322), .A2(new_n1324), .A3(KEYINPUT61), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1318), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1317), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1285), .A2(new_n1276), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1321), .A2(new_n1320), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  AOI21_X1  g1131(.A(KEYINPUT126), .B1(new_n1330), .B2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1298), .A2(KEYINPUT62), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT62), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1285), .A2(new_n1334), .A3(new_n1297), .A4(new_n1276), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1333), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1327), .B1(new_n1332), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1326), .A2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1274), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1184), .B2(G375), .ZN(new_n1340));
  OR2_X1    g1140(.A1(new_n1340), .A2(new_n1297), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1297), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  XNOR2_X1  g1143(.A(new_n1343), .B(new_n1327), .ZN(G402));
endmodule


