//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(KEYINPUT67), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT64), .B(G238), .ZN(new_n209));
  AOI22_X1  g0009(.A1(new_n209), .A2(G68), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G77), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  NAND2_X1  g0016(.A1(G107), .A2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G58), .A2(G232), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n208), .B1(new_n221), .B2(new_n203), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n222), .B(new_n223), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n224), .C1(new_n227), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n235), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n225), .ZN(new_n250));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G68), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n253), .B(KEYINPUT74), .Z(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n256), .A2(new_n211), .B1(new_n226), .B2(G68), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n226), .A2(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n213), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n250), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT11), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G68), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT12), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n254), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT68), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT68), .A2(G41), .ZN(new_n270));
  AOI21_X1  g0070(.A(G45), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G1), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(G33), .A2(G97), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n237), .A2(G1698), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G226), .B2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n276), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G1), .A3(G13), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n275), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G238), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n288), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n288), .B(new_n295), .C1(new_n289), .C2(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n268), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n297), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(G179), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT76), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(KEYINPUT75), .B2(KEYINPUT14), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n297), .A2(G169), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(KEYINPUT14), .ZN(new_n308));
  AND3_X1   g0108(.A1(new_n297), .A2(G169), .A3(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n304), .B(new_n307), .C1(new_n309), .C2(new_n306), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n303), .B1(new_n310), .B2(new_n267), .ZN(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT3), .B(G33), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G222), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G223), .A2(G1698), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n287), .C1(G77), .C2(new_n312), .ZN(new_n317));
  INV_X1    g0117(.A(new_n275), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(new_n212), .C2(new_n292), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n319), .A2(G179), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n319), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n252), .A2(G50), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n263), .A2(new_n211), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n229), .B2(G50), .ZN(new_n325));
  INV_X1    g0125(.A(G150), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(new_n256), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT70), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT69), .B(G58), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT8), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G58), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT69), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G58), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT70), .A3(KEYINPUT8), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n330), .A2(KEYINPUT71), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n330), .A2(KEYINPUT71), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n338), .A2(G58), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n258), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n327), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n250), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n323), .B(new_n324), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n322), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n319), .A2(new_n298), .ZN(new_n347));
  OR2_X1    g0147(.A1(new_n345), .A2(KEYINPUT9), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(KEYINPUT9), .ZN(new_n349));
  AOI211_X1 g0149(.A(KEYINPUT73), .B(new_n347), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n319), .A2(G200), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(KEYINPUT10), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT10), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n350), .B2(new_n351), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n311), .B(new_n346), .C1(new_n353), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT17), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT78), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n333), .A2(new_n335), .A3(G68), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n226), .B1(new_n359), .B2(new_n229), .ZN(new_n360));
  INV_X1    g0160(.A(G159), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n256), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n358), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT7), .B1(new_n283), .B2(new_n226), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  AOI211_X1 g0165(.A(new_n365), .B(G20), .C1(new_n280), .C2(new_n282), .ZN(new_n366));
  OAI21_X1  g0166(.A(G68), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n362), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n228), .B1(new_n329), .B2(G68), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT78), .B(new_n368), .C1(new_n369), .C2(new_n226), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT16), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n365), .B1(new_n312), .B2(G20), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n281), .A2(G33), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n376));
  OAI211_X1 g0176(.A(KEYINPUT7), .B(new_n226), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n374), .A2(KEYINPUT77), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT77), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n366), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(G68), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n363), .A4(new_n370), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n373), .A2(new_n250), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n341), .A2(new_n252), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n262), .B2(new_n341), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n212), .A2(G1698), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n280), .A2(new_n387), .A3(new_n282), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n287), .ZN(new_n392));
  INV_X1    g0192(.A(G45), .ZN(new_n393));
  INV_X1    g0193(.A(new_n270), .ZN(new_n394));
  NOR2_X1   g0194(.A1(KEYINPUT68), .A2(G41), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n291), .A2(G232), .B1(new_n396), .B2(new_n273), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT79), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n392), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n286), .B1(new_n389), .B2(new_n390), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n286), .A2(G232), .A3(new_n290), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n271), .B2(new_n274), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT79), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(G200), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n400), .A2(new_n402), .A3(G190), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n386), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n357), .B1(new_n383), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n398), .B1(new_n392), .B2(new_n397), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT79), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n301), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n405), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n385), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n373), .A2(new_n382), .A3(new_n250), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(KEYINPUT17), .A3(new_n413), .ZN(new_n414));
  AND3_X1   g0214(.A1(new_n407), .A2(KEYINPUT80), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT80), .B1(new_n407), .B2(new_n414), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n209), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n418), .B(new_n312), .C1(new_n237), .C2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n287), .C1(G107), .C2(new_n312), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n291), .A2(G244), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n318), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n422), .A2(new_n298), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(G200), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT8), .B(G58), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n256), .B1(new_n226), .B2(new_n213), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n258), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n250), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n252), .A2(G77), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n263), .A2(new_n213), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n423), .B(new_n424), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n422), .A2(new_n321), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n433), .C1(G179), .C2(new_n422), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n413), .A2(new_n386), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n400), .A2(new_n402), .A3(G179), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n399), .A2(new_n403), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(new_n321), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n440), .A2(new_n446), .A3(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n417), .A2(new_n439), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n356), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n279), .A2(G1), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n263), .A2(new_n250), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G107), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n456), .A2(KEYINPUT86), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n226), .B2(G107), .ZN(new_n458));
  INV_X1    g0258(.A(G116), .ZN(new_n459));
  INV_X1    g0259(.A(G107), .ZN(new_n460));
  AOI22_X1  g0260(.A1(KEYINPUT86), .A2(new_n456), .B1(new_n460), .B2(G20), .ZN(new_n461));
  OAI221_X1 g0261(.A(new_n458), .B1(new_n459), .B2(new_n258), .C1(new_n461), .C2(new_n457), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n280), .A2(new_n282), .A3(new_n226), .A4(G87), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT85), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT85), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n312), .A2(new_n466), .A3(new_n226), .A4(G87), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT22), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT24), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g0273(.A(KEYINPUT24), .B(new_n463), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n250), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G41), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT5), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n393), .A2(G1), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT68), .B(G41), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n477), .B(new_n478), .C1(new_n479), .C2(KEYINPUT5), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n480), .A2(new_n286), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G264), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n312), .B1(G257), .B2(new_n313), .ZN(new_n483));
  NOR2_X1   g0283(.A1(G250), .A2(G1698), .ZN(new_n484));
  INV_X1    g0284(.A(G294), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n483), .A2(new_n484), .B1(new_n279), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n287), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n480), .A2(new_n272), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(G190), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n262), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT25), .ZN(new_n492));
  AND4_X1   g0292(.A1(new_n455), .A2(new_n475), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n482), .A2(new_n489), .A3(new_n487), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G200), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n475), .A2(new_n455), .A3(new_n492), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n494), .A2(new_n321), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(G179), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n493), .A2(new_n495), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n280), .A2(new_n282), .A3(G244), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n502), .A2(G1698), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n312), .A2(G244), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G33), .A2(G283), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n312), .A2(G250), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n313), .B1(new_n508), .B2(KEYINPUT4), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n287), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n480), .A2(G257), .A3(new_n286), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n489), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(G169), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n510), .A2(G179), .A3(new_n489), .A4(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(G107), .B1(new_n364), .B2(new_n366), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n460), .A2(KEYINPUT6), .A3(G97), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n518), .A2(new_n460), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n517), .B1(new_n521), .B2(KEYINPUT6), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G20), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n255), .A2(G77), .ZN(new_n524));
  XOR2_X1   g0324(.A(new_n524), .B(KEYINPUT81), .Z(new_n525));
  NAND3_X1  g0325(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n250), .B1(new_n518), .B2(new_n263), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n454), .A2(G97), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n515), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n501), .A2(new_n502), .B1(G33), .B2(G283), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n502), .B1(new_n312), .B2(G250), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n505), .C1(new_n313), .C2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(new_n287), .B1(new_n481), .B2(G257), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(G190), .A3(new_n489), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n512), .A2(G200), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n527), .A4(new_n528), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT82), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n393), .B2(G1), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n251), .A2(new_n272), .A3(G45), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n286), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n289), .A2(new_n313), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n214), .A2(G1698), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n312), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n543), .B1(new_n548), .B2(new_n287), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n538), .B1(new_n549), .B2(G190), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n286), .B1(new_n546), .B2(new_n547), .ZN(new_n551));
  NOR4_X1   g0351(.A1(new_n551), .A2(KEYINPUT82), .A3(new_n298), .A4(new_n543), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G200), .B1(new_n551), .B2(new_n543), .ZN(new_n554));
  INV_X1    g0354(.A(G87), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n520), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n276), .A2(new_n226), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(KEYINPUT19), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n280), .A2(new_n282), .A3(new_n226), .A4(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n276), .B2(G20), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n250), .B1(new_n263), .B2(new_n427), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n454), .A2(G87), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n554), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n548), .A2(new_n287), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n542), .ZN(new_n567));
  INV_X1    g0367(.A(new_n427), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n454), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n567), .A2(new_n321), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G179), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n549), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n553), .A2(new_n565), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n530), .A2(new_n537), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT83), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT83), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n530), .A2(new_n537), .A3(new_n573), .A4(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G264), .A2(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n313), .A2(G257), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n312), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n580), .B(new_n287), .C1(G303), .C2(new_n312), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n480), .A2(G270), .A3(new_n286), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n489), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n506), .B(new_n226), .C1(G33), .C2(new_n518), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n459), .A2(G20), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n250), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT20), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n588), .A2(KEYINPUT84), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n454), .A2(G116), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n586), .A2(new_n592), .A3(new_n587), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n263), .A2(new_n459), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n583), .B(G169), .C1(new_n590), .C2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n583), .A2(new_n571), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n588), .A2(KEYINPUT84), .A3(new_n589), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n600), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n601), .A2(KEYINPUT21), .A3(G169), .A4(new_n583), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n601), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n583), .A2(new_n298), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(G200), .B2(new_n583), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n604), .B1(new_n605), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n500), .A2(new_n575), .A3(new_n577), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n452), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT87), .ZN(G372));
  INV_X1    g0411(.A(new_n346), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n310), .A2(new_n267), .ZN(new_n613));
  XOR2_X1   g0413(.A(new_n438), .B(KEYINPUT89), .Z(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(new_n303), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n417), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n449), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n352), .B(KEYINPUT10), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT82), .B1(new_n567), .B2(new_n298), .ZN(new_n620));
  INV_X1    g0420(.A(new_n552), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n565), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n570), .A2(new_n572), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT26), .B1(new_n530), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n623), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n321), .B1(new_n534), .B2(new_n489), .ZN(new_n628));
  INV_X1    g0428(.A(new_n514), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT88), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n513), .A2(new_n631), .A3(new_n514), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n630), .A2(new_n573), .A3(new_n529), .A4(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n493), .A2(new_n495), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n530), .A2(new_n537), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n573), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n496), .A2(new_n499), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n598), .A2(new_n602), .A3(new_n603), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n627), .B(new_n634), .C1(new_n637), .C2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n619), .B1(new_n452), .B2(new_n643), .ZN(G369));
  INV_X1    g0444(.A(G13), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G20), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n251), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n605), .A2(new_n653), .ZN(new_n654));
  MUX2_X1   g0454(.A(new_n608), .B(new_n604), .S(new_n654), .Z(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n638), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n496), .A2(new_n652), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n657), .B1(new_n635), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n657), .B2(new_n653), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n604), .A2(new_n653), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n500), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n657), .B2(new_n653), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n479), .ZN(new_n669));
  INV_X1    g0469(.A(new_n204), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n520), .A2(new_n555), .A3(new_n459), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n230), .B2(new_n672), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n583), .A2(new_n571), .A3(new_n567), .ZN(new_n678));
  INV_X1    g0478(.A(new_n512), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(new_n488), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT30), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT30), .A4(new_n488), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n583), .A2(new_n571), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n512), .A3(new_n567), .A4(new_n494), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n652), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT31), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n689), .B(new_n690), .C1(new_n609), .C2(new_n652), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n691), .A2(G330), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n642), .A2(new_n653), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n640), .A2(KEYINPUT91), .ZN(new_n696));
  INV_X1    g0496(.A(new_n495), .ZN(new_n697));
  INV_X1    g0497(.A(new_n490), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n496), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n699), .A2(new_n574), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT91), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n638), .A2(new_n639), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT26), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n573), .A2(new_n705), .A3(new_n515), .A4(new_n529), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT90), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n623), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n704), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n572), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n703), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .A3(new_n653), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n692), .B1(new_n695), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n677), .B1(new_n713), .B2(G1), .ZN(G364));
  NAND2_X1  g0514(.A1(new_n646), .A2(G45), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n672), .A2(G1), .A3(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n656), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(G330), .B2(new_n655), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  XOR2_X1   g0520(.A(new_n720), .B(KEYINPUT92), .Z(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT95), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n655), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n571), .A2(new_n301), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n226), .A2(G190), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(G179), .A2(G200), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G159), .ZN(new_n733));
  OAI221_X1 g0533(.A(new_n312), .B1(new_n264), .B2(new_n729), .C1(new_n733), .C2(KEYINPUT32), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(KEYINPUT32), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n226), .A2(new_n298), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n301), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n226), .B1(new_n730), .B2(G190), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n738), .A2(new_n555), .B1(new_n739), .B2(new_n518), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n571), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n737), .A2(new_n728), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n742), .A2(new_n336), .B1(new_n743), .B2(new_n460), .ZN(new_n744));
  NOR4_X1   g0544(.A1(new_n734), .A2(new_n735), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n736), .A2(new_n727), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n728), .A2(new_n741), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n745), .B1(new_n211), .B2(new_n746), .C1(new_n213), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n738), .B(KEYINPUT93), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n283), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT94), .ZN(new_n752));
  INV_X1    g0552(.A(new_n742), .ZN(new_n753));
  AOI22_X1  g0553(.A1(G322), .A2(new_n753), .B1(new_n732), .B2(G329), .ZN(new_n754));
  INV_X1    g0554(.A(G311), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT33), .B(G317), .Z(new_n756));
  OAI221_X1 g0556(.A(new_n754), .B1(new_n755), .B2(new_n747), .C1(new_n729), .C2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n746), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n757), .B1(G326), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n752), .B(new_n759), .C1(new_n485), .C2(new_n739), .ZN(new_n760));
  INV_X1    g0560(.A(G283), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n743), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n748), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n225), .B1(G20), .B2(new_n321), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n231), .A2(new_n393), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n670), .A2(new_n312), .ZN(new_n767));
  OAI211_X1 g0567(.A(new_n766), .B(new_n767), .C1(new_n244), .C2(new_n393), .ZN(new_n768));
  INV_X1    g0568(.A(G355), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n312), .A2(new_n204), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n768), .B1(G116), .B2(new_n204), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n723), .A2(new_n764), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n726), .A2(new_n765), .A3(new_n773), .A4(new_n717), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n719), .A2(new_n774), .ZN(G396));
  AOI21_X1  g0575(.A(new_n626), .B1(new_n700), .B2(new_n640), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n652), .B1(new_n776), .B2(new_n634), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n433), .A2(new_n652), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n439), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n614), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g0581(.A(KEYINPUT97), .B1(new_n777), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n692), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n777), .A2(new_n781), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n783), .B(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(new_n716), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n781), .A2(new_n722), .ZN(new_n787));
  INV_X1    g0587(.A(new_n764), .ZN(new_n788));
  INV_X1    g0588(.A(new_n747), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G143), .A2(new_n753), .B1(new_n789), .B2(G159), .ZN(new_n790));
  INV_X1    g0590(.A(G137), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n790), .B1(new_n791), .B2(new_n746), .C1(new_n326), .C2(new_n729), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT96), .Z(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n739), .A2(new_n336), .ZN(new_n795));
  INV_X1    g0595(.A(new_n743), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G68), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n312), .C1(new_n798), .C2(new_n731), .ZN(new_n799));
  INV_X1    g0599(.A(new_n749), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n795), .B(new_n799), .C1(G50), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n794), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n739), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n800), .A2(G107), .B1(G97), .B2(new_n804), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n805), .B1(new_n555), .B2(new_n743), .C1(new_n755), .C2(new_n731), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n746), .A2(new_n750), .B1(new_n747), .B2(new_n459), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n806), .A2(new_n312), .A3(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n808), .B1(new_n761), .B2(new_n729), .C1(new_n485), .C2(new_n742), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n788), .B1(new_n803), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n764), .A2(new_n720), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G77), .ZN(new_n813));
  NOR4_X1   g0613(.A1(new_n787), .A2(new_n810), .A3(new_n716), .A4(new_n813), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n786), .A2(new_n814), .ZN(G384));
  INV_X1    g0615(.A(KEYINPUT38), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n381), .A2(new_n363), .A3(new_n370), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n344), .B1(new_n817), .B2(new_n372), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT101), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n382), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n818), .A2(new_n819), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n386), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n650), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(new_n417), .B2(new_n449), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n440), .A2(new_n824), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n412), .A2(new_n413), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n444), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n822), .ZN(new_n832));
  INV_X1    g0632(.A(new_n382), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n818), .B2(new_n819), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n385), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n443), .A2(new_n824), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n829), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n831), .B1(new_n837), .B2(KEYINPUT37), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n816), .B1(new_n826), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT80), .ZN(new_n840));
  NOR3_X1   g0640(.A1(new_n383), .A2(new_n406), .A3(new_n357), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT17), .B1(new_n412), .B2(new_n413), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n407), .A2(KEYINPUT80), .A3(new_n414), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n843), .A2(new_n445), .A3(new_n447), .A4(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n824), .A3(new_n823), .ZN(new_n846));
  INV_X1    g0646(.A(new_n836), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n823), .A2(new_n847), .B1(new_n413), .B2(new_n412), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n830), .B1(new_n848), .B2(new_n828), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n846), .A2(new_n849), .A3(KEYINPUT38), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n839), .A2(KEYINPUT102), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n438), .A2(new_n652), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n781), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n693), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n267), .A2(new_n652), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n311), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n310), .A2(new_n267), .A3(new_n652), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT102), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n846), .A2(new_n849), .A3(new_n860), .A4(KEYINPUT38), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n851), .A2(new_n855), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n449), .B2(new_n824), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n613), .A2(new_n652), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n851), .A2(KEYINPUT39), .A3(new_n861), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n444), .A2(new_n827), .A3(new_n829), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT103), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n830), .ZN(new_n870));
  OR3_X1    g0670(.A1(new_n867), .A2(new_n869), .A3(KEYINPUT37), .ZN(new_n871));
  AND4_X1   g0671(.A1(new_n445), .A2(new_n447), .A3(new_n407), .A4(new_n414), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(new_n871), .C1(new_n827), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n816), .ZN(new_n874));
  XNOR2_X1  g0674(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n850), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n865), .B1(new_n866), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n863), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT106), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n695), .A2(new_n712), .A3(new_n451), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n619), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n879), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n451), .A2(new_n691), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT105), .Z(new_n884));
  AND3_X1   g0684(.A1(new_n691), .A2(new_n859), .A3(new_n781), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n851), .A2(new_n885), .A3(new_n861), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT40), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n874), .B2(new_n850), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n886), .A2(new_n887), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n884), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(G330), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n882), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n251), .B2(new_n646), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n231), .A2(G77), .A3(new_n359), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT99), .Z(new_n895));
  NAND2_X1  g0695(.A1(new_n211), .A2(G68), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT100), .ZN(new_n897));
  OAI211_X1 g0697(.A(G1), .B(new_n645), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n459), .B1(new_n522), .B2(KEYINPUT35), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n899), .B(new_n227), .C1(KEYINPUT35), .C2(new_n522), .ZN(new_n900));
  XOR2_X1   g0700(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n901));
  XNOR2_X1  g0701(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n893), .A2(new_n898), .A3(new_n902), .ZN(G367));
  NAND4_X1  g0703(.A1(new_n630), .A2(new_n529), .A3(new_n632), .A4(new_n652), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT107), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n529), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n636), .B1(new_n907), .B2(new_n653), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n905), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n661), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT108), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n563), .A2(new_n564), .ZN(new_n913));
  OR3_X1    g0713(.A1(new_n623), .A2(new_n913), .A3(new_n653), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n653), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n914), .B1(new_n624), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n912), .B(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n666), .A2(new_n910), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT42), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n910), .A2(new_n657), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n652), .B1(new_n922), .B2(new_n530), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n919), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n918), .B(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n671), .B(KEYINPUT41), .Z(new_n926));
  NOR2_X1   g0726(.A1(new_n667), .A2(new_n910), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT44), .Z(new_n928));
  NAND2_X1  g0728(.A1(new_n667), .A2(new_n910), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT45), .ZN(new_n930));
  OR3_X1    g0730(.A1(new_n928), .A2(new_n661), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n661), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  OAI211_X1 g0732(.A(KEYINPUT109), .B(new_n665), .C1(new_n660), .C2(new_n664), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT109), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n656), .B1(new_n934), .B2(new_n666), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n933), .A2(new_n935), .B1(new_n661), .B2(KEYINPUT109), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n713), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n932), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n926), .B1(new_n939), .B2(new_n713), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n715), .A2(G1), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n925), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n767), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n772), .B1(new_n204), .B2(new_n427), .C1(new_n235), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n717), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT110), .ZN(new_n946));
  XNOR2_X1  g0746(.A(KEYINPUT111), .B(G317), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n731), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT46), .B1(new_n749), .B2(new_n459), .ZN(new_n949));
  OR3_X1    g0749(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n459), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n283), .B1(new_n742), .B2(new_n750), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G311), .B2(new_n758), .ZN(new_n953));
  INV_X1    g0753(.A(new_n729), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n954), .A2(G294), .B1(new_n796), .B2(G97), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n804), .A2(G107), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n951), .A2(new_n953), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n948), .B(new_n957), .C1(G283), .C2(new_n789), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n743), .A2(new_n213), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n739), .A2(new_n264), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G143), .B2(new_n758), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n791), .B2(new_n731), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G159), .B2(new_n954), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n326), .B2(new_n742), .C1(new_n336), .C2(new_n738), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n959), .B(new_n964), .C1(G50), .C2(new_n789), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n958), .B1(new_n965), .B2(new_n312), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT47), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n946), .B1(new_n967), .B2(new_n788), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT112), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n725), .B2(new_n916), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n942), .A2(new_n970), .ZN(G387));
  AOI22_X1  g0771(.A1(G311), .A2(new_n954), .B1(new_n789), .B2(G303), .ZN(new_n972));
  INV_X1    g0772(.A(G322), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n972), .B1(new_n973), .B2(new_n746), .C1(new_n742), .C2(new_n947), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT48), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n738), .A2(new_n485), .B1(new_n739), .B2(new_n761), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT114), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT49), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n312), .B1(new_n732), .B2(G326), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n459), .C2(new_n743), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n742), .A2(new_n211), .B1(new_n743), .B2(new_n518), .ZN(new_n984));
  INV_X1    g0784(.A(new_n738), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(G77), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n732), .A2(G150), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n804), .A2(new_n568), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n986), .A2(new_n987), .A3(new_n988), .A4(new_n312), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n984), .B(new_n989), .C1(new_n341), .C2(new_n954), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n990), .B1(new_n264), .B2(new_n747), .C1(new_n361), .C2(new_n746), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n788), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n717), .B1(new_n660), .B2(new_n725), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n240), .A2(G45), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT113), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n425), .A2(G50), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  AOI21_X1  g0797(.A(G45), .B1(G68), .B2(G77), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n674), .A3(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n995), .A2(new_n767), .A3(new_n999), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(G107), .B2(new_n204), .C1(new_n674), .C2(new_n770), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n992), .B(new_n993), .C1(new_n772), .C2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n936), .B2(new_n941), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n671), .B1(new_n936), .B2(new_n713), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1003), .B1(new_n938), .B2(new_n1004), .ZN(G393));
  NAND2_X1  g0805(.A1(new_n931), .A2(new_n932), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n672), .B1(new_n1006), .B2(new_n937), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1007), .A2(new_n939), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G107), .A2(new_n796), .B1(new_n789), .B2(G294), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n750), .B2(new_n729), .C1(new_n973), .C2(new_n731), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n312), .B(new_n1010), .C1(G283), .C2(new_n985), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G317), .A2(new_n758), .B1(new_n753), .B2(G311), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT52), .Z(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1013), .C1(new_n459), .C2(new_n739), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT116), .Z(new_n1015));
  OAI22_X1  g0815(.A1(new_n746), .A2(new_n326), .B1(new_n742), .B2(new_n361), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT51), .Z(new_n1017));
  AOI21_X1  g0817(.A(new_n283), .B1(new_n732), .B2(G143), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n264), .B2(new_n738), .C1(new_n555), .C2(new_n743), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT115), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G77), .B2(new_n804), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n747), .A2(new_n425), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1017), .B(new_n1023), .C1(G50), .C2(new_n954), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n764), .B1(new_n1015), .B2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n772), .B1(new_n518), .B2(new_n204), .C1(new_n247), .C2(new_n943), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n906), .A2(new_n908), .A3(new_n723), .A4(new_n909), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1025), .A2(new_n717), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n941), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1028), .B1(new_n1006), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1008), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(G390));
  AOI21_X1  g0832(.A(new_n852), .B1(new_n777), .B2(new_n781), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n859), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n865), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n866), .A2(new_n876), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n864), .B1(new_n874), .B2(new_n850), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n711), .A2(new_n781), .A3(new_n653), .ZN(new_n1038));
  AND2_X1   g0838(.A1(new_n1038), .A2(new_n853), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1037), .B1(new_n1039), .B2(new_n1034), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n691), .A2(new_n859), .A3(G330), .A4(new_n781), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1036), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n866), .A2(new_n721), .A3(new_n876), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n954), .A2(G137), .B1(new_n804), .B2(G159), .ZN(new_n1049));
  XOR2_X1   g0849(.A(KEYINPUT54), .B(G143), .Z(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n747), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT119), .Z(new_n1053));
  AOI22_X1  g0853(.A1(new_n758), .A2(G128), .B1(new_n732), .B2(G125), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n1053), .A2(new_n312), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n796), .A2(G50), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n753), .A2(G132), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n738), .A2(new_n326), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT53), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n797), .B1(new_n213), .B2(new_n739), .C1(new_n485), .C2(new_n731), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n749), .A2(new_n555), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n742), .A2(new_n459), .B1(new_n747), .B2(new_n518), .ZN(new_n1063));
  NOR4_X1   g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n312), .A4(new_n1063), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1064), .B1(new_n460), .B2(new_n729), .C1(new_n761), .C2(new_n746), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n788), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n341), .A2(new_n812), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n1066), .A2(new_n716), .A3(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT120), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n1047), .A2(new_n941), .B1(new_n1048), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT118), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n451), .A2(G330), .A3(new_n691), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n880), .A2(new_n619), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n691), .A2(G330), .A3(new_n781), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n1034), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1039), .A2(new_n1042), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1033), .B1(new_n1076), .B2(new_n1042), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT117), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(new_n1042), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n855), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1039), .A2(new_n1042), .A3(new_n1076), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1073), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n672), .B1(new_n1087), .B2(new_n1046), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1044), .A2(new_n1045), .A3(new_n1084), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1071), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1085), .B1(new_n1091), .B2(new_n1074), .ZN(new_n1092));
  AOI211_X1 g0892(.A(KEYINPUT117), .B(new_n1073), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1042), .B1(new_n1036), .B2(new_n1040), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1036), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n1092), .A2(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AND4_X1   g0896(.A1(new_n1071), .A2(new_n1096), .A3(new_n671), .A4(new_n1089), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1070), .B1(new_n1090), .B2(new_n1097), .ZN(G378));
  NAND2_X1  g0898(.A1(new_n886), .A2(new_n887), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n888), .A2(new_n885), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1099), .A2(G330), .A3(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1102));
  NOR2_X1   g0902(.A1(new_n353), .A2(new_n355), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n612), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1102), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n618), .A2(new_n346), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n345), .A2(new_n824), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1104), .A2(new_n1106), .A3(new_n345), .A4(new_n824), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n889), .A2(G330), .A3(new_n1111), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1113), .A2(new_n878), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n878), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT122), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n863), .A2(new_n877), .ZN(new_n1118));
  AND4_X1   g0918(.A1(G330), .A2(new_n1111), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1111), .B1(new_n889), .B2(G330), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT122), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1117), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT123), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1095), .A2(new_n1094), .A3(new_n1079), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n1073), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1074), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT57), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT57), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1113), .A2(new_n878), .A3(new_n1114), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1131), .B1(new_n1121), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1074), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT123), .B1(new_n1089), .B2(new_n1074), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n671), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1130), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1111), .A2(new_n722), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n669), .A2(new_n312), .ZN(new_n1140));
  AOI211_X1 g0940(.A(G50), .B(new_n1140), .C1(new_n279), .C2(new_n476), .ZN(new_n1141));
  INV_X1    g0941(.A(G128), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n742), .A2(new_n1142), .B1(new_n747), .B2(new_n791), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1051), .A2(new_n738), .B1(new_n326), .B2(new_n739), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G125), .C2(new_n758), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n798), .B2(new_n729), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(G124), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n279), .B(new_n476), .C1(new_n731), .C2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G159), .B2(new_n796), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1141), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n986), .B1(new_n731), .B2(new_n761), .C1(new_n459), .C2(new_n746), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n954), .A2(G97), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n753), .A2(G107), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n796), .A2(new_n329), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1140), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n747), .A2(new_n427), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1153), .A2(new_n1157), .A3(new_n960), .A4(new_n1158), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT58), .Z(new_n1160));
  AOI21_X1  g0960(.A(new_n788), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n812), .A2(G50), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1139), .A2(new_n716), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1124), .B2(new_n941), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1138), .A2(new_n1164), .ZN(G375));
  NOR2_X1   g0965(.A1(new_n747), .A2(new_n326), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n739), .A2(new_n211), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n749), .A2(new_n361), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1156), .B1(new_n729), .B2(new_n1051), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n312), .B1(new_n731), .B2(new_n1142), .C1(new_n746), .C2(new_n798), .ZN(new_n1170));
  OR4_X1    g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1166), .B(new_n1171), .C1(G137), .C2(new_n753), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n959), .B1(G283), .B2(new_n753), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n283), .C1(new_n749), .C2(new_n518), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n746), .A2(new_n485), .B1(new_n747), .B2(new_n460), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1175), .B1(G116), .B2(new_n954), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT125), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n988), .B1(new_n750), .B2(new_n731), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1174), .B(new_n1178), .C1(new_n1177), .C2(new_n1176), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n764), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n720), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n717), .B(new_n1180), .C1(new_n859), .C2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n264), .B2(new_n811), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n941), .B(KEYINPUT124), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1091), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1082), .A2(new_n1073), .A3(new_n1083), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1087), .A2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1187), .B2(new_n926), .ZN(G381));
  INV_X1    g0988(.A(G375), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1190));
  AND2_X1   g0990(.A1(new_n1190), .A2(new_n1070), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G381), .A2(G384), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1031), .A2(new_n942), .A3(new_n970), .ZN(new_n1195));
  OR3_X1    g0995(.A1(new_n1195), .A2(G396), .A3(G393), .ZN(new_n1196));
  OR3_X1    g0996(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .ZN(G407));
  NAND3_X1  g0997(.A1(new_n1189), .A2(new_n651), .A3(new_n1191), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT126), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(G407), .A2(new_n1198), .A3(new_n1199), .A4(G213), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1192), .A2(new_n1194), .A3(new_n1196), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1198), .A2(G213), .ZN(new_n1202));
  OAI21_X1  g1002(.A(KEYINPUT126), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1200), .A2(new_n1203), .ZN(G409));
  NOR2_X1   g1004(.A1(new_n786), .A2(new_n814), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT60), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n672), .B1(new_n1186), .B2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n1079), .C1(new_n1206), .C2(new_n1186), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1185), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1205), .A2(new_n1209), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1213), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1212), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1210), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(G378), .B(new_n1164), .C1(new_n1130), .C2(new_n1137), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1121), .A2(new_n1132), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1163), .B1(new_n1220), .B2(new_n1184), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1123), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1122), .B1(new_n1121), .B2(new_n1132), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1222), .A2(new_n1223), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1224), .B2(new_n926), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1191), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1219), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n651), .A2(G213), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1218), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT127), .B1(new_n1229), .B2(KEYINPUT61), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT127), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT61), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1219), .A2(new_n1226), .B1(G213), .B2(new_n651), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1231), .B(new_n1232), .C1(new_n1233), .C2(new_n1218), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1216), .A2(new_n1210), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT62), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT62), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1233), .A2(new_n1238), .A3(new_n1235), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1230), .A2(new_n1234), .A3(new_n1237), .A4(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G390), .A2(G387), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1195), .ZN(new_n1242));
  XOR2_X1   g1042(.A(G393), .B(G396), .Z(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1243), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1241), .A2(new_n1195), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1240), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1236), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1247), .B1(new_n1249), .B2(KEYINPUT63), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1236), .B1(new_n1229), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(new_n1232), .A3(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1248), .A2(new_n1253), .ZN(G405));
  NAND2_X1  g1054(.A1(G375), .A2(new_n1191), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1219), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1247), .A2(new_n1219), .A3(new_n1255), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1235), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1257), .A2(new_n1258), .A3(new_n1235), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(G402));
endmodule


