//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G141gat), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208));
  AND2_X1   g007(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n210));
  INV_X1    g009(.A(G162gat), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n207), .B(new_n208), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(new_n208), .ZN(new_n215));
  XNOR2_X1  g014(.A(G141gat), .B(G148gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(KEYINPUT2), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(G197gat), .B(G204gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT22), .ZN(new_n220));
  INV_X1    g019(.A(G211gat), .ZN(new_n221));
  INV_X1    g020(.A(G218gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G211gat), .B(G218gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n219), .A3(new_n223), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT29), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n218), .B1(new_n229), .B2(KEYINPUT3), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n202), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n233), .A3(new_n217), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT72), .B(KEYINPUT29), .Z(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT71), .ZN(new_n238));
  INV_X1    g037(.A(new_n228), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n225), .B1(new_n223), .B2(new_n219), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n227), .A2(KEYINPUT71), .A3(new_n228), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  OAI211_X1 g043(.A(KEYINPUT80), .B(new_n218), .C1(new_n229), .C2(KEYINPUT3), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n232), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT79), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT79), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n249), .B(new_n236), .C1(new_n239), .C2(new_n240), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n233), .A3(new_n250), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n251), .A2(new_n218), .B1(new_n243), .B2(new_n237), .ZN(new_n252));
  INV_X1    g051(.A(new_n202), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n246), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255));
  OAI21_X1  g054(.A(G22gat), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G78gat), .B(G106gat), .Z(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n254), .B2(new_n255), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n251), .A2(new_n218), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(new_n244), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n202), .ZN(new_n264));
  INV_X1    g063(.A(G22gat), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n264), .A2(KEYINPUT81), .A3(new_n265), .A4(new_n246), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n256), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n261), .B1(new_n256), .B2(new_n266), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G64gat), .B(G92gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G36gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT73), .ZN(new_n272));
  INV_X1    g071(.A(G8gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G226gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NOR3_X1   g076(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n278));
  AND2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  AND2_X1   g084(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n287));
  OAI211_X1 g086(.A(KEYINPUT28), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n291), .A2(KEYINPUT67), .A3(KEYINPUT28), .A4(new_n285), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT65), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n284), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n279), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  OAI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n283), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT25), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n283), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT64), .B1(new_n283), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT64), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n313), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT23), .ZN(new_n316));
  INV_X1    g115(.A(G169gat), .ZN(new_n317));
  INV_X1    g116(.A(G176gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n279), .B1(new_n319), .B2(new_n302), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n309), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n277), .B1(new_n300), .B2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n282), .A2(new_n283), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n290), .A2(new_n292), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n323), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n235), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n243), .B(new_n324), .C1(new_n330), .C2(new_n277), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n299), .A2(new_n290), .A3(new_n292), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n323), .B1(new_n333), .B2(new_n325), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n276), .B1(new_n334), .B2(KEYINPUT29), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n243), .B1(new_n335), .B2(new_n324), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n275), .B1(new_n332), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT30), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n276), .B1(new_n328), .B2(new_n329), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n341), .B1(new_n300), .B2(new_n323), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n340), .B1(new_n276), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n331), .B1(new_n343), .B2(new_n243), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n275), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n338), .A2(new_n339), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n344), .A2(KEYINPUT30), .A3(new_n275), .ZN(new_n348));
  INV_X1    g147(.A(new_n243), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n328), .A2(new_n329), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n277), .B1(new_n350), .B2(new_n341), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n349), .B1(new_n351), .B2(new_n340), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n331), .A3(new_n274), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G120gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(G113gat), .ZN(new_n357));
  INV_X1    g156(.A(G113gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G120gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT1), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G134gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G127gat), .ZN(new_n364));
  INV_X1    g163(.A(G127gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(G134gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G127gat), .B(G134gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(new_n369), .A3(new_n361), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT4), .B1(new_n218), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n208), .B1(new_n213), .B2(new_n207), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT75), .A2(G155gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(G162gat), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n216), .B1(new_n376), .B2(KEYINPUT2), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n377), .B2(new_n208), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n360), .A2(new_n369), .A3(new_n361), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n360), .A2(new_n361), .B1(new_n364), .B2(new_n366), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT76), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n380), .B2(new_n381), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n385), .A2(new_n234), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n384), .A2(new_n389), .A3(KEYINPUT5), .A4(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n384), .A2(new_n389), .A3(new_n390), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT5), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n382), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n386), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n378), .ZN(new_n396));
  INV_X1    g195(.A(new_n390), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n391), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G57gat), .B(G85gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n403), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n402), .A2(new_n406), .ZN(new_n408));
  OAI221_X1 g207(.A(new_n391), .B1(new_n407), .B2(new_n408), .C1(new_n392), .C2(new_n398), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT78), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n399), .A2(new_n404), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT6), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT6), .B1(new_n399), .B2(new_n404), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT78), .A3(new_n409), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n269), .B1(new_n355), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT68), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT69), .ZN(new_n422));
  XOR2_X1   g221(.A(G15gat), .B(G43gat), .Z(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n371), .B1(new_n300), .B2(new_n323), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n328), .A2(new_n382), .A3(new_n329), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n424), .B1(new_n428), .B2(KEYINPUT33), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT70), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n426), .A2(new_n425), .A3(new_n427), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n430), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n424), .C1(KEYINPUT33), .C2(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT32), .ZN(new_n436));
  OR3_X1    g235(.A1(new_n428), .A2(new_n436), .A3(KEYINPUT34), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT34), .B1(new_n428), .B2(new_n436), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n432), .A2(new_n434), .A3(new_n438), .A4(new_n437), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n440), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n419), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT40), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n390), .B1(new_n384), .B2(new_n389), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n396), .A2(new_n397), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NOR3_X1   g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n218), .A2(new_n371), .A3(KEYINPUT4), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n379), .B1(new_n378), .B2(new_n382), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n234), .A2(new_n386), .A3(new_n388), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n233), .B1(new_n214), .B2(new_n217), .ZN(new_n457));
  OAI22_X1  g256(.A1(new_n454), .A2(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n452), .A3(new_n397), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT82), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n408), .B2(new_n407), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n449), .B1(new_n453), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n462), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n391), .B(new_n466), .C1(new_n392), .C2(new_n398), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n458), .A2(new_n397), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n396), .A2(new_n397), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT39), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(KEYINPUT40), .A3(new_n463), .A4(new_n459), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n465), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n448), .B1(new_n355), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT37), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n331), .C1(new_n343), .C2(new_n243), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n352), .B2(new_n331), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n274), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT38), .ZN(new_n479));
  AOI211_X1 g278(.A(KEYINPUT74), .B(new_n274), .C1(new_n352), .C2(new_n331), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n345), .B1(new_n344), .B2(new_n275), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n416), .A2(new_n467), .B1(new_n414), .B2(KEYINPUT6), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n349), .B(new_n324), .C1(new_n330), .C2(new_n277), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n484), .B1(new_n343), .B2(new_n349), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n475), .B1(new_n485), .B2(new_n474), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT38), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n274), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n479), .A2(new_n482), .A3(new_n483), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n347), .A2(new_n354), .ZN(new_n490));
  INV_X1    g289(.A(new_n472), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT83), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n473), .A2(new_n269), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n269), .A2(new_n442), .ZN(new_n494));
  INV_X1    g293(.A(new_n483), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n496));
  NAND4_X1  g295(.A1(new_n494), .A2(new_n355), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n355), .A2(new_n418), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n269), .A2(new_n442), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT35), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n447), .A2(new_n493), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n502));
  XNOR2_X1  g301(.A(KEYINPUT87), .B(G169gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT86), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT12), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G43gat), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(G50gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(G50gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT15), .A3(new_n513), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT89), .B(G50gat), .Z(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n511), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT15), .B1(new_n516), .B2(new_n512), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT88), .B(G29gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  OR3_X1    g320(.A1(new_n520), .A2(G29gat), .A3(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n514), .B1(new_n517), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n514), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT17), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528));
  XOR2_X1   g327(.A(G15gat), .B(G22gat), .Z(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n533));
  INV_X1    g332(.A(G1gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT16), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(G1gat), .B1(new_n531), .B2(new_n533), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n528), .B(new_n273), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n531), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n534), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n528), .A2(new_n273), .ZN(new_n541));
  NAND2_X1  g340(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n524), .A2(new_n546), .A3(new_n525), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n524), .A2(new_n525), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n538), .A3(new_n544), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT18), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n545), .A2(new_n526), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n551), .B(KEYINPUT13), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n548), .A2(KEYINPUT18), .A3(new_n550), .A4(new_n551), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n554), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n510), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n509), .A2(new_n559), .A3(new_n554), .A4(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT92), .B1(new_n501), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n493), .A2(new_n447), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n497), .A2(new_n500), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n564), .ZN(new_n571));
  XNOR2_X1  g370(.A(G127gat), .B(G155gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT20), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  INV_X1    g374(.A(G64gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G57gat), .ZN(new_n577));
  INV_X1    g376(.A(G57gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(G64gat), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n581), .A2(KEYINPUT93), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(KEYINPUT93), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G71gat), .B(G78gat), .Z(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n585), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n587), .B(new_n580), .C1(new_n583), .C2(new_n582), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n586), .A2(new_n588), .A3(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n545), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n590), .B(KEYINPUT96), .ZN(new_n591));
  INV_X1    g390(.A(G231gat), .ZN(new_n592));
  INV_X1    g391(.A(G233gat), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n590), .B(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(G231gat), .A3(G233gat), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n574), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G183gat), .B(G211gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT95), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT19), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n588), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n602), .B(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n594), .A2(new_n597), .A3(new_n574), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n606), .ZN(new_n609));
  INV_X1    g408(.A(new_n607), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n609), .B1(new_n610), .B2(new_n598), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  INV_X1    g413(.A(G92gat), .ZN(new_n615));
  AOI22_X1  g414(.A1(KEYINPUT8), .A2(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n614), .B2(new_n615), .ZN(new_n618));
  NAND3_X1  g417(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G99gat), .B(G106gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n527), .A2(new_n622), .A3(new_n547), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n620), .A2(new_n621), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n620), .A2(new_n621), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(G232gat), .A2(G233gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(new_n549), .A2(new_n626), .B1(KEYINPUT41), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G190gat), .B(G218gat), .Z(new_n629));
  NAND3_X1  g428(.A1(new_n623), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G134gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n211), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n629), .B1(new_n623), .B2(new_n628), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n630), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n623), .A2(new_n628), .ZN(new_n637));
  INV_X1    g436(.A(new_n633), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n637), .B(new_n629), .C1(KEYINPUT98), .C2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n636), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n640), .B1(new_n636), .B2(new_n639), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n612), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G230gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n593), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n588), .A3(new_n586), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT10), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n603), .A2(new_n622), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n626), .A2(KEYINPUT10), .A3(new_n588), .A4(new_n586), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n646), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n649), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n646), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(new_n318), .ZN(new_n658));
  INV_X1    g457(.A(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n653), .A2(new_n655), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n566), .A2(new_n571), .A3(new_n644), .A4(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n418), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT99), .B(G1gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1324gat));
  OAI21_X1  g468(.A(G8gat), .B1(new_n666), .B2(new_n355), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT100), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT16), .ZN(new_n672));
  AOI211_X1 g471(.A(new_n355), .B(new_n666), .C1(new_n672), .C2(new_n273), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  NAND2_X1  g473(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n674), .B1(new_n673), .B2(new_n675), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(G1325gat));
  AND3_X1   g477(.A1(new_n440), .A2(KEYINPUT36), .A3(new_n441), .ZN(new_n679));
  AOI21_X1  g478(.A(KEYINPUT36), .B1(new_n440), .B2(new_n441), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n666), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n442), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n683), .A2(G15gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n666), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT101), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n666), .A2(new_n269), .ZN(new_n687));
  XOR2_X1   g486(.A(KEYINPUT43), .B(G22gat), .Z(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n643), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n501), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n489), .A2(new_n269), .ZN(new_n693));
  AOI211_X1 g492(.A(new_n448), .B(new_n472), .C1(new_n347), .C2(new_n354), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT83), .B1(new_n490), .B2(new_n491), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n416), .A2(KEYINPUT78), .A3(new_n409), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT78), .B1(new_n416), .B2(new_n409), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n490), .B1(new_n699), .B2(new_n415), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n681), .B1(new_n700), .B2(new_n269), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT102), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n493), .A2(new_n447), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n568), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n643), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n692), .B1(new_n706), .B2(new_n690), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n608), .A2(new_n611), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n664), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n418), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n564), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT103), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT103), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n710), .A2(new_n714), .A3(new_n711), .A4(new_n564), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n518), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n566), .A2(new_n571), .A3(new_n643), .A4(new_n709), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n717), .A2(new_n418), .A3(new_n518), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT45), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1328gat));
  NOR2_X1   g519(.A1(new_n717), .A2(G36gat), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n490), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT104), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n724), .A3(new_n490), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n707), .A2(new_n490), .A3(new_n564), .A4(new_n709), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT105), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(G36gat), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n723), .A2(KEYINPUT46), .A3(new_n725), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n728), .A2(new_n733), .A3(new_n734), .ZN(G1329gat));
  NOR3_X1   g534(.A1(new_n717), .A2(G43gat), .A3(new_n683), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n707), .A2(new_n446), .A3(new_n564), .A4(new_n709), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G43gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g538(.A1(new_n717), .A2(new_n515), .A3(new_n269), .ZN(new_n740));
  INV_X1    g539(.A(new_n269), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n707), .A2(new_n741), .A3(new_n564), .A4(new_n709), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(new_n515), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g543(.A1(new_n612), .A2(new_n643), .A3(new_n564), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n705), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n664), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n418), .ZN(new_n748));
  XNOR2_X1  g547(.A(KEYINPUT106), .B(G57gat), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n748), .B(new_n749), .ZN(G1332gat));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n664), .A3(new_n490), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OR3_X1    g551(.A1(new_n751), .A2(KEYINPUT107), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(new_n751), .B2(new_n752), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n755), .B(new_n756), .ZN(G1333gat));
  AND4_X1   g556(.A1(G71gat), .A2(new_n705), .A3(new_n664), .A4(new_n745), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n758), .A2(KEYINPUT108), .A3(new_n446), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT108), .B1(new_n758), .B2(new_n446), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n747), .A2(new_n683), .ZN(new_n761));
  OAI22_X1  g560(.A1(new_n759), .A2(new_n760), .B1(new_n761), .B2(G71gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n747), .A2(new_n269), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g564(.A1(new_n708), .A2(new_n564), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n705), .A2(new_n643), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n643), .A4(new_n766), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n665), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n711), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT44), .B1(new_n705), .B2(new_n643), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n766), .A2(new_n664), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n773), .A2(new_n692), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n418), .A2(new_n614), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n770), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n664), .A3(new_n490), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n615), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n775), .A2(G92gat), .A3(new_n490), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(G92gat), .B1(new_n771), .B2(new_n490), .ZN(new_n786));
  INV_X1    g585(.A(new_n774), .ZN(new_n787));
  AND4_X1   g586(.A1(G92gat), .A2(new_n707), .A3(new_n490), .A4(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n781), .B(KEYINPUT52), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n785), .A2(new_n789), .ZN(G1337gat));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n446), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(G99gat), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(G99gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n771), .A2(new_n795), .A3(new_n442), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n794), .A2(new_n796), .ZN(G1338gat));
  INV_X1    g596(.A(KEYINPUT111), .ZN(new_n798));
  NOR4_X1   g597(.A1(new_n773), .A2(new_n692), .A3(new_n269), .A4(new_n774), .ZN(new_n799));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n706), .A2(new_n690), .ZN(new_n802));
  INV_X1    g601(.A(new_n692), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n802), .A2(new_n741), .A3(new_n803), .A4(new_n787), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n804), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n269), .A2(G106gat), .A3(new_n665), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT112), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n778), .A2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n801), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n804), .A2(G106gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n778), .A2(new_n806), .ZN(new_n812));
  AND4_X1   g611(.A1(KEYINPUT113), .A2(new_n811), .A3(new_n810), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n804), .B2(G106gat), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n814), .B2(new_n812), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n809), .A2(new_n810), .B1(new_n813), .B2(new_n815), .ZN(G1339gat));
  NAND3_X1  g615(.A1(new_n650), .A2(new_n651), .A3(new_n646), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n662), .B1(new_n652), .B2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(KEYINPUT55), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n820), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n564), .A2(new_n663), .A3(new_n821), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n550), .A2(new_n555), .A3(new_n557), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n550), .A2(new_n555), .A3(KEYINPUT115), .A4(new_n557), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n548), .A2(new_n550), .ZN(new_n831));
  INV_X1    g630(.A(new_n551), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT114), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834));
  AOI211_X1 g633(.A(new_n834), .B(new_n551), .C1(new_n548), .C2(new_n550), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n830), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n508), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n664), .B(new_n563), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n643), .B1(new_n825), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n831), .A2(new_n832), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n834), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n831), .A2(KEYINPUT114), .A3(new_n832), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n508), .B1(new_n843), .B2(new_n830), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n844), .B(new_n563), .C1(new_n641), .C2(new_n642), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n824), .A2(new_n663), .A3(new_n821), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n612), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n708), .A2(new_n691), .A3(new_n665), .A4(new_n565), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n499), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n711), .A3(new_n355), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n565), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(new_n358), .ZN(G1340gat));
  OAI21_X1  g652(.A(G120gat), .B1(new_n851), .B2(new_n665), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n664), .A2(new_n356), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT116), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n854), .B1(new_n851), .B2(new_n856), .ZN(G1341gat));
  NOR2_X1   g656(.A1(new_n851), .A2(new_n612), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n858), .B(new_n365), .ZN(G1342gat));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n363), .ZN(new_n861));
  OR3_X1    g660(.A1(new_n851), .A2(new_n691), .A3(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT117), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n363), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n863), .B(new_n864), .ZN(G1343gat));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n838), .A2(KEYINPUT118), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n844), .A2(new_n868), .A3(new_n664), .A4(new_n563), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n825), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n847), .B1(new_n870), .B2(new_n691), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n849), .B1(new_n871), .B2(new_n708), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n866), .B1(new_n872), .B2(new_n741), .ZN(new_n873));
  AOI211_X1 g672(.A(KEYINPUT57), .B(new_n269), .C1(new_n848), .C2(new_n849), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n711), .A2(new_n355), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n446), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR4_X1   g676(.A1(new_n873), .A2(new_n874), .A3(new_n565), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT119), .B1(new_n878), .B2(new_n205), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n870), .A2(new_n691), .ZN(new_n882));
  INV_X1    g681(.A(new_n847), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n708), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n849), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n741), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n269), .B1(new_n848), .B2(new_n849), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n866), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n887), .A2(new_n564), .A3(new_n876), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G141gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n848), .A2(new_n849), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n741), .ZN(new_n893));
  NOR4_X1   g692(.A1(new_n893), .A2(G141gat), .A3(new_n565), .A4(new_n877), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n881), .B1(new_n891), .B2(new_n895), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT120), .B(new_n894), .C1(new_n890), .C2(G141gat), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n880), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n895), .B1(new_n878), .B2(new_n205), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT120), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT58), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n891), .B2(KEYINPUT119), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n891), .A2(new_n881), .A3(new_n895), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n898), .A2(new_n904), .ZN(G1344gat));
  NOR2_X1   g704(.A1(new_n893), .A2(new_n877), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(new_n203), .A3(new_n664), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n866), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n872), .B2(new_n741), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n664), .B(new_n876), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n203), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n908), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n887), .A2(new_n876), .A3(new_n889), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n908), .B1(new_n916), .B2(new_n665), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n203), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n907), .B1(new_n915), .B2(new_n918), .ZN(G1345gat));
  NOR2_X1   g718(.A1(new_n209), .A2(new_n210), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n906), .B2(new_n708), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n916), .A2(new_n612), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n922), .B2(new_n920), .ZN(G1346gat));
  AOI21_X1  g722(.A(G162gat), .B1(new_n906), .B2(new_n643), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n916), .A2(new_n691), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n711), .A2(new_n355), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n850), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(new_n565), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(new_n317), .ZN(G1348gat));
  NOR2_X1   g729(.A1(new_n928), .A2(new_n665), .ZN(new_n931));
  XOR2_X1   g730(.A(KEYINPUT122), .B(G176gat), .Z(new_n932));
  XNOR2_X1  g731(.A(new_n931), .B(new_n932), .ZN(G1349gat));
  INV_X1    g732(.A(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g733(.A(G183gat), .B1(new_n928), .B2(new_n612), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(new_n291), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n928), .A2(new_n612), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n928), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n708), .A3(new_n291), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n941), .A2(KEYINPUT123), .A3(new_n935), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(KEYINPUT60), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n936), .A2(new_n938), .A3(KEYINPUT60), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(KEYINPUT124), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n945), .B1(new_n947), .B2(new_n943), .ZN(G1350gat));
  NAND2_X1  g747(.A1(new_n940), .A2(new_n643), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G190gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT61), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n950), .B(KEYINPUT125), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n953), .B(new_n956), .C1(G190gat), .C2(new_n949), .ZN(G1351gat));
  OR2_X1    g756(.A1(new_n909), .A2(new_n910), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n446), .A2(new_n711), .A3(new_n355), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT126), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(G197gat), .B1(new_n961), .B2(new_n565), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n888), .A2(new_n959), .ZN(new_n963));
  INV_X1    g762(.A(G197gat), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n964), .A3(new_n564), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1352gat));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n659), .A3(new_n664), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n967), .B(KEYINPUT62), .Z(new_n968));
  NAND3_X1  g767(.A1(new_n958), .A2(new_n664), .A3(new_n960), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n970), .B2(new_n659), .ZN(G1353gat));
  NAND3_X1  g770(.A1(new_n963), .A2(new_n221), .A3(new_n708), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n958), .A2(new_n708), .A3(new_n960), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n973), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n973), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n972), .B1(new_n974), .B2(new_n975), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n961), .B2(new_n691), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n963), .A2(new_n222), .A3(new_n643), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(G1355gat));
endmodule


