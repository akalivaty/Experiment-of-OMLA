//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n462), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n462), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n476), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT69), .Z(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n485), .B(new_n486), .C1(new_n464), .C2(new_n463), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n462), .A2(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n473), .B2(new_n474), .ZN(new_n489));
  XOR2_X1   g064(.A(KEYINPUT71), .B(KEYINPUT4), .Z(new_n490));
  OAI21_X1  g065(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT70), .B1(new_n462), .B2(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n492), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT72), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(KEYINPUT72), .A2(KEYINPUT6), .A3(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n507), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT5), .B(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n509), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n514), .A2(new_n517), .ZN(G166));
  NAND2_X1  g093(.A1(new_n508), .A2(G51), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(KEYINPUT7), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n519), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(KEYINPUT5), .A2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n506), .B2(new_n507), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n528), .A2(G90), .B1(new_n533), .B2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n508), .A2(G52), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  AOI22_X1  g112(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n538), .A2(new_n516), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n508), .A2(G43), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n528), .A2(G81), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  AOI22_X1  g123(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n516), .ZN(new_n550));
  INV_X1    g125(.A(G53), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(KEYINPUT9), .ZN(new_n553));
  OAI211_X1 g128(.A(new_n508), .B(new_n553), .C1(new_n552), .C2(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT9), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n511), .A2(G543), .ZN(new_n556));
  OAI211_X1 g131(.A(KEYINPUT73), .B(new_n555), .C1(new_n556), .C2(new_n551), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n528), .A2(G91), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n550), .A2(new_n554), .A3(new_n557), .A4(new_n558), .ZN(G299));
  INV_X1    g134(.A(G168), .ZN(G286));
  INV_X1    g135(.A(G166), .ZN(G303));
  NAND3_X1  g136(.A1(new_n511), .A2(G87), .A3(new_n512), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  INV_X1    g140(.A(G49), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n556), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n508), .A2(KEYINPUT74), .A3(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n564), .A2(KEYINPUT75), .A3(new_n567), .A4(new_n568), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n511), .A2(G86), .A3(new_n512), .ZN(new_n575));
  INV_X1    g150(.A(new_n507), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT6), .B1(KEYINPUT72), .B2(G651), .ZN(new_n577));
  OAI211_X1 g152(.A(G48), .B(G543), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AND2_X1   g153(.A1(G73), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n512), .B2(G61), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n575), .B(new_n578), .C1(new_n580), .C2(new_n516), .ZN(G305));
  NAND2_X1  g156(.A1(new_n528), .A2(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n508), .A2(G47), .ZN(new_n583));
  NAND2_X1  g158(.A1(G72), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G60), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n527), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n583), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(KEYINPUT76), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n528), .A2(G85), .B1(new_n586), .B2(G651), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n583), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OR3_X1    g171(.A1(new_n513), .A2(KEYINPUT77), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT77), .B1(new_n513), .B2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(KEYINPUT10), .A3(new_n598), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n527), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(G651), .B1(G54), .B2(new_n508), .ZN(new_n606));
  AND3_X1   g181(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n595), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT78), .Z(G297));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n542), .A2(new_n610), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n618), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n473), .A2(new_n474), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n469), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT80), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n475), .A2(G135), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT81), .Z(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI22_X1  g209(.A1(new_n631), .A2(new_n632), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  AOI22_X1  g210(.A1(new_n633), .A2(new_n635), .B1(new_n477), .B2(G123), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G2096), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(new_n638), .B1(new_n625), .B2(new_n626), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n628), .B(new_n639), .C1(new_n638), .C2(new_n637), .ZN(G156));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT14), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n647), .B(new_n651), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n647), .B(new_n651), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n653), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n655), .A2(new_n657), .A3(G14), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT83), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n660));
  NAND4_X1  g235(.A1(new_n655), .A2(new_n657), .A3(new_n660), .A4(G14), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT17), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n666), .A2(new_n667), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n668), .B2(new_n664), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n671), .B(new_n673), .Z(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(KEYINPUT86), .B(KEYINPUT87), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1961), .B(G1966), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT85), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(new_n684), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n686), .A2(new_n687), .ZN(new_n690));
  MUX2_X1   g265(.A(new_n684), .B(new_n689), .S(new_n690), .Z(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n684), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n691), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n696), .B1(new_n691), .B2(new_n694), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n682), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1981), .B(G1986), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(new_n694), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(new_n695), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n681), .A3(new_n697), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n702), .B1(new_n700), .B2(new_n705), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n680), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n698), .A2(new_n682), .A3(new_n699), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n681), .B1(new_n704), .B2(new_n697), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n701), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n712), .A2(new_n679), .A3(new_n706), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(G229));
  NOR2_X1   g290(.A1(G4), .A2(G16), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n607), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT91), .B(G1348), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  AOI22_X1  g295(.A1(new_n475), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n477), .A2(G129), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT26), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n725), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(KEYINPUT95), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n731), .B(KEYINPUT95), .C1(G29), .C2(G32), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT27), .B(G1996), .Z(new_n734));
  AND3_X1   g309(.A1(new_n732), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n732), .B2(new_n733), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n719), .B(new_n720), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G35), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT97), .Z(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(new_n482), .B2(G29), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2090), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n637), .A2(G29), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT96), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n739), .A2(G27), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G164), .B2(new_n739), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n475), .A2(G139), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n621), .A2(G127), .ZN(new_n757));
  NAND2_X1  g332(.A1(G115), .A2(G2104), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n462), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(G29), .B1(new_n756), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G33), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(G29), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2072), .Z(new_n763));
  AND2_X1   g338(.A1(KEYINPUT24), .A2(G34), .ZN(new_n764));
  NOR2_X1   g339(.A1(KEYINPUT24), .A2(G34), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n739), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT93), .Z(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G29), .B2(G160), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n763), .B1(G2084), .B2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G16), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n770), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G1966), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(G28), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n739), .B1(new_n774), .B2(G28), .ZN(new_n776));
  AND2_X1   g351(.A1(KEYINPUT31), .A2(G11), .ZN(new_n777));
  NOR2_X1   g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  OAI22_X1  g353(.A1(new_n775), .A2(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n768), .B2(G2084), .ZN(new_n780));
  NOR2_X1   g355(.A1(G171), .A2(new_n770), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G5), .B2(new_n770), .ZN(new_n782));
  INV_X1    g357(.A(G1961), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n752), .A2(new_n769), .A3(new_n773), .A4(new_n784), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n770), .A2(G20), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT23), .ZN(new_n788));
  INV_X1    g363(.A(G299), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n770), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(G1956), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n770), .A2(G19), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n543), .B2(new_n770), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1341), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n739), .A2(G26), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n475), .A2(G140), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n477), .A2(G128), .ZN(new_n799));
  OR2_X1    g374(.A1(G104), .A2(G2105), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n798), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n797), .B1(new_n803), .B2(new_n739), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  NOR4_X1   g380(.A1(new_n786), .A2(new_n791), .A3(new_n794), .A4(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n738), .A2(new_n745), .A3(new_n785), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n770), .A2(G23), .ZN(new_n808));
  INV_X1    g383(.A(new_n569), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n770), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n770), .A2(G22), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G166), .B2(new_n770), .ZN(new_n814));
  INV_X1    g389(.A(G1971), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  MUX2_X1   g391(.A(G6), .B(G305), .S(G16), .Z(new_n817));
  XOR2_X1   g392(.A(KEYINPUT32), .B(G1981), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n812), .A2(new_n816), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT34), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n593), .A2(G16), .ZN(new_n822));
  OR2_X1    g397(.A1(G16), .A2(G24), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n822), .A2(G1986), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(G1986), .B1(new_n822), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  NOR3_X1   g402(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n828));
  OAI221_X1 g403(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n475), .A2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n477), .A2(G119), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  MUX2_X1   g407(.A(G25), .B(new_n832), .S(G29), .Z(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT89), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n824), .A2(new_n825), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT34), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n812), .A2(new_n838), .A3(new_n816), .A4(new_n819), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(KEYINPUT90), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT90), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n821), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(KEYINPUT36), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n807), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT99), .ZN(G311));
  XNOR2_X1  g421(.A(new_n845), .B(KEYINPUT100), .ZN(G150));
  NAND2_X1  g422(.A1(new_n508), .A2(G55), .ZN(new_n848));
  INV_X1    g423(.A(G93), .ZN(new_n849));
  AOI22_X1  g424(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n850));
  OAI221_X1 g425(.A(new_n848), .B1(new_n513), .B2(new_n849), .C1(new_n850), .C2(new_n516), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n852), .A2(new_n542), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n542), .A2(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n607), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n859));
  AOI21_X1  g434(.A(G860), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(new_n859), .B2(new_n858), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n852), .A2(G860), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT37), .Z(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(G145));
  XNOR2_X1  g439(.A(new_n729), .B(new_n803), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n477), .A2(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n462), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(G142), .B2(new_n475), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n865), .B(new_n870), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n756), .A2(KEYINPUT104), .A3(new_n759), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n499), .A2(new_n873), .A3(new_n500), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n873), .B1(new_n499), .B2(new_n500), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n491), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n872), .B(new_n876), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n624), .B(new_n832), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n871), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(G160), .B(KEYINPUT102), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n482), .B(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(new_n637), .Z(new_n883));
  AOI21_X1  g458(.A(G37), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n884), .B1(new_n883), .B2(new_n880), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g461(.A1(new_n588), .A2(KEYINPUT76), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n591), .A2(new_n590), .A3(new_n583), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n887), .A2(KEYINPUT105), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT105), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n889), .A2(new_n890), .A3(new_n809), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n589), .B2(new_n592), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT105), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n569), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(G166), .B(G305), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n891), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n809), .B1(new_n889), .B2(new_n890), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(new_n569), .A3(new_n894), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(KEYINPUT42), .B1(new_n897), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT106), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n891), .B2(new_n895), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n898), .A3(new_n900), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT106), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT42), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n607), .A2(new_n789), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n617), .A2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT41), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(KEYINPUT41), .A3(new_n911), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n855), .A2(new_n618), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n853), .B(new_n854), .C1(G559), .C2(new_n617), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n914), .A2(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n906), .B2(KEYINPUT42), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT42), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n904), .A2(KEYINPUT107), .A3(new_n923), .A4(new_n905), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n909), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n920), .B1(new_n909), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n852), .A2(new_n610), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(G295));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n928), .A2(new_n931), .A3(new_n929), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n931), .B1(new_n928), .B2(new_n929), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(G331));
  INV_X1    g509(.A(G37), .ZN(new_n935));
  XNOR2_X1  g510(.A(G171), .B(G168), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(new_n853), .A3(new_n854), .ZN(new_n937));
  INV_X1    g512(.A(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n855), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n914), .A2(new_n915), .A3(new_n937), .A4(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n937), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n936), .B1(new_n853), .B2(new_n854), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n911), .B(new_n910), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n906), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n935), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n945), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n949), .A2(KEYINPUT109), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT109), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n944), .B2(new_n945), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n947), .B(new_n948), .C1(new_n950), .C2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n949), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT43), .B1(new_n954), .B2(new_n946), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n947), .B(KEYINPUT43), .C1(new_n950), .C2(new_n952), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n948), .B1(new_n954), .B2(new_n946), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n958), .B1(new_n957), .B2(new_n961), .ZN(G397));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n876), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(new_n492), .B2(new_n501), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n465), .A2(new_n466), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G2105), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n468), .A2(new_n470), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(G40), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n972), .A2(G2084), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT45), .B1(new_n876), .B2(new_n964), .ZN(new_n974));
  NAND2_X1  g549(.A1(G160), .A2(G40), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT119), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT119), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n501), .A2(KEYINPUT103), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n499), .A2(new_n873), .A3(new_n500), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n980), .B2(new_n491), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n977), .B(new_n971), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(new_n501), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n983), .B2(new_n491), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT45), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n976), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1966), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n973), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(G168), .A2(G8), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2090), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n991), .A2(new_n965), .A3(new_n967), .A4(new_n971), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n975), .B1(new_n966), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n995));
  AOI21_X1  g570(.A(G1971), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(G8), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  NOR2_X1   g573(.A1(G166), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT55), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1000), .B(G8), .C1(new_n996), .C2(new_n992), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(KEYINPUT63), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  NAND2_X1  g580(.A1(G305), .A2(G1981), .ZN(new_n1006));
  INV_X1    g581(.A(G61), .ZN(new_n1007));
  OR2_X1    g582(.A1(KEYINPUT5), .A2(G543), .ZN(new_n1008));
  NAND2_X1  g583(.A1(KEYINPUT5), .A2(G543), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(G651), .B1(new_n1010), .B2(new_n579), .ZN(new_n1011));
  INV_X1    g586(.A(G1981), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n575), .A4(new_n578), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(KEYINPUT115), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT115), .ZN(new_n1015));
  NAND3_X1  g590(.A1(G305), .A2(new_n1015), .A3(G1981), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1005), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n876), .A2(new_n971), .A3(new_n964), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G8), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1014), .A2(new_n1005), .A3(new_n1016), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n564), .A2(G1976), .A3(new_n567), .A4(new_n568), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n571), .A2(new_n572), .A3(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1019), .A2(G8), .A3(new_n1025), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1023), .A2(new_n1028), .A3(KEYINPUT116), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(new_n1024), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1033), .B2(new_n1029), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1014), .A2(new_n1005), .A3(new_n1016), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1035), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1004), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT118), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1023), .A2(new_n1028), .A3(KEYINPUT118), .A4(new_n1030), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n963), .B1(new_n876), .B2(new_n964), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n963), .B(new_n964), .C1(new_n492), .C2(new_n501), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n971), .ZN(new_n1046));
  NOR3_X1   g621(.A1(new_n1044), .A2(new_n1046), .A3(G2090), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1043), .B1(new_n1047), .B2(new_n996), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n964), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n971), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n815), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n975), .B1(new_n984), .B2(new_n963), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(new_n991), .C1(new_n963), .C2(new_n981), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1053), .A3(KEYINPUT117), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1048), .A2(G8), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1001), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1042), .A2(new_n1056), .A3(new_n1003), .A4(new_n990), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n990), .A2(new_n1038), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1003), .B1(new_n1037), .B2(new_n1031), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1026), .B(new_n573), .C1(new_n1035), .C2(new_n1017), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1020), .B1(new_n1061), .B2(new_n1013), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT121), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1004), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1037), .A2(new_n1031), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n990), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1063), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1003), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1073), .B1(new_n1001), .B2(new_n1055), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n1042), .ZN(new_n1075));
  INV_X1    g650(.A(new_n974), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n969), .A2(KEYINPUT53), .A3(G40), .A4(new_n750), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n970), .A2(KEYINPUT123), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1076), .A2(new_n995), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(new_n1081), .B(KEYINPUT124), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT53), .B1(new_n1083), .B2(new_n750), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n783), .B2(new_n972), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(G301), .B(KEYINPUT54), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n986), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1091), .A3(new_n1087), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1075), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(G299), .B(KEYINPUT57), .Z(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  AND2_X1   g671(.A1(new_n1083), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(G1956), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1095), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1019), .ZN(new_n1102));
  INV_X1    g677(.A(G2067), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n972), .A2(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1100), .B1(new_n617), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1083), .A2(new_n1096), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n1094), .C1(G1956), .C2(new_n1098), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  AND3_X1   g684(.A1(new_n1100), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1100), .B2(new_n1107), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n994), .A2(new_n995), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT58), .B(G1341), .ZN(new_n1114));
  OAI22_X1  g689(.A1(new_n1113), .A2(G1996), .B1(new_n1102), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n1116), .A3(new_n543), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n617), .B1(new_n1104), .B2(KEYINPUT60), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(KEYINPUT60), .B2(new_n1104), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n617), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1108), .B1(new_n1112), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n988), .A2(G168), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G8), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n988), .A2(G168), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT51), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n998), .B1(new_n988), .B2(G168), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT51), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1093), .A2(new_n1125), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1128), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1131), .B1(new_n1135), .B2(new_n1130), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1132), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT62), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1129), .A2(new_n1139), .A3(new_n1132), .ZN(new_n1140));
  AOI21_X1  g715(.A(G301), .B1(new_n1085), .B2(new_n1091), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1074), .A2(new_n1141), .A3(new_n1042), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1065), .A2(new_n1072), .A3(new_n1134), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n974), .A2(new_n971), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT112), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n802), .B(G2067), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT113), .ZN(new_n1150));
  INV_X1    g725(.A(new_n834), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n832), .A2(new_n1151), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n832), .A2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1147), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OR2_X1    g729(.A1(new_n1145), .A2(G1996), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1155), .A2(KEYINPUT111), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(KEYINPUT111), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1146), .A2(new_n730), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1158), .A2(new_n730), .B1(new_n1159), .B2(G1996), .ZN(new_n1160));
  OR2_X1    g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  NAND2_X1  g736(.A1(G290), .A2(G1986), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(KEYINPUT110), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1145), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1163), .B(new_n1164), .C1(KEYINPUT110), .C2(new_n1162), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1150), .A2(new_n1154), .A3(new_n1160), .A4(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(KEYINPUT114), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1144), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1158), .A2(KEYINPUT46), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1156), .A2(new_n1170), .A3(new_n1157), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1147), .B1(new_n729), .B2(new_n1148), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1169), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1150), .A2(new_n1154), .A3(new_n1160), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1161), .A2(new_n1145), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT125), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1177), .B(KEYINPUT48), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1174), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1150), .A2(new_n1152), .A3(new_n1160), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n803), .A2(new_n1103), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1146), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1168), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1186));
  OAI21_X1  g760(.A(new_n460), .B1(new_n676), .B2(new_n677), .ZN(new_n1187));
  INV_X1    g761(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n662), .B2(new_n1188), .ZN(new_n1189));
  AOI211_X1 g763(.A(KEYINPUT126), .B(new_n1187), .C1(new_n659), .C2(new_n661), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g765(.A(KEYINPUT127), .B1(new_n714), .B2(new_n1191), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n714), .A2(new_n1191), .A3(KEYINPUT127), .ZN(new_n1193));
  OAI211_X1 g767(.A(new_n956), .B(new_n885), .C1(new_n1192), .C2(new_n1193), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


