//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n209), .B1(new_n215), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n209), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(new_n207), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n203), .A2(G50), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT65), .Z(new_n234));
  AOI211_X1 g0034(.A(new_n223), .B(new_n226), .C1(new_n232), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G58), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT66), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n217), .A2(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G97), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G107), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G116), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g0053(.A(new_n247), .B(new_n253), .Z(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n231), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n230), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G77), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g0061(.A1(new_n261), .A2(new_n211), .B1(new_n207), .B2(G68), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n256), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  XOR2_X1   g0064(.A(KEYINPUT71), .B(KEYINPUT11), .Z(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n207), .A3(G1), .ZN(new_n269));
  AOI211_X1 g0069(.A(KEYINPUT72), .B(KEYINPUT12), .C1(new_n269), .C2(new_n202), .ZN(new_n270));
  INV_X1    g0070(.A(new_n269), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n271), .A2(G68), .A3(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n256), .B1(new_n206), .B2(G20), .ZN(new_n274));
  AOI211_X1 g0074(.A(new_n270), .B(new_n273), .C1(G68), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(new_n267), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n281), .A2(new_n277), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n279), .B1(new_n282), .B2(G238), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  INV_X1    g0084(.A(G1698), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n286), .A2(new_n212), .B1(new_n287), .B2(new_n249), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(KEYINPUT3), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(new_n285), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n288), .B1(G232), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n283), .B1(new_n294), .B2(new_n281), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT14), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G179), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n295), .B(KEYINPUT13), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT14), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n303), .A3(G169), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n276), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n276), .B1(new_n297), .B2(G190), .ZN(new_n307));
  INV_X1    g0107(.A(G200), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(new_n297), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n279), .B1(new_n282), .B2(G244), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n293), .A2(G238), .B1(G107), .B2(new_n292), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n292), .A2(G1698), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G232), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n310), .B1(new_n314), .B2(new_n281), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G200), .ZN(new_n316));
  INV_X1    g0116(.A(new_n256), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT8), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G58), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n230), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n322), .A2(new_n260), .B1(new_n323), .B2(G77), .ZN(new_n324));
  XOR2_X1   g0124(.A(KEYINPUT15), .B(G87), .Z(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G33), .A3(new_n230), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n317), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n274), .A2(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G77), .B2(new_n271), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G190), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n316), .B(new_n330), .C1(new_n331), .C2(new_n315), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n315), .A2(G179), .ZN(new_n333));
  XNOR2_X1  g0133(.A(new_n333), .B(KEYINPUT70), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n330), .B1(new_n315), .B2(new_n298), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n306), .A2(new_n309), .A3(new_n332), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n312), .A2(G222), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n293), .A2(G223), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n338), .B(new_n339), .C1(new_n258), .C2(new_n284), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n280), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n279), .B1(new_n282), .B2(G226), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n343), .A2(new_n331), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(G200), .B2(new_n343), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n274), .A2(G50), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(G50), .B2(new_n271), .ZN(new_n347));
  OAI21_X1  g0147(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n348));
  INV_X1    g0148(.A(G150), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n261), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n319), .B(KEYINPUT69), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT67), .B(G58), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT68), .B1(new_n354), .B2(new_n318), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT68), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n353), .A2(new_n356), .A3(KEYINPUT8), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n352), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n351), .B1(new_n358), .B2(new_n257), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n347), .B1(new_n359), .B2(new_n256), .ZN(new_n360));
  OR2_X1    g0160(.A1(new_n360), .A2(KEYINPUT9), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(KEYINPUT9), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n345), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n363), .B(KEYINPUT10), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n343), .A2(G179), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n298), .B2(new_n343), .ZN(new_n366));
  INV_X1    g0166(.A(new_n360), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n292), .A2(new_n371), .A3(new_n207), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n227), .A2(new_n229), .B1(new_n289), .B2(new_n291), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n372), .B(G68), .C1(new_n373), .C2(new_n371), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n203), .B1(new_n353), .B2(new_n202), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT73), .ZN(new_n378));
  INV_X1    g0178(.A(G159), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n261), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n260), .A2(KEYINPUT73), .A3(G159), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n377), .A2(G20), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n374), .A2(new_n375), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n370), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(KEYINPUT7), .B1(new_n284), .B2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n230), .A2(new_n292), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n386), .B(G68), .C1(new_n387), .C2(KEYINPUT7), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n388), .A2(new_n382), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n317), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n358), .A2(new_n274), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n358), .A2(new_n271), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n385), .A2(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n289), .A2(new_n291), .A3(G226), .A4(G1698), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n289), .A2(new_n291), .A3(G223), .A4(new_n285), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT75), .A4(new_n398), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n402), .A3(new_n280), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n279), .B1(new_n282), .B2(G232), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n331), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n404), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n405), .A2(KEYINPUT76), .B1(new_n406), .B2(new_n308), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n403), .A2(new_n408), .A3(new_n331), .A4(new_n404), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT77), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(KEYINPUT76), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n406), .A2(new_n308), .ZN(new_n412));
  AND4_X1   g0212(.A1(KEYINPUT77), .A2(new_n411), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n393), .B(new_n395), .C1(new_n410), .C2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n385), .A2(new_n390), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n391), .A2(new_n392), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n411), .A2(new_n409), .A3(new_n412), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n407), .A2(KEYINPUT77), .A3(new_n409), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n418), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n414), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n406), .A2(new_n300), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n298), .B1(new_n403), .B2(new_n404), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n393), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT18), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n393), .B2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n424), .A2(new_n432), .ZN(new_n433));
  NOR3_X1   g0233(.A1(new_n337), .A2(new_n369), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n284), .A2(G250), .A3(new_n285), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n284), .A2(G257), .A3(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G294), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT84), .A4(new_n437), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n440), .A2(new_n280), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT5), .B(G41), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n443), .A2(G274), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n445), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n281), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n446), .B1(new_n448), .B2(new_n218), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n442), .A2(new_n331), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT85), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n281), .B1(new_n438), .B2(new_n439), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n449), .B1(new_n454), .B2(new_n441), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(KEYINPUT85), .A3(new_n331), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n442), .A2(new_n450), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n308), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n453), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT25), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n271), .A2(new_n460), .A3(G107), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n271), .B2(G107), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n206), .A2(G33), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n271), .A2(new_n317), .A3(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n462), .A2(new_n463), .B1(G107), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G116), .ZN(new_n468));
  OR2_X1    g0268(.A1(KEYINPUT23), .A2(G107), .ZN(new_n469));
  OAI221_X1 g0269(.A(new_n467), .B1(G20), .B2(new_n468), .C1(new_n230), .C2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n230), .A2(new_n284), .A3(G87), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT22), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT22), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n230), .A2(new_n284), .A3(new_n473), .A4(G87), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n470), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(KEYINPUT24), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n256), .B1(new_n475), .B2(KEYINPUT24), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n459), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n271), .A2(G97), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n481), .B1(new_n465), .B2(G97), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n251), .B2(KEYINPUT6), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n484), .A2(new_n323), .B1(G77), .B2(new_n260), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n372), .B(G107), .C1(new_n373), .C2(new_n371), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT79), .B1(new_n487), .B2(new_n256), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT79), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n317), .C1(new_n485), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n482), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n312), .A2(G244), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n284), .A2(G244), .A3(new_n285), .ZN(new_n496));
  INV_X1    g0296(.A(new_n494), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n492), .A2(new_n493), .B1(G33), .B2(G283), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n495), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n280), .B1(new_n445), .B2(new_n443), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n501), .A2(new_n280), .B1(G257), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n300), .A3(new_n446), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n499), .B(new_n500), .C1(new_n496), .C2(new_n497), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n494), .B1(new_n312), .B2(G244), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n280), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(G257), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n446), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n298), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n491), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n488), .A2(new_n490), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n503), .A2(G190), .A3(new_n446), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n509), .A2(G200), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n482), .A4(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n271), .A2(new_n325), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n230), .A2(new_n284), .A3(G68), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n213), .A2(new_n249), .A3(new_n217), .ZN(new_n518));
  AND3_X1   g0318(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n323), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n257), .A2(new_n249), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n517), .B(new_n520), .C1(new_n521), .C2(KEYINPUT19), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n516), .B1(new_n522), .B2(new_n256), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n465), .A2(new_n325), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n445), .A2(new_n214), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n281), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n445), .A2(G274), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n289), .A2(new_n291), .A3(G238), .A4(new_n285), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT81), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT81), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n284), .A2(new_n532), .A3(G238), .A4(new_n285), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n289), .A2(new_n291), .A3(G244), .A4(G1698), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n468), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n529), .B1(new_n538), .B2(new_n280), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n300), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n536), .B1(new_n533), .B2(new_n531), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n528), .B(new_n527), .C1(new_n541), .C2(new_n281), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n298), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n525), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n542), .B2(new_n331), .ZN(new_n546));
  AND4_X1   g0346(.A1(G87), .A2(new_n317), .A3(new_n271), .A4(new_n464), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n516), .B(new_n547), .C1(new_n522), .C2(new_n256), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n539), .A2(KEYINPUT82), .A3(G190), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n542), .A2(G200), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n546), .A2(new_n548), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  AND4_X1   g0351(.A1(new_n511), .A2(new_n515), .A3(new_n544), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n455), .A2(new_n300), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n457), .A2(new_n298), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n478), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n255), .A2(new_n231), .B1(G20), .B2(new_n219), .ZN(new_n556));
  NAND2_X1  g0356(.A1(G33), .A2(G283), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n249), .B2(G33), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n323), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(KEYINPUT20), .B(new_n556), .C1(new_n323), .C2(new_n558), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n271), .A2(G116), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n465), .B2(G116), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n289), .A2(new_n291), .A3(G257), .A4(new_n285), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT83), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT83), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n284), .A2(new_n569), .A3(G257), .A4(new_n285), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n284), .A2(G264), .A3(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n292), .A2(G303), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n568), .A2(new_n570), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n280), .ZN(new_n574));
  INV_X1    g0374(.A(new_n446), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n502), .B2(G270), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n566), .A2(new_n577), .A3(G169), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n574), .A2(new_n576), .A3(G179), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n566), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n566), .A2(new_n577), .A3(KEYINPUT21), .A4(G169), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(new_n566), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n574), .A2(new_n576), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n585), .B1(new_n586), .B2(new_n308), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n577), .A2(new_n331), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n555), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  AND4_X1   g0390(.A1(new_n434), .A2(new_n480), .A3(new_n552), .A4(new_n590), .ZN(G372));
  INV_X1    g0391(.A(new_n306), .ZN(new_n592));
  INV_X1    g0392(.A(new_n336), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n424), .B(new_n309), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n432), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(new_n364), .B1(new_n367), .B2(new_n366), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n551), .A2(new_n544), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n597), .A2(new_n480), .A3(new_n511), .A4(new_n515), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n555), .A2(new_n584), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n544), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT26), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n551), .A2(new_n544), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(new_n511), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n491), .A2(new_n504), .A3(new_n510), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n605), .A2(KEYINPUT26), .A3(new_n544), .A4(new_n551), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n434), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n596), .A2(new_n609), .ZN(G369));
  NOR2_X1   g0410(.A1(new_n323), .A2(new_n268), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n206), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT27), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n614), .A3(new_n206), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(G213), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT86), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G343), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n555), .ZN(new_n623));
  INV_X1    g0423(.A(G343), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n566), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(new_n584), .ZN(new_n627));
  INV_X1    g0427(.A(G330), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n627), .A2(new_n628), .A3(new_n589), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n622), .A2(new_n584), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n480), .B1(new_n622), .B2(new_n479), .ZN(new_n632));
  INV_X1    g0432(.A(new_n555), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n623), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n623), .B1(new_n631), .B2(new_n636), .ZN(G399));
  INV_X1    g0437(.A(G41), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n224), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n518), .A2(G116), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G1), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n234), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(new_n639), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n643), .B(KEYINPUT28), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n625), .B1(new_n601), .B2(new_n607), .ZN(new_n645));
  OR3_X1    g0445(.A1(new_n645), .A2(KEYINPUT90), .A3(KEYINPUT29), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT90), .B1(new_n645), .B2(KEYINPUT29), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n607), .A2(KEYINPUT91), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n597), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n605), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n649), .B(new_n544), .C1(new_n598), .C2(new_n599), .ZN(new_n650));
  OAI211_X1 g0450(.A(KEYINPUT29), .B(new_n622), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n646), .A2(new_n647), .A3(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n552), .A2(new_n590), .A3(new_n480), .A4(new_n622), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n581), .A2(new_n503), .A3(new_n455), .A4(new_n539), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT87), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT30), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n507), .A2(new_n508), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n542), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n658), .A2(KEYINPUT87), .A3(new_n455), .A4(new_n581), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n586), .A2(new_n539), .A3(G179), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n455), .B1(new_n446), .B2(new_n503), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n656), .A2(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT30), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n654), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n622), .B1(new_n662), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n653), .B1(new_n666), .B2(KEYINPUT31), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n625), .A2(KEYINPUT31), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n654), .A2(new_n655), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n669), .A2(new_n659), .A3(new_n663), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n661), .A2(new_n660), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n664), .B1(new_n672), .B2(KEYINPUT88), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n662), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n668), .B1(new_n673), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(G330), .B1(new_n667), .B2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n625), .B1(new_n672), .B2(new_n664), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT31), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n665), .B1(new_n662), .B2(new_n674), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n672), .A2(KEYINPUT88), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI211_X1 g0485(.A(new_n682), .B(new_n653), .C1(new_n685), .C2(new_n668), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT89), .B1(new_n686), .B2(G330), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n679), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n652), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n644), .B1(new_n690), .B2(G1), .ZN(G364));
  INV_X1    g0491(.A(G311), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n230), .A2(new_n300), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n331), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G200), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n308), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  XOR2_X1   g0498(.A(KEYINPUT33), .B(G317), .Z(new_n699));
  OAI22_X1  g0499(.A1(new_n692), .A2(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G303), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n308), .A2(G179), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(G20), .A3(G190), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n331), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n300), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n323), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G294), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n292), .B1(new_n701), .B2(new_n703), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n693), .A2(new_n704), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n709), .B1(G322), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G283), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n323), .A2(new_n331), .A3(new_n702), .ZN(new_n714));
  INV_X1    g0514(.A(G326), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n693), .A2(G190), .A3(G200), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n712), .B1(new_n713), .B2(new_n714), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  NOR4_X1   g0517(.A1(new_n230), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n700), .B(new_n717), .C1(G329), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n721), .A2(new_n379), .ZN(new_n724));
  XNOR2_X1  g0524(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(KEYINPUT32), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n707), .A2(new_n249), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n714), .A2(new_n217), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n703), .A2(new_n213), .ZN(new_n729));
  OR4_X1    g0529(.A1(new_n292), .A2(new_n727), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n716), .A2(new_n211), .B1(new_n710), .B2(new_n353), .ZN(new_n731));
  OAI22_X1  g0531(.A1(new_n202), .A2(new_n698), .B1(new_n696), .B2(new_n258), .ZN(new_n732));
  NOR4_X1   g0532(.A1(new_n726), .A2(new_n730), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n725), .A2(KEYINPUT32), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n723), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n231), .B1(G20), .B2(new_n298), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n206), .B1(new_n611), .B2(G45), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n639), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n224), .A2(new_n284), .ZN(new_n745));
  INV_X1    g0545(.A(G355), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n745), .A2(new_n746), .B1(G116), .B2(new_n224), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n224), .A2(new_n292), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT93), .Z(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n444), .B2(new_n234), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n247), .A2(G45), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n736), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n744), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n738), .A2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT96), .Z(new_n761));
  OAI21_X1  g0561(.A(new_n756), .B1(new_n627), .B2(new_n589), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n628), .B1(new_n627), .B2(new_n589), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n629), .A2(new_n742), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(G396));
  NAND2_X1  g0566(.A1(new_n593), .A2(new_n622), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n332), .B1(new_n622), .B2(new_n330), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n336), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n688), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n677), .A2(new_n678), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n686), .A2(KEYINPUT89), .A3(G330), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n645), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n742), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n771), .A2(new_n645), .A3(new_n775), .ZN(new_n778));
  AND2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n736), .A2(new_n754), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n744), .B1(G77), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n770), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n755), .ZN(new_n784));
  INV_X1    g0584(.A(new_n716), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G283), .A2(new_n697), .B1(new_n785), .B2(G303), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n219), .B2(new_n696), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT97), .Z(new_n788));
  OAI22_X1  g0588(.A1(new_n721), .A2(new_n692), .B1(new_n213), .B2(new_n714), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT98), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n292), .B1(new_n703), .B2(new_n217), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n793), .B(new_n727), .C1(G294), .C2(new_n711), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n791), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n785), .A2(G137), .B1(new_n711), .B2(G143), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n698), .B2(new_n349), .C1(new_n379), .C2(new_n696), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n714), .A2(new_n202), .B1(new_n211), .B2(new_n703), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT99), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n292), .B1(new_n706), .B2(new_n354), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n722), .A2(G132), .B1(new_n801), .B2(new_n800), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n799), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n797), .A2(new_n798), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n788), .A2(new_n795), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n782), .B(new_n784), .C1(new_n736), .C2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n779), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G384));
  INV_X1    g0610(.A(KEYINPUT38), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n390), .B1(KEYINPUT16), .B2(new_n389), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(new_n417), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n621), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n424), .B2(new_n432), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n393), .B1(new_n410), .B2(new_n413), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n620), .A2(new_n427), .B1(new_n812), .B2(new_n417), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n620), .A2(new_n427), .B1(new_n416), .B2(new_n417), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n423), .A2(KEYINPUT37), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n811), .B1(new_n815), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n821), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n817), .A2(new_n825), .A3(new_n816), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT37), .B1(new_n423), .B2(new_n818), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n415), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n817), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n830), .A2(new_n414), .B1(new_n431), .B2(new_n429), .ZN(new_n831));
  OAI211_X1 g0631(.A(KEYINPUT38), .B(new_n828), .C1(new_n831), .C2(new_n814), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n824), .A2(KEYINPUT101), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n815), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT101), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT38), .A4(new_n828), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n833), .A2(KEYINPUT39), .A3(new_n836), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n393), .B(new_n620), .C1(new_n424), .C2(new_n432), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n816), .B1(new_n817), .B2(new_n825), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n822), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n811), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT39), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n832), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n837), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n592), .A2(new_n622), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n833), .A2(new_n836), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n604), .A2(new_n606), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n622), .B(new_n769), .C1(new_n600), .C2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n767), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n625), .A2(new_n276), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n306), .A2(new_n309), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n276), .B(new_n625), .C1(new_n302), .C2(new_n305), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n848), .A2(new_n856), .B1(new_n432), .B2(new_n621), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n847), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n646), .A2(new_n647), .A3(new_n434), .A4(new_n651), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n596), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n858), .B(new_n860), .Z(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n680), .A2(new_n862), .A3(new_n681), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n666), .B1(KEYINPUT102), .B2(KEYINPUT31), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n653), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n855), .A2(new_n865), .A3(new_n783), .ZN(new_n866));
  NOR3_X1   g0666(.A1(new_n848), .A2(KEYINPUT40), .A3(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT40), .ZN(new_n868));
  INV_X1    g0668(.A(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n841), .A2(new_n832), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n434), .A3(new_n865), .ZN(new_n873));
  OAI21_X1  g0673(.A(G330), .B1(new_n867), .B2(new_n871), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n434), .A2(G330), .A3(new_n865), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n861), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n861), .A2(new_n877), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n878), .B(new_n879), .C1(new_n206), .C2(new_n611), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n484), .A2(KEYINPUT35), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(G116), .A3(new_n232), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(KEYINPUT35), .B2(new_n484), .ZN(new_n883));
  XOR2_X1   g0683(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n884));
  OR2_X1    g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(G77), .B1(new_n353), .B2(new_n202), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n642), .A2(new_n886), .B1(G50), .B2(new_n202), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(G1), .A3(new_n268), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n884), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n880), .A2(new_n885), .A3(new_n888), .A4(new_n889), .ZN(G367));
  OR2_X1    g0690(.A1(new_n622), .A2(new_n548), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(new_n544), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n597), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n756), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n714), .A2(new_n249), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n284), .B(new_n897), .C1(new_n722), .C2(G317), .ZN(new_n898));
  OR2_X1    g0698(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n900));
  OAI22_X1  g0700(.A1(new_n713), .A2(new_n696), .B1(new_n698), .B2(new_n708), .ZN(new_n901));
  INV_X1    g0701(.A(new_n703), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(KEYINPUT46), .A3(G116), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT46), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n703), .B2(new_n219), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n903), .B(new_n905), .C1(new_n707), .C2(new_n217), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n716), .A2(new_n692), .B1(new_n710), .B2(new_n701), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n901), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n899), .A2(new_n900), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(G137), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n721), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n284), .B1(new_n703), .B2(new_n353), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n714), .A2(new_n258), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n912), .B(new_n913), .C1(G68), .C2(new_n706), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n785), .A2(G143), .B1(new_n711), .B2(G150), .ZN(new_n915));
  AOI22_X1  g0715(.A1(G50), .A2(new_n695), .B1(new_n697), .B2(G159), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n909), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT47), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n737), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n325), .ZN(new_n923));
  OAI221_X1 g0723(.A(new_n757), .B1(new_n224), .B2(new_n923), .C1(new_n750), .C2(new_n242), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n896), .A2(new_n744), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n631), .B(new_n636), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n689), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n635), .A2(new_n630), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n625), .A2(new_n491), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n511), .A3(new_n515), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n625), .A2(new_n605), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n928), .A2(new_n623), .A3(new_n932), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT45), .Z(new_n934));
  AOI21_X1  g0734(.A(new_n932), .B1(new_n928), .B2(new_n623), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT44), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n629), .A2(new_n635), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n927), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n690), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n639), .B(KEYINPUT41), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n740), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n635), .A2(new_n630), .A3(new_n932), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n511), .B1(new_n930), .B2(new_n633), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT103), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n625), .B1(new_n946), .B2(KEYINPUT103), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n944), .A2(KEYINPUT42), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n945), .A2(new_n949), .B1(KEYINPUT43), .B2(new_n894), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n894), .A2(KEYINPUT43), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n950), .B(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n932), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n938), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n952), .B(new_n954), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n925), .B1(new_n943), .B2(new_n955), .ZN(G387));
  NOR2_X1   g0756(.A1(new_n926), .A2(new_n739), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n745), .A2(new_n640), .B1(G107), .B2(new_n224), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n959));
  NAND3_X1  g0759(.A1(new_n322), .A2(new_n959), .A3(new_n211), .ZN(new_n960));
  INV_X1    g0760(.A(new_n959), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n321), .B2(G50), .ZN(new_n962));
  AOI21_X1  g0762(.A(G45), .B1(G68), .B2(G77), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n960), .A2(new_n962), .A3(new_n640), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT106), .B1(new_n749), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G45), .B2(new_n239), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n749), .A2(KEYINPUT106), .A3(new_n964), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n958), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n358), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n969), .A2(new_n697), .B1(new_n695), .B2(G68), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT107), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n721), .A2(new_n349), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n706), .A2(new_n325), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n902), .A2(G77), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n284), .A3(new_n976), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n716), .A2(new_n379), .B1(new_n710), .B2(new_n211), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n974), .A2(new_n897), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n972), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n785), .A2(G322), .B1(new_n711), .B2(G317), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n698), .B2(new_n692), .C1(new_n701), .C2(new_n696), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT48), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n983), .B1(new_n713), .B2(new_n707), .C1(new_n708), .C2(new_n703), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n292), .B1(new_n219), .B2(new_n714), .C1(new_n721), .C2(new_n715), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n985), .B2(new_n986), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n980), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n744), .B1(new_n758), .B2(new_n968), .C1(new_n990), .C2(new_n737), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT109), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n636), .A2(new_n756), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n957), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n927), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(KEYINPUT110), .A3(new_n741), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n689), .A2(new_n926), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT110), .B1(new_n995), .B2(new_n741), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n994), .B1(new_n998), .B2(new_n999), .ZN(G393));
  XNOR2_X1  g0800(.A(new_n937), .B(new_n938), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n741), .B(new_n940), .C1(new_n1001), .C2(new_n927), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n953), .A2(new_n756), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n757), .B1(new_n249), .B2(new_n224), .C1(new_n750), .C2(new_n253), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT111), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n743), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n1005), .B2(new_n1004), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n284), .B(new_n728), .C1(G283), .C2(new_n902), .ZN(new_n1008));
  INV_X1    g0808(.A(G322), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n1009), .B2(new_n721), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT114), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n785), .A2(G317), .B1(new_n711), .B2(G311), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT52), .Z(new_n1013));
  OAI22_X1  g0813(.A1(new_n698), .A2(new_n701), .B1(new_n219), .B2(new_n707), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(G294), .B2(new_n695), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1010), .A2(KEYINPUT114), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n292), .B1(new_n902), .B2(G68), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n213), .B2(new_n714), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n722), .B2(G143), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT112), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n716), .A2(new_n349), .B1(new_n710), .B2(new_n379), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT51), .Z(new_n1024));
  NOR2_X1   g0824(.A1(new_n707), .A2(new_n258), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n322), .B2(new_n695), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n211), .B2(new_n698), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1022), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1018), .B1(new_n1029), .B2(KEYINPUT113), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT113), .B2(new_n1029), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1007), .B1(new_n1031), .B2(new_n736), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1001), .A2(new_n740), .B1(new_n1003), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1002), .A2(new_n1033), .ZN(G390));
  NAND2_X1  g0834(.A1(new_n856), .A2(new_n846), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n837), .A2(new_n843), .A3(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n783), .B(new_n855), .C1(new_n679), .C2(new_n687), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n622), .B(new_n769), .C1(new_n648), .C2(new_n650), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n767), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n855), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n870), .A2(new_n1040), .A3(new_n846), .ZN(new_n1041));
  AND3_X1   g0841(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n869), .A2(G330), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT115), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1036), .A2(new_n1037), .A3(new_n1041), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT115), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n859), .A2(new_n596), .A3(new_n875), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1043), .B1(new_n774), .B2(new_n855), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n851), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n865), .A2(G330), .A3(new_n783), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n855), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1039), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1037), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1050), .B1(new_n1052), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(KEYINPUT117), .B1(new_n1049), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1059), .A2(new_n639), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1045), .A2(new_n1048), .A3(new_n1057), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT116), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n1045), .A2(new_n1057), .A3(KEYINPUT116), .A4(new_n1048), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1049), .A2(KEYINPUT117), .A3(new_n1058), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1049), .A2(new_n739), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n845), .A2(new_n754), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n744), .B1(new_n969), .B2(new_n781), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n722), .A2(G294), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G97), .A2(new_n695), .B1(new_n697), .B2(G107), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n714), .A2(new_n202), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1025), .A2(new_n1073), .A3(new_n284), .A4(new_n729), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n785), .A2(G283), .B1(new_n711), .B2(G116), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n722), .A2(G125), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT54), .B(G143), .Z(new_n1078));
  AOI22_X1  g0878(.A1(G137), .A2(new_n697), .B1(new_n695), .B2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n703), .A2(new_n349), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1081));
  OAI22_X1  g0881(.A1(new_n707), .A2(new_n379), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n785), .A2(G128), .B1(new_n711), .B2(G132), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1077), .A2(new_n1079), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n284), .B1(new_n714), .B2(new_n211), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT118), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1076), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1070), .B1(new_n1088), .B2(new_n736), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1068), .B1(new_n1069), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1067), .A2(new_n1090), .ZN(G378));
  INV_X1    g0891(.A(new_n1050), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1065), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n364), .A2(KEYINPUT120), .A3(new_n368), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT120), .B1(new_n364), .B2(new_n368), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n620), .A2(new_n360), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1099));
  AND3_X1   g0899(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1098), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n874), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n874), .A2(new_n1102), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n1104), .A2(new_n1105), .B1(new_n847), .B2(new_n857), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1105), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n858), .A3(new_n1103), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1093), .A2(KEYINPUT57), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT57), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1050), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1110), .A2(new_n741), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n754), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n742), .B1(G50), .B2(new_n781), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n287), .A2(new_n638), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n211), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n638), .B2(new_n292), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n714), .A2(new_n353), .ZN(new_n1121));
  AOI211_X1 g0921(.A(G41), .B(new_n284), .C1(new_n902), .C2(G77), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n202), .B2(new_n707), .C1(new_n217), .C2(new_n710), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n1121), .B(new_n1123), .C1(G116), .C2(new_n785), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G97), .A2(new_n697), .B1(new_n695), .B2(new_n325), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n713), .C2(new_n721), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT58), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1120), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n902), .A2(new_n1078), .ZN(new_n1129));
  INV_X1    g0929(.A(G128), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1129), .B1(new_n710), .B2(new_n1130), .C1(new_n349), .C2(new_n707), .ZN(new_n1131));
  INV_X1    g0931(.A(G132), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n1132), .A2(new_n698), .B1(new_n696), .B2(new_n910), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(G125), .C2(new_n785), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(KEYINPUT59), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n722), .A2(G124), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n714), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1138), .B2(G159), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT59), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1137), .B(new_n1139), .C1(new_n1134), .C2(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1128), .B1(new_n1127), .B2(new_n1126), .C1(new_n1136), .C2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1117), .B1(new_n1142), .B2(new_n736), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1109), .A2(new_n740), .B1(new_n1116), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1115), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT121), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT121), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1115), .A2(new_n1147), .A3(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(G375));
  NAND2_X1  g0949(.A1(new_n697), .A2(new_n1078), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n696), .B2(new_n349), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n284), .B1(new_n703), .B2(new_n379), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1152), .B(new_n1121), .C1(G50), .C2(new_n706), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n1132), .B2(new_n716), .C1(new_n910), .C2(new_n710), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1151), .B(new_n1154), .C1(G128), .C2(new_n722), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n975), .B1(new_n710), .B2(new_n713), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT123), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n721), .A2(new_n701), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n284), .B(new_n913), .C1(G97), .C2(new_n902), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G107), .A2(new_n695), .B1(new_n697), .B2(G116), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n708), .C2(new_n716), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1158), .B(new_n1161), .C1(new_n1157), .C2(new_n1156), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n736), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n743), .B1(new_n202), .B2(new_n780), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n855), .C2(new_n755), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1052), .A2(new_n1056), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n739), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1050), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT122), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1058), .A2(new_n942), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(G381));
  INV_X1    g0972(.A(G378), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1146), .A2(new_n1173), .A3(new_n1148), .ZN(new_n1174));
  OR2_X1    g0974(.A1(G387), .A2(G390), .ZN(new_n1175));
  OR2_X1    g0975(.A1(G393), .A2(G396), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(G384), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT124), .ZN(new_n1178));
  OR4_X1    g0978(.A1(G381), .A2(new_n1174), .A3(new_n1175), .A4(new_n1178), .ZN(G407));
  INV_X1    g0979(.A(new_n1148), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1147), .B1(new_n1115), .B2(new_n1144), .ZN(new_n1181));
  NOR3_X1   g0981(.A1(new_n1180), .A2(new_n1181), .A3(G378), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n624), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(G407), .A2(G213), .A3(new_n1183), .ZN(G409));
  NAND2_X1  g0984(.A1(new_n1145), .A2(G378), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1067), .A2(new_n1144), .A3(new_n1090), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1093), .A2(new_n942), .A3(new_n1109), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1186), .A2(new_n1187), .B1(G213), .B2(new_n624), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT60), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n741), .B1(new_n1169), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT122), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1169), .B(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1057), .A2(new_n1190), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1191), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n809), .B1(new_n1196), .B2(new_n1167), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1170), .A2(new_n1194), .ZN(new_n1198));
  OAI211_X1 g0998(.A(G384), .B(new_n1168), .C1(new_n1198), .C2(new_n1191), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n624), .A2(G213), .A3(G2897), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1200), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT61), .B1(new_n1189), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1185), .A2(new_n1188), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT63), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(G387), .B(G390), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT125), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(G393), .B(G396), .ZN(new_n1212));
  OR3_X1    g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1214));
  INV_X1    g1014(.A(G390), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT126), .ZN(new_n1216));
  OR3_X1    g1016(.A1(new_n1215), .A2(G387), .A3(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(G387), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1215), .B2(G387), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1217), .A2(new_n1212), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1213), .A2(new_n1214), .A3(new_n1220), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1185), .A2(KEYINPUT63), .A3(new_n1188), .A4(new_n1206), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1204), .A2(new_n1209), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT62), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1185), .A2(new_n1224), .A3(new_n1188), .A4(new_n1206), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1207), .A2(KEYINPUT62), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1204), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1223), .B1(new_n1227), .B2(new_n1221), .ZN(G405));
  INV_X1    g1028(.A(KEYINPUT127), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1221), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1221), .A2(new_n1229), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1174), .A2(new_n1185), .A3(new_n1206), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1206), .B1(new_n1174), .B2(new_n1185), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1230), .B(new_n1231), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1185), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1205), .B1(new_n1182), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1174), .A2(new_n1185), .A3(new_n1206), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1236), .A2(new_n1229), .A3(new_n1221), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(G402));
endmodule


