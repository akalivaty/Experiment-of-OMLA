//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n560,
    new_n561, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT67), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n453), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  INV_X1    g034(.A(new_n455), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G125), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .B1(G113), .B2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n471), .B1(new_n478), .B2(G2105), .ZN(G160));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n473), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT69), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n480), .A2(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT70), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n467), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT70), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  OR2_X1    g065(.A1(G100), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n483), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n468), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n486), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n472), .B2(new_n473), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n501), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT71), .B1(new_n501), .B2(KEYINPUT4), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n500), .B(new_n505), .C1(new_n473), .C2(new_n472), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n467), .A2(KEYINPUT72), .A3(new_n505), .A4(new_n500), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n498), .B1(new_n504), .B2(new_n510), .ZN(G164));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT73), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n512), .A2(new_n513), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT5), .B(G543), .Z(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n525), .A2(new_n518), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(G651), .B1(new_n528), .B2(G88), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n523), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n515), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n514), .A2(G89), .ZN(new_n536));
  NAND2_X1  g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n525), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g113(.A1(new_n535), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  XNOR2_X1  g115(.A(KEYINPUT5), .B(G543), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(KEYINPUT74), .B(G52), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n520), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT75), .B(G90), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n528), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n514), .A2(new_n541), .ZN(new_n552));
  INV_X1    g127(.A(G81), .ZN(new_n553));
  OAI22_X1  g128(.A1(new_n551), .A2(new_n515), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n541), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n543), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n520), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n525), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n528), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  OR2_X1    g144(.A1(new_n541), .A2(G74), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n570), .A2(G651), .B1(new_n520), .B2(G49), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n528), .A2(G87), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(new_n520), .A2(G48), .ZN(new_n574));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n541), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  OAI221_X1 g151(.A(new_n574), .B1(new_n552), .B2(new_n575), .C1(new_n543), .C2(new_n576), .ZN(G305));
  INV_X1    g152(.A(G47), .ZN(new_n578));
  INV_X1    g153(.A(G85), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n578), .A2(new_n515), .B1(new_n552), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n541), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n528), .A2(G92), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n525), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G284));
  OAI21_X1  g168(.A(new_n585), .B1(new_n592), .B2(G868), .ZN(G321));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  NAND3_X1  g170(.A1(G286), .A2(new_n595), .A3(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(G868), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n595), .B1(G286), .B2(G868), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n596), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G297));
  XNOR2_X1  g177(.A(new_n601), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n592), .B1(new_n604), .B2(G860), .ZN(G148));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n554), .B2(new_n556), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n587), .A2(new_n591), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n609), .B2(new_n606), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n481), .A2(G135), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT79), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n489), .A2(G123), .ZN(new_n615));
  OR2_X1    g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n616), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G2096), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n467), .A2(new_n465), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  NOR2_X1   g199(.A1(KEYINPUT78), .A2(G2100), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n620), .B(new_n626), .C1(new_n624), .C2(new_n621), .ZN(G156));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XOR2_X1   g204(.A(G2443), .B(G2446), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT82), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT83), .Z(G401));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT84), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  XOR2_X1   g228(.A(new_n651), .B(KEYINPUT17), .Z(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n648), .B1(new_n650), .B2(new_n651), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n656), .B1(new_n658), .B2(KEYINPUT85), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(KEYINPUT85), .B2(new_n658), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n619), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT86), .B(G2100), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  INV_X1    g259(.A(KEYINPUT36), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G24), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(new_n583), .B2(new_n686), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(G1986), .Z(new_n689));
  NOR2_X1   g264(.A1(G25), .A2(G29), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT35), .B(G1991), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n485), .A2(G119), .A3(new_n488), .ZN(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n695));
  INV_X1    g270(.A(G107), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G2105), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n481), .B2(G131), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n694), .A2(KEYINPUT87), .A3(new_n698), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n691), .B(new_n693), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n691), .B1(new_n703), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(new_n692), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n689), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT88), .B(KEYINPUT34), .Z(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G1976), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n686), .B1(new_n571), .B2(new_n572), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n686), .A2(G23), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT33), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n712), .A2(KEYINPUT33), .A3(new_n714), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(new_n717), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n719), .A2(G1976), .A3(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n686), .A2(G22), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT90), .Z(new_n724));
  OAI211_X1 g299(.A(new_n722), .B(new_n724), .C1(G166), .C2(new_n686), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n686), .A2(G6), .ZN(new_n726));
  INV_X1    g301(.A(G48), .ZN(new_n727));
  OAI22_X1  g302(.A1(new_n727), .A2(new_n515), .B1(new_n552), .B2(new_n575), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n576), .A2(new_n543), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n726), .B1(new_n730), .B2(new_n686), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT32), .B(G1981), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT89), .Z(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n686), .B1(new_n523), .B2(new_n529), .ZN(new_n736));
  INV_X1    g311(.A(new_n724), .ZN(new_n737));
  OAI21_X1  g312(.A(G1971), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n726), .B(new_n733), .C1(new_n730), .C2(new_n686), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n725), .A2(new_n735), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n710), .B1(new_n721), .B2(new_n740), .ZN(new_n741));
  AND4_X1   g316(.A1(new_n725), .A2(new_n735), .A3(new_n738), .A4(new_n739), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n742), .A2(new_n709), .A3(new_n720), .A4(new_n718), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n708), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n685), .B1(new_n744), .B2(KEYINPUT91), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT91), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n741), .A2(new_n708), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(KEYINPUT92), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n745), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n741), .A2(new_n708), .A3(new_n743), .A4(new_n685), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n686), .A2(G4), .ZN(new_n755));
  OAI211_X1 g330(.A(G1348), .B(new_n755), .C1(new_n592), .C2(new_n686), .ZN(new_n756));
  INV_X1    g331(.A(G1348), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n686), .B1(new_n587), .B2(new_n591), .ZN(new_n758));
  INV_X1    g333(.A(new_n755), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n618), .A2(new_n704), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n557), .A2(G16), .ZN(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n763), .A2(G1341), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT31), .B(G11), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT97), .ZN(new_n768));
  INV_X1    g343(.A(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n769), .B2(KEYINPUT30), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(G286), .A2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n686), .A2(G21), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  AND4_X1   g351(.A1(new_n762), .A2(new_n766), .A3(new_n772), .A4(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n704), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n489), .A2(G129), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n465), .A2(G105), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT26), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n780), .B(new_n782), .C1(G141), .C2(new_n481), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n778), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n686), .A2(G5), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G301), .B2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n774), .B1(new_n773), .B2(new_n775), .ZN(new_n792));
  AOI21_X1  g367(.A(G1341), .B1(new_n763), .B2(new_n765), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n761), .A2(new_n777), .A3(new_n787), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n686), .A2(G20), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT23), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G299), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1956), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n789), .A2(new_n790), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT98), .ZN(new_n802));
  NOR2_X1   g377(.A1(G27), .A2(G29), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G164), .B2(G29), .ZN(new_n804));
  INV_X1    g379(.A(G2078), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n800), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n795), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n809));
  INV_X1    g384(.A(G35), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G29), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(new_n493), .B2(G29), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT29), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AOI211_X1 g389(.A(KEYINPUT29), .B(new_n811), .C1(new_n493), .C2(G29), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2090), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI211_X1 g393(.A(KEYINPUT99), .B(G2090), .C1(new_n814), .C2(new_n815), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n814), .A2(new_n815), .A3(G2090), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n704), .A2(G26), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT28), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n489), .A2(G128), .ZN(new_n825));
  NOR2_X1   g400(.A1(G104), .A2(G2105), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT94), .Z(new_n827));
  INV_X1    g402(.A(G116), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n464), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n827), .A2(new_n829), .B1(new_n481), .B2(G140), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n824), .B1(new_n831), .B2(G29), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G2067), .ZN(new_n833));
  INV_X1    g408(.A(G2067), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n704), .B1(new_n825), .B2(new_n830), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n835), .B2(new_n824), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT24), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n704), .B1(new_n838), .B2(G34), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(G34), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G160), .B2(G29), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(G2084), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n704), .A2(G33), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(G139), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n847), .B2(new_n469), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n467), .A2(G127), .ZN(new_n849));
  NAND2_X1  g424(.A1(G115), .A2(G2104), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n468), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n843), .B1(new_n852), .B2(new_n704), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT95), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(KEYINPUT95), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(G2072), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n841), .A2(G2084), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n837), .A2(new_n842), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(G2072), .B1(new_n854), .B2(new_n855), .ZN(new_n859));
  OR2_X1    g434(.A1(new_n859), .A2(KEYINPUT96), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(KEYINPUT96), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n808), .A2(new_n820), .A3(new_n822), .A4(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI211_X1 g440(.A(new_n821), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n866), .A2(KEYINPUT100), .A3(new_n820), .A4(new_n808), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n754), .A2(new_n868), .ZN(G311));
  NAND2_X1  g444(.A1(new_n753), .A2(new_n751), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n750), .B1(new_n745), .B2(new_n747), .ZN(new_n871));
  OAI211_X1 g446(.A(KEYINPUT101), .B(new_n868), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT101), .B1(new_n754), .B2(new_n868), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(G150));
  XNOR2_X1  g450(.A(KEYINPUT104), .B(G860), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n608), .A2(new_n604), .ZN(new_n878));
  XNOR2_X1  g453(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(G93), .ZN(new_n881));
  XOR2_X1   g456(.A(KEYINPUT103), .B(G55), .Z(new_n882));
  OAI22_X1  g457(.A1(new_n881), .A2(new_n552), .B1(new_n515), .B2(new_n882), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n541), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n884), .A2(new_n543), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n557), .B(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n880), .B(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n877), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(KEYINPUT39), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n886), .A2(new_n876), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(KEYINPUT37), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(G145));
  XNOR2_X1  g468(.A(new_n618), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(G162), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n468), .B2(G118), .ZN(new_n898));
  OAI211_X1 g473(.A(KEYINPUT106), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n899));
  INV_X1    g474(.A(G118), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(KEYINPUT105), .A3(G2105), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI22_X1  g480(.A1(G142), .A2(new_n481), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n485), .A2(new_n488), .ZN(new_n907));
  INV_X1    g482(.A(G130), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n909), .B(KEYINPUT107), .Z(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(new_n623), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT71), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n468), .A2(G138), .ZN(new_n913));
  OR2_X1    g488(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n914));
  NAND2_X1  g489(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n912), .B1(new_n916), .B2(new_n505), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n501), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n508), .A3(new_n509), .A4(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n498), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n852), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n911), .B(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n784), .B(new_n831), .ZN(new_n924));
  INV_X1    g499(.A(new_n703), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n923), .A2(new_n926), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n896), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n923), .A2(new_n926), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n895), .A3(new_n927), .ZN(new_n932));
  INV_X1    g507(.A(G37), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  XOR2_X1   g509(.A(KEYINPUT108), .B(KEYINPUT40), .Z(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(G395));
  XNOR2_X1  g511(.A(new_n609), .B(new_n887), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n608), .A2(G299), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n597), .A2(new_n587), .A3(new_n591), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n940), .B1(new_n938), .B2(new_n939), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n608), .A2(G299), .ZN(new_n945));
  AOI22_X1  g520(.A1(new_n587), .A2(new_n591), .B1(new_n564), .B2(new_n568), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT41), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n947), .A2(KEYINPUT109), .ZN(new_n948));
  OAI211_X1 g523(.A(KEYINPUT110), .B(new_n937), .C1(new_n944), .C2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n949), .B1(new_n937), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n947), .A2(KEYINPUT109), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n942), .A2(new_n943), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n954), .A3(new_n941), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT110), .B1(new_n955), .B2(new_n937), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT112), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n952), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n957), .B1(new_n952), .B2(new_n956), .ZN(new_n959));
  XNOR2_X1  g534(.A(G290), .B(G303), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n730), .B(G288), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n963), .B(KEYINPUT42), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n958), .B1(new_n959), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n952), .A2(new_n956), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n966), .A2(KEYINPUT112), .A3(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(G868), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n606), .B1(new_n883), .B2(new_n885), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(G295));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n969), .ZN(G331));
  XNOR2_X1  g546(.A(G286), .B(G301), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(new_n887), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n887), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n955), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n962), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(KEYINPUT113), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n972), .A2(new_n887), .A3(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n978), .A2(new_n973), .A3(new_n950), .A4(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n977), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n973), .A3(new_n980), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n947), .A2(new_n941), .A3(KEYINPUT114), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n983), .B(new_n984), .C1(KEYINPUT114), .C2(new_n947), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n973), .A2(new_n950), .A3(new_n974), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n977), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT115), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n982), .B(new_n933), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  AOI211_X1 g564(.A(KEYINPUT115), .B(new_n977), .C1(new_n985), .C2(new_n986), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NOR3_X1   g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n982), .A2(new_n933), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n976), .A2(new_n981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n962), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT43), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n992), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n989), .A2(new_n990), .A3(KEYINPUT43), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n991), .B1(new_n993), .B2(new_n995), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(G397));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(G164), .B2(G1384), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G160), .A2(G40), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n831), .B(new_n834), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n784), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n925), .A2(new_n692), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n703), .A2(new_n693), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n583), .B(G1986), .Z(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G40), .ZN(new_n1018));
  AOI211_X1 g593(.A(new_n1018), .B(new_n471), .C1(new_n478), .C2(G2105), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1384), .B1(new_n919), .B2(new_n920), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1019), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI211_X1 g597(.A(KEYINPUT50), .B(G1384), .C1(new_n919), .C2(new_n920), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(KEYINPUT45), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1004), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n817), .A2(new_n1024), .B1(new_n1026), .B2(new_n722), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1017), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT49), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n730), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(G305), .A2(G1981), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1030), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n730), .A2(new_n1031), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G305), .A2(G1981), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1034), .A2(G8), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n571), .A2(G1976), .A3(new_n572), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT52), .B1(G288), .B2(new_n711), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1035), .A2(G8), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1035), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1045), .A2(new_n1028), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1044), .B1(new_n1046), .B2(new_n1040), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1017), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1020), .A2(KEYINPUT45), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1003), .B(G1384), .C1(new_n919), .C2(new_n920), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1050), .A2(new_n1051), .A3(new_n1005), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(G1971), .ZN(new_n1053));
  INV_X1    g628(.A(G1384), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n921), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1019), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(G2090), .ZN(new_n1059));
  OAI211_X1 g634(.A(G8), .B(new_n1049), .C1(new_n1053), .C2(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1029), .A2(new_n1048), .A3(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1022), .A2(new_n1023), .A3(G2084), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1026), .A2(new_n774), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1028), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1061), .A2(G168), .A3(new_n1065), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1029), .A2(new_n1048), .A3(new_n1060), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1065), .A2(G168), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1066), .B(new_n1067), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(KEYINPUT118), .A2(KEYINPUT63), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1046), .B(KEYINPUT117), .ZN(new_n1075));
  NOR2_X1   g650(.A1(G288), .A2(G1976), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1033), .B1(new_n1039), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1060), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1078), .B1(new_n1079), .B2(new_n1048), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n1081));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n568), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G299), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n564), .B(new_n568), .C1(new_n1081), .C2(KEYINPUT57), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1004), .A2(new_n1019), .A3(new_n1025), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1087), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n757), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1045), .A2(new_n834), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n608), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n608), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1096), .A2(new_n1097), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n592), .A2(KEYINPUT60), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1096), .A2(new_n1097), .A3(KEYINPUT60), .A4(new_n592), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT61), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1085), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1094), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n557), .A2(KEYINPUT122), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1004), .A2(new_n1008), .A3(new_n1019), .A4(new_n1025), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  NAND2_X1  g689(.A1(new_n1035), .A2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1113), .A2(KEYINPUT121), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT121), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1112), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(KEYINPUT59), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1120), .B(new_n1112), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1111), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1093), .A2(KEYINPUT61), .A3(new_n1095), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1100), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT54), .B1(G301), .B2(KEYINPUT125), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1026), .B2(G2078), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n805), .A2(KEYINPUT53), .ZN(new_n1130));
  OAI22_X1  g705(.A1(new_n1024), .A2(G1961), .B1(new_n1026), .B2(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1129), .A2(new_n1131), .A3(G171), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1127), .A2(G2078), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n1052), .A2(new_n1133), .B1(new_n1058), .B2(new_n790), .ZN(new_n1134));
  AOI21_X1  g709(.A(G301), .B1(new_n1134), .B2(new_n1128), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1126), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(G171), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(G301), .A3(new_n1128), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n1138), .A3(new_n1125), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1070), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  INV_X1    g716(.A(G2084), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1142), .A2(new_n1024), .B1(new_n1026), .B2(new_n774), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1141), .B1(new_n1143), .B2(new_n1028), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1966), .B1(new_n1145), .B2(new_n1019), .ZN(new_n1146));
  OAI211_X1 g721(.A(KEYINPUT124), .B(G8), .C1(new_n1146), .C2(new_n1062), .ZN(new_n1147));
  NAND2_X1  g722(.A1(G286), .A2(G8), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT51), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1144), .A2(new_n1147), .A3(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1148), .B(KEYINPUT123), .Z(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1143), .B2(new_n1028), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT51), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1143), .A2(new_n1148), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1140), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1074), .B(new_n1080), .C1(new_n1124), .C2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1157), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  OAI21_X1  g738(.A(KEYINPUT126), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1135), .A2(new_n1029), .A3(new_n1048), .A4(new_n1060), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1165), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n1167));
  OAI21_X1  g742(.A(G8), .B1(new_n1146), .B2(new_n1062), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1150), .B1(new_n1168), .B2(new_n1141), .ZN(new_n1169));
  AOI22_X1  g744(.A1(new_n1169), .A2(new_n1147), .B1(KEYINPUT51), .B2(new_n1154), .ZN(new_n1170));
  OAI211_X1 g745(.A(new_n1167), .B(KEYINPUT62), .C1(new_n1170), .C2(new_n1157), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1164), .A2(new_n1166), .A3(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1014), .B1(new_n1161), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1174));
  OR2_X1    g749(.A1(new_n1174), .A2(KEYINPUT46), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(KEYINPUT46), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1007), .A2(new_n779), .A3(new_n783), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1175), .A2(new_n1176), .B1(new_n1006), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1178), .B(KEYINPUT47), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n1012), .A2(new_n1006), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1180), .A2(KEYINPUT127), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1180), .A2(KEYINPUT127), .ZN(new_n1182));
  NOR4_X1   g757(.A1(new_n1004), .A2(G1986), .A3(G290), .A4(new_n1005), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  NOR3_X1   g759(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1186), .A2(new_n1010), .B1(G2067), .B2(new_n831), .ZN(new_n1187));
  AOI211_X1 g762(.A(new_n1179), .B(new_n1185), .C1(new_n1006), .C2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1173), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g764(.A1(G401), .A2(new_n462), .ZN(new_n1191));
  AND3_X1   g765(.A1(new_n683), .A2(new_n665), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1192), .B(new_n934), .C1(new_n999), .C2(new_n1000), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


