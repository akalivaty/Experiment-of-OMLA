//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  AOI211_X1 g0013(.A(new_n205), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n214), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(KEYINPUT0), .B2(new_n214), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT65), .B(G244), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n225), .B1(G77), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n209), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n221), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n215), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT71), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G58), .ZN(new_n258));
  OR2_X1    g0058(.A1(KEYINPUT72), .A2(KEYINPUT8), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT72), .A2(KEYINPUT8), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT8), .ZN(new_n262));
  OAI21_X1  g0062(.A(KEYINPUT73), .B1(new_n262), .B2(G58), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT73), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(new_n265), .B2(new_n261), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n207), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT74), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G68), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n223), .A2(new_n258), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G20), .A2(G33), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n272), .A2(G20), .B1(G150), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n257), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT75), .ZN(new_n276));
  OR2_X1    g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n276), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n257), .B1(G1), .B2(new_n207), .ZN(new_n282));
  MUX2_X1   g0082(.A(new_n281), .B(new_n282), .S(G50), .Z(new_n283));
  NAND3_X1  g0083(.A1(new_n277), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT3), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT70), .ZN(new_n290));
  AND3_X1   g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n287), .B2(new_n289), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1698), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n293), .A2(G222), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G77), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n295), .B1(new_n296), .B2(new_n293), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  AOI21_X1  g0105(.A(G1), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n300), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(KEYINPUT69), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n309), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n308), .B1(new_n315), .B2(G226), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n301), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(KEYINPUT76), .B1(new_n285), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT76), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n284), .B(new_n321), .C1(G169), .C2(new_n318), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT77), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT77), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n320), .A2(new_n327), .A3(new_n322), .A4(new_n324), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT78), .ZN(new_n331));
  INV_X1    g0131(.A(new_n273), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n267), .B(KEYINPUT74), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n334), .B1(new_n207), .B2(new_n296), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n255), .ZN(new_n338));
  INV_X1    g0138(.A(new_n255), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n281), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT79), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(G77), .C1(G1), .C2(new_n207), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n279), .A2(new_n207), .A3(G1), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(new_n296), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n315), .A2(new_n226), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n307), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n293), .A2(G232), .A3(new_n294), .ZN(new_n348));
  INV_X1    g0148(.A(G107), .ZN(new_n349));
  INV_X1    g0149(.A(G238), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n348), .B1(new_n349), .B2(new_n293), .C1(new_n297), .C2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n347), .B1(new_n351), .B2(new_n300), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n345), .B1(new_n352), .B2(G169), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT81), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n345), .B(KEYINPUT81), .C1(G169), .C2(new_n352), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(new_n323), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT80), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n352), .A2(KEYINPUT80), .A3(new_n323), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n355), .A2(new_n356), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n352), .A2(G190), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n352), .A2(new_n363), .ZN(new_n364));
  OR3_X1    g0164(.A1(new_n362), .A2(new_n364), .A3(new_n345), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n284), .A2(KEYINPUT9), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT9), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n277), .A2(new_n368), .A3(new_n278), .A4(new_n283), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n317), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(G200), .B2(new_n317), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT10), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n370), .A2(new_n376), .A3(new_n373), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n366), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n288), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT70), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NOR3_X1   g0183(.A1(new_n383), .A2(new_n237), .A3(new_n294), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n381), .A2(G226), .A3(new_n294), .A4(new_n382), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G97), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n300), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n308), .B1(new_n315), .B2(G238), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT13), .ZN(new_n390));
  AND3_X1   g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n390), .B1(new_n388), .B2(new_n389), .ZN(new_n392));
  OAI21_X1  g0192(.A(G200), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n389), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT13), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n395), .A2(G190), .A3(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n335), .A2(new_n296), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n332), .A2(new_n223), .B1(new_n207), .B2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n256), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT11), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n341), .B(G68), .C1(G1), .C2(new_n207), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n343), .A2(new_n271), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n393), .A2(new_n397), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT82), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n393), .A2(new_n397), .A3(new_n408), .A4(KEYINPUT82), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n414), .B(G169), .C1(new_n391), .C2(new_n392), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n395), .A2(new_n396), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n415), .B1(new_n323), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n416), .B2(G169), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n407), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n329), .A2(new_n378), .A3(new_n413), .A4(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(G223), .A2(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n224), .B2(G1698), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT3), .B(G33), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n422), .A2(new_n423), .B1(G33), .B2(G87), .ZN(new_n424));
  OAI221_X1 g0224(.A(new_n307), .B1(new_n424), .B2(new_n309), .C1(new_n237), .C2(new_n314), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(new_n323), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(G169), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT84), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT84), .B1(new_n426), .B2(new_n427), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n266), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n343), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n282), .B2(new_n432), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n258), .A2(new_n271), .ZN(new_n436));
  NOR2_X1   g0236(.A1(G58), .A2(G68), .ZN(new_n437));
  OAI21_X1  g0237(.A(G20), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n273), .A2(G159), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT7), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n423), .B2(G20), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n287), .A2(new_n289), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n440), .B1(new_n445), .B2(G68), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n339), .B1(new_n446), .B2(KEYINPUT16), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT83), .ZN(new_n448));
  AOI21_X1  g0248(.A(G20), .B1(new_n381), .B2(new_n382), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n444), .B1(new_n449), .B2(KEYINPUT7), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n440), .B1(new_n450), .B2(G68), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n447), .B(new_n448), .C1(new_n451), .C2(KEYINPUT16), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n440), .ZN(new_n454));
  INV_X1    g0254(.A(new_n444), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n207), .B1(new_n291), .B2(new_n292), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(new_n441), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(new_n271), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT16), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n448), .B1(new_n460), .B2(new_n447), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n435), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n431), .B(new_n462), .C1(KEYINPUT85), .C2(KEYINPUT18), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n464));
  INV_X1    g0264(.A(new_n430), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n428), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n447), .B1(new_n451), .B2(KEYINPUT16), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT83), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n434), .B1(new_n468), .B2(new_n452), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n464), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT85), .A2(KEYINPUT18), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n463), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n425), .A2(new_n363), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n315), .A2(G232), .ZN(new_n475));
  OR2_X1    g0275(.A1(new_n424), .A2(new_n309), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n475), .A2(new_n476), .A3(new_n371), .A4(new_n307), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n435), .C1(new_n453), .C2(new_n461), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT17), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n469), .A2(KEYINPUT17), .A3(new_n479), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT86), .B1(new_n482), .B2(new_n483), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n473), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n420), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT90), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n305), .A2(G1), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G250), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n488), .B1(new_n491), .B2(new_n300), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n309), .A2(KEYINPUT90), .A3(G250), .A4(new_n490), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n492), .A2(new_n493), .B1(new_n303), .B2(new_n489), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n423), .A2(G244), .ZN(new_n495));
  INV_X1    g0295(.A(G116), .ZN(new_n496));
  OAI22_X1  g0296(.A1(new_n495), .A2(new_n294), .B1(new_n286), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n423), .A2(G238), .A3(new_n294), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT91), .ZN(new_n499));
  OR2_X1    g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n494), .B1(new_n502), .B2(new_n309), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G200), .ZN(new_n504));
  OAI211_X1 g0304(.A(G190), .B(new_n494), .C1(new_n502), .C2(new_n309), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT19), .B1(new_n269), .B2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT19), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n207), .B1(new_n386), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(G87), .B2(new_n203), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n423), .A2(new_n207), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n271), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n255), .B1(new_n506), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n336), .A2(new_n343), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n286), .A2(G1), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n343), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n257), .A2(G87), .A3(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n504), .A2(new_n505), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G169), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n503), .A2(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n323), .B(new_n494), .C1(new_n502), .C2(new_n309), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n257), .A2(new_n515), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n512), .B(new_n513), .C1(new_n336), .C2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n281), .A2(G97), .ZN(new_n526));
  XNOR2_X1  g0326(.A(new_n526), .B(KEYINPUT87), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n527), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n349), .A2(KEYINPUT6), .A3(G97), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n528), .A2(new_n349), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n202), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n532), .B2(KEYINPUT6), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n533), .A2(G20), .B1(G77), .B2(new_n273), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n457), .B2(new_n349), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n529), .B1(new_n255), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  XNOR2_X1  g0337(.A(KEYINPUT5), .B(G41), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n538), .A2(new_n489), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n303), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n489), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n309), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n540), .B1(new_n212), .B2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n381), .A2(G250), .A3(G1698), .A4(new_n382), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT4), .ZN(new_n545));
  INV_X1    g0345(.A(G244), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n381), .A2(new_n294), .A3(new_n382), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n423), .A2(G244), .A3(new_n294), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n545), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G283), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n544), .A2(new_n548), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n543), .B1(new_n552), .B2(new_n300), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n323), .ZN(new_n554));
  INV_X1    g0354(.A(new_n553), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n519), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n537), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(G190), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n559));
  OAI21_X1  g0359(.A(G200), .B1(new_n553), .B2(KEYINPUT88), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n558), .B(new_n536), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT89), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n525), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n557), .A2(new_n561), .A3(KEYINPUT89), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT92), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT92), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n341), .B(G116), .C1(G1), .C2(new_n286), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n551), .B(new_n207), .C1(G33), .C2(new_n528), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n496), .A2(G20), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n255), .A3(new_n572), .ZN(new_n573));
  XOR2_X1   g0373(.A(new_n573), .B(KEYINPUT20), .Z(new_n574));
  INV_X1    g0374(.A(new_n280), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n570), .B(new_n574), .C1(new_n575), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n383), .A2(G303), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n213), .A2(G1698), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n423), .B(new_n578), .C1(G257), .C2(G1698), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n309), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G270), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n540), .B1(new_n581), .B2(new_n542), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n519), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n576), .A2(KEYINPUT21), .A3(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n580), .A2(new_n323), .A3(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n576), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT21), .B1(new_n576), .B2(new_n584), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n583), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n576), .B1(G200), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n371), .B2(new_n591), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G87), .ZN(new_n595));
  OAI21_X1  g0395(.A(KEYINPUT22), .B1(new_n510), .B2(new_n595), .ZN(new_n596));
  OR3_X1    g0396(.A1(new_n595), .A2(KEYINPUT22), .A3(G20), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n383), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n286), .A2(new_n496), .A3(G20), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT23), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(G20), .B2(new_n349), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n207), .A2(KEYINPUT23), .A3(G107), .ZN(new_n603));
  AND2_X1   g0403(.A1(KEYINPUT93), .A2(KEYINPUT24), .ZN(new_n604));
  NOR4_X1   g0404(.A1(new_n600), .A2(new_n602), .A3(new_n603), .A4(new_n604), .ZN(new_n605));
  AND3_X1   g0405(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n599), .B1(new_n598), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n255), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n257), .A2(G107), .A3(new_n515), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n281), .A2(G107), .ZN(new_n610));
  XNOR2_X1  g0410(.A(new_n610), .B(KEYINPUT25), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n608), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(G250), .A2(G1698), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n615), .B1(new_n212), .B2(G1698), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n616), .A2(new_n423), .B1(G33), .B2(G294), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n617), .A2(new_n309), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n541), .A2(G264), .A3(new_n309), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n618), .A2(new_n323), .A3(new_n540), .A4(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n540), .B(new_n619), .C1(new_n309), .C2(new_n617), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n519), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n614), .A2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT94), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n614), .A2(KEYINPUT94), .A3(new_n624), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n621), .A2(new_n371), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(G200), .B2(new_n621), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(new_n608), .A3(new_n613), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT95), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT94), .B1(new_n614), .B2(new_n624), .ZN(new_n634));
  AOI211_X1 g0434(.A(new_n626), .B(new_n623), .C1(new_n608), .C2(new_n613), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT95), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n631), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n594), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n487), .A2(new_n567), .A3(new_n569), .A4(new_n639), .ZN(G372));
  NAND2_X1  g0440(.A1(new_n426), .A2(new_n427), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(KEYINPUT18), .B1(new_n469), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT18), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n462), .A2(new_n644), .A3(new_n641), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n361), .B1(new_n411), .B2(new_n412), .ZN(new_n648));
  INV_X1    g0448(.A(new_n419), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT99), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n482), .A2(new_n483), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT86), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n482), .A2(KEYINPUT86), .A3(new_n483), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n649), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n647), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n375), .A2(new_n377), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(new_n329), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n524), .A2(new_n518), .A3(KEYINPUT96), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT96), .B1(new_n518), .B2(new_n524), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n537), .A2(new_n554), .A3(KEYINPUT98), .A4(new_n556), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT98), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n557), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n664), .A2(new_n665), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n524), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n525), .A2(new_n557), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  INV_X1    g0472(.A(new_n625), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT97), .B1(new_n588), .B2(new_n589), .ZN(new_n674));
  INV_X1    g0474(.A(new_n589), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT97), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n587), .A4(new_n585), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n673), .B1(new_n674), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n557), .A2(new_n561), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n664), .A2(new_n679), .A3(new_n631), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n669), .B(new_n672), .C1(new_n678), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n487), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n661), .A2(new_n682), .ZN(G369));
  NAND2_X1  g0483(.A1(new_n280), .A2(new_n207), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT100), .Z(new_n686));
  INV_X1    g0486(.A(G213), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n684), .B2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n625), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n633), .A2(new_n638), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n614), .A2(new_n691), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n576), .A2(new_n691), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n674), .A2(new_n677), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n594), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n696), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n625), .A2(new_n691), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n692), .B1(new_n588), .B2(new_n589), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n704), .B1(new_n694), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n703), .A2(new_n707), .ZN(G399));
  NOR2_X1   g0508(.A1(new_n211), .A2(G41), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G1), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n217), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT29), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n681), .A2(new_n715), .A3(new_n692), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT96), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n525), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n518), .A2(new_n524), .A3(KEYINPUT96), .ZN(new_n719));
  AND4_X1   g0519(.A1(new_n679), .A2(new_n631), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n636), .A2(new_n590), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n670), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n671), .A2(new_n665), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n718), .A2(new_n668), .A3(new_n666), .A4(new_n719), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n665), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n691), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n716), .B1(new_n726), .B2(new_n715), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n639), .A2(new_n567), .A3(new_n569), .A4(new_n692), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n618), .A2(new_n619), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n503), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(new_n553), .A3(new_n586), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n731), .A2(KEYINPUT30), .A3(new_n553), .A4(new_n586), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n621), .A2(new_n323), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n555), .A2(new_n591), .A3(new_n503), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n738), .B2(new_n691), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n728), .B1(new_n729), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n727), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n714), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(new_n701), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n700), .A2(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n279), .A2(G20), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n206), .B1(new_n748), .B2(G45), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n709), .A2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n746), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT101), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n371), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n207), .ZN(new_n755));
  INV_X1    g0555(.A(G294), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n207), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(new_n371), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n755), .A2(new_n756), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(G20), .A2(G179), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n761), .A2(new_n371), .A3(new_n363), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(G326), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n761), .A2(new_n371), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G322), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n763), .A2(new_n764), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G190), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n768), .B1(G329), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n761), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n769), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n761), .A2(new_n363), .A3(G190), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n775), .A2(G311), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n772), .A2(new_n383), .A3(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n760), .B(new_n779), .C1(G303), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n783), .A2(KEYINPUT103), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(KEYINPUT103), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n383), .B1(G87), .B2(new_n781), .ZN(new_n786));
  INV_X1    g0586(.A(G159), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n770), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT32), .ZN(new_n789));
  INV_X1    g0589(.A(new_n776), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n258), .A2(new_n766), .B1(new_n790), .B2(new_n271), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n763), .A2(new_n223), .B1(new_n774), .B2(new_n296), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n755), .A2(new_n528), .ZN(new_n794));
  INV_X1    g0594(.A(new_n758), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n794), .B1(G107), .B2(new_n795), .ZN(new_n796));
  AND4_X1   g0596(.A1(new_n786), .A2(new_n789), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n784), .A2(new_n785), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n215), .B1(G20), .B2(new_n519), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n751), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G13), .A2(G33), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n700), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n210), .A2(G116), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n211), .A2(new_n423), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n808), .B1(G45), .B2(new_n217), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n249), .B2(G45), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n211), .A2(new_n383), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n807), .B(new_n810), .C1(G355), .C2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT102), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n804), .B(new_n799), .C1(new_n812), .C2(KEYINPUT102), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n801), .B(new_n806), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n753), .A2(new_n815), .ZN(G396));
  INV_X1    g0616(.A(new_n751), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G137), .A2(new_n762), .B1(new_n765), .B2(G143), .ZN(new_n818));
  INV_X1    g0618(.A(G150), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n818), .B1(new_n819), .B2(new_n790), .C1(new_n787), .C2(new_n774), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT34), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(G132), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n423), .B1(new_n770), .B2(new_n823), .C1(new_n271), .C2(new_n758), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n755), .A2(new_n258), .B1(new_n780), .B2(new_n223), .ZN(new_n825));
  NOR3_X1   g0625(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n820), .A2(new_n821), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n758), .A2(new_n595), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n829), .B(new_n794), .C1(G107), .C2(new_n781), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n790), .A2(new_n759), .B1(new_n770), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(G303), .B2(new_n762), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n775), .A2(G116), .B1(G294), .B2(new_n765), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n830), .A2(new_n383), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n800), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n799), .A2(new_n802), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n817), .B(new_n836), .C1(new_n296), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n345), .A2(new_n691), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n353), .A2(new_n354), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n365), .B(new_n839), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n361), .B2(new_n839), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n838), .B1(new_n843), .B2(new_n803), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n681), .A2(new_n692), .ZN(new_n845));
  INV_X1    g0645(.A(new_n843), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT104), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n681), .A2(new_n692), .A3(new_n843), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(KEYINPUT104), .A3(new_n846), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n743), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n817), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n844), .B1(new_n855), .B2(new_n856), .ZN(G384));
  OR2_X1    g0657(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n533), .A2(KEYINPUT35), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(G116), .A3(new_n216), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  OAI211_X1 g0661(.A(new_n218), .B(G77), .C1(new_n258), .C2(new_n271), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n223), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n206), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT109), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n649), .A2(new_n692), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT106), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n257), .B1(new_n446), .B2(KEYINPUT16), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(KEYINPUT16), .B2(new_n446), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n435), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n689), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n641), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n870), .B1(new_n480), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n469), .A2(new_n689), .ZN(new_n877));
  AOI211_X1 g0677(.A(new_n434), .B(new_n478), .C1(new_n468), .C2(new_n452), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(KEYINPUT105), .B(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n431), .B2(new_n462), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n876), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n873), .A2(new_n874), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n869), .B(new_n883), .C1(new_n486), .C2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n886), .A2(KEYINPUT39), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n482), .A2(new_n643), .A3(new_n645), .A4(new_n483), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n877), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n879), .A2(new_n882), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n462), .A2(new_n641), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n462), .A2(new_n874), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(new_n892), .A3(new_n480), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n881), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n889), .A2(KEYINPUT107), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(new_n896), .A3(new_n877), .ZN(new_n897));
  AOI211_X1 g0697(.A(KEYINPUT108), .B(KEYINPUT38), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT108), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(KEYINPUT107), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n894), .A2(new_n890), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n900), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n899), .B1(new_n902), .B2(new_n869), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n887), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n884), .B1(new_n655), .B2(new_n473), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n869), .B1(new_n905), .B2(new_n883), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n486), .A2(new_n885), .ZN(new_n907));
  INV_X1    g0707(.A(new_n883), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n868), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n407), .A2(new_n691), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n413), .A2(new_n419), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n913), .B1(new_n413), .B2(new_n419), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n361), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n692), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n849), .B2(new_n918), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n910), .A2(new_n919), .B1(new_n646), .B2(new_n689), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n866), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n906), .B2(new_n909), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n888), .A2(new_n896), .A3(new_n877), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n896), .B1(new_n888), .B2(new_n877), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n881), .A2(new_n893), .B1(new_n879), .B2(new_n882), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT108), .B1(new_n928), .B2(KEYINPUT38), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n902), .A2(new_n899), .A3(new_n869), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n924), .B1(new_n931), .B2(new_n887), .ZN(new_n932));
  OAI211_X1 g0732(.A(KEYINPUT109), .B(new_n920), .C1(new_n932), .C2(new_n868), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n922), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n487), .A2(new_n727), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n661), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  OAI21_X1  g0737(.A(new_n909), .B1(new_n898), .B2(new_n903), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n843), .B1(new_n914), .B2(new_n915), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT110), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n739), .B1(new_n741), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n738), .A2(KEYINPUT110), .A3(KEYINPUT31), .A4(new_n691), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n939), .B1(new_n729), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT40), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n907), .B2(new_n908), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n944), .B1(new_n948), .B2(new_n886), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n729), .A2(new_n943), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n487), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n954), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(G330), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n937), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n206), .B2(new_n748), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n937), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n865), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT111), .ZN(G367));
  OAI21_X1  g0762(.A(new_n561), .B1(new_n634), .B2(new_n635), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n691), .B1(new_n963), .B2(new_n557), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT42), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n637), .B1(new_n636), .B2(new_n631), .ZN(new_n966));
  AND4_X1   g0766(.A1(new_n637), .A2(new_n627), .A3(new_n628), .A4(new_n631), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n706), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n557), .A2(new_n692), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n537), .A2(new_n691), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n969), .B1(new_n679), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n965), .B1(new_n968), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n705), .B1(new_n633), .B2(new_n638), .ZN(new_n973));
  INV_X1    g0773(.A(new_n971), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n973), .A2(KEYINPUT42), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n964), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n692), .A2(new_n517), .ZN(new_n977));
  MUX2_X1   g0777(.A(new_n664), .B(new_n670), .S(new_n977), .Z(new_n978));
  NOR2_X1   g0778(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n979));
  AND2_X1   g0779(.A1(new_n978), .A2(KEYINPUT43), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n976), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT112), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n976), .A2(new_n982), .A3(new_n979), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(new_n976), .B2(new_n979), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n702), .A2(new_n974), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n986), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n981), .B(new_n988), .C1(new_n983), .C2(new_n984), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n709), .B(KEYINPUT41), .Z(new_n990));
  INV_X1    g0790(.A(new_n704), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n968), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(KEYINPUT44), .B1(new_n992), .B2(new_n971), .ZN(new_n993));
  OAI211_X1 g0793(.A(KEYINPUT44), .B(new_n971), .C1(new_n973), .C2(new_n704), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT45), .B1(new_n707), .B2(new_n974), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n973), .A2(new_n997), .A3(new_n704), .A4(new_n971), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n993), .A2(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n702), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n968), .A2(KEYINPUT113), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT113), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n973), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n693), .B(new_n706), .C1(new_n694), .C2(new_n695), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n746), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n696), .A2(new_n705), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1007), .A2(new_n1001), .A3(new_n701), .A4(new_n1003), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n997), .B1(new_n992), .B2(new_n971), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n974), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n707), .B2(new_n974), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n994), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1015), .A3(new_n703), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1000), .A2(new_n744), .A3(new_n1009), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n990), .B1(new_n1017), .B2(new_n744), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n987), .B(new_n989), .C1(new_n1018), .C2(new_n750), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n804), .A2(new_n799), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n808), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1020), .B1(new_n210), .B2(new_n336), .C1(new_n1021), .C2(new_n243), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1022), .A2(new_n751), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n758), .A2(new_n296), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n755), .A2(new_n271), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G58), .C2(new_n781), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n766), .A2(new_n819), .B1(new_n774), .B2(new_n223), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G143), .B2(new_n762), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(KEYINPUT116), .B(G137), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n771), .A2(new_n1030), .B1(G159), .B2(new_n776), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1026), .A2(new_n293), .A3(new_n1028), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n755), .A2(new_n349), .B1(new_n774), .B2(new_n759), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT114), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n758), .A2(new_n528), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n443), .B1(new_n763), .B2(new_n831), .ZN(new_n1037));
  INV_X1    g0837(.A(G303), .ZN(new_n1038));
  INV_X1    g0838(.A(G317), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n766), .A2(new_n1038), .B1(new_n770), .B2(new_n1039), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT115), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n781), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT46), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n780), .B2(new_n496), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(new_n756), .C2(new_n790), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1041), .B1(new_n1034), .B2(new_n1033), .C1(new_n1042), .C2(new_n1046), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n1046), .A2(new_n1042), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1032), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT47), .Z(new_n1050));
  OAI221_X1 g0850(.A(new_n1023), .B1(new_n800), .B2(new_n1050), .C1(new_n978), .C2(new_n805), .ZN(new_n1051));
  AND3_X1   g0851(.A1(new_n1019), .A2(KEYINPUT117), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT117), .B1(new_n1019), .B2(new_n1051), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1052), .A2(new_n1053), .ZN(G387));
  NAND2_X1  g0854(.A1(new_n1009), .A2(new_n750), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n696), .A2(new_n804), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n443), .B1(new_n770), .B2(new_n764), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n755), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1058), .A2(G283), .B1(new_n781), .B2(G294), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n766), .A2(new_n1039), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n790), .A2(new_n831), .B1(new_n774), .B2(new_n1038), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1060), .B(new_n1061), .C1(G322), .C2(new_n762), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1059), .B1(new_n1062), .B2(KEYINPUT48), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(KEYINPUT48), .B2(new_n1062), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT49), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n1057), .B(new_n1065), .C1(G116), .C2(new_n795), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n443), .B(new_n1036), .C1(G150), .C2(new_n771), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n766), .A2(new_n223), .B1(new_n774), .B2(new_n271), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G159), .B2(new_n762), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n755), .A2(new_n336), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G77), .B2(new_n781), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n266), .B2(new_n776), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n799), .B1(new_n1066), .B2(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n240), .A2(new_n305), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n711), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1075), .A2(new_n808), .B1(new_n1076), .B2(new_n811), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT50), .B1(new_n330), .B2(G50), .ZN(new_n1078));
  AOI21_X1  g0878(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n711), .A3(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n330), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1077), .A2(new_n1082), .B1(G107), .B2(new_n210), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n817), .B1(new_n1083), .B2(new_n1020), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1056), .A2(new_n1074), .A3(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n744), .A2(new_n1009), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n709), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n744), .A2(new_n1009), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1055), .B(new_n1085), .C1(new_n1087), .C2(new_n1088), .ZN(G393));
  AND3_X1   g0889(.A1(new_n1012), .A2(new_n1015), .A3(new_n703), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n703), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1086), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n709), .A3(new_n1017), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n971), .A2(new_n804), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n780), .A2(new_n759), .B1(new_n770), .B2(new_n767), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT119), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n383), .B1(new_n349), .B2(new_n758), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n1097), .B2(new_n1096), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT120), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G317), .A2(new_n762), .B1(new_n765), .B2(G311), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT52), .Z(new_n1102));
  OAI22_X1  g0902(.A1(new_n790), .A2(new_n1038), .B1(new_n774), .B2(new_n756), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G116), .B2(new_n1058), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(G150), .A2(new_n762), .B1(new_n765), .B2(G159), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT51), .Z(new_n1107));
  OAI22_X1  g0907(.A1(new_n790), .A2(new_n223), .B1(new_n774), .B2(new_n330), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT118), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n443), .B(new_n829), .C1(G143), .C2(new_n771), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n755), .A2(new_n296), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G68), .B2(new_n781), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n800), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1020), .B1(new_n528), .B2(new_n210), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n808), .B2(new_n252), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(new_n817), .A3(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1094), .A2(new_n750), .B1(new_n1095), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1093), .A2(new_n1118), .ZN(G390));
  NAND2_X1  g0919(.A1(new_n953), .A2(G330), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1120), .A2(new_n939), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n849), .A2(new_n918), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n916), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n868), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n904), .A2(new_n1126), .A3(new_n911), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n868), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n721), .A2(new_n679), .A3(new_n631), .A4(new_n664), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n725), .A2(new_n1129), .A3(new_n524), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n692), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n918), .B1(new_n1131), .B2(new_n846), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1128), .B1(new_n1132), .B2(new_n1124), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n938), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1122), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT121), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n904), .A2(new_n911), .A3(new_n1126), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n743), .A2(new_n843), .A3(new_n1124), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n886), .B1(new_n929), .B2(new_n930), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n726), .A2(new_n843), .B1(new_n917), .B2(new_n692), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n868), .B1(new_n1140), .B2(new_n916), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1138), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1136), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n743), .A2(new_n843), .A3(new_n1124), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n938), .B2(new_n1133), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(KEYINPUT121), .A3(new_n1127), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1135), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n750), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n932), .A2(new_n802), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n817), .B1(new_n432), .B2(new_n837), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n383), .B1(new_n528), .B2(new_n774), .C1(new_n756), .C2(new_n770), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G283), .A2(new_n762), .B1(new_n765), .B2(G116), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1152), .B1(new_n349), .B2(new_n790), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n271), .A2(new_n758), .B1(new_n780), .B2(new_n595), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1111), .A4(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n771), .A2(G125), .B1(G128), .B2(new_n762), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n823), .B2(new_n766), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n293), .B1(new_n223), .B2(new_n758), .C1(new_n787), .C2(new_n755), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT122), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n790), .A2(new_n1029), .B1(new_n1160), .B2(new_n774), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1157), .B(new_n1158), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  OR3_X1    g0962(.A1(new_n780), .A2(KEYINPUT53), .A3(new_n819), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT53), .B1(new_n780), .B2(new_n819), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n1161), .C2(new_n1159), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1155), .B1(new_n1162), .B2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1149), .B(new_n1150), .C1(new_n800), .C2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n487), .A2(G330), .A3(new_n953), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1169), .A2(new_n935), .A3(new_n660), .A4(new_n329), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1124), .B1(new_n743), .B2(new_n843), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1123), .B1(new_n1121), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n916), .B1(new_n1120), .B2(new_n846), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n1140), .A3(new_n1138), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1170), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n709), .B1(new_n1147), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1121), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1145), .A2(KEYINPUT121), .A3(new_n1127), .ZN(new_n1179));
  AOI21_X1  g0979(.A(KEYINPUT121), .B1(new_n1145), .B2(new_n1127), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1178), .B(new_n1175), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1148), .B(new_n1168), .C1(new_n1176), .C2(new_n1182), .ZN(G378));
  OAI211_X1 g0983(.A(new_n951), .B(G330), .C1(new_n1139), .C2(new_n945), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n285), .A2(new_n689), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n659), .A2(new_n325), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1186), .B1(new_n659), .B2(new_n325), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n1190), .B(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1184), .A2(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n947), .A2(new_n1192), .A3(G330), .A4(new_n951), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n934), .A2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n922), .A2(new_n1194), .A3(new_n933), .A4(new_n1195), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n750), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n817), .B1(new_n223), .B2(new_n837), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n443), .A2(new_n304), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(G97), .B2(new_n776), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n349), .B2(new_n766), .C1(new_n496), .C2(new_n763), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n774), .A2(new_n336), .B1(new_n770), .B2(new_n759), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n258), .A2(new_n758), .B1(new_n780), .B2(new_n296), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1203), .A2(new_n1025), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT58), .Z(new_n1207));
  AOI22_X1  g1007(.A1(new_n775), .A2(G137), .B1(G128), .B2(new_n765), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(G125), .A2(new_n762), .B1(new_n776), .B2(G132), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n755), .A2(new_n819), .B1(new_n780), .B2(new_n1160), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n795), .A2(G159), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n771), .C2(G124), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1201), .B(new_n223), .C1(G33), .C2(G41), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1207), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1221), .A2(KEYINPUT123), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n799), .B1(new_n1221), .B2(KEYINPUT123), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1200), .B1(new_n1222), .B2(new_n1223), .C1(new_n1192), .C2(new_n803), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1199), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1174), .A2(new_n1172), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1170), .B1(new_n1147), .B2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1197), .A2(KEYINPUT57), .A3(new_n1198), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n709), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AND4_X1   g1030(.A1(new_n922), .A2(new_n1194), .A3(new_n933), .A4(new_n1195), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n922), .A2(new_n933), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1170), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1181), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT57), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1226), .B1(new_n1230), .B2(new_n1236), .ZN(G375));
  NOR2_X1   g1037(.A1(new_n1227), .A2(new_n1234), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(new_n990), .A3(new_n1175), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1227), .A2(new_n750), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n817), .B1(new_n271), .B2(new_n837), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n766), .A2(new_n1029), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n763), .A2(new_n823), .B1(new_n790), .B2(new_n1160), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G128), .C2(new_n771), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n423), .B1(new_n774), .B2(new_n819), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n755), .A2(new_n223), .B1(new_n780), .B2(new_n787), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(G58), .C2(new_n795), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(G294), .A2(new_n762), .B1(new_n776), .B2(G116), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(new_n349), .B2(new_n774), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n766), .A2(new_n759), .B1(new_n770), .B2(new_n1038), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1249), .A2(new_n293), .A3(new_n1250), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1024), .B(new_n1070), .C1(G97), .C2(new_n781), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1244), .A2(new_n1247), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1241), .B1(new_n800), .B2(new_n1253), .C1(new_n1124), .C2(new_n803), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1240), .A2(new_n1254), .ZN(new_n1255));
  OR2_X1    g1055(.A1(new_n1239), .A2(new_n1255), .ZN(G381));
  OR2_X1    g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  OR4_X1    g1057(.A1(G384), .A2(G381), .A3(new_n1257), .A4(G390), .ZN(new_n1258));
  OR4_X1    g1058(.A1(G387), .A2(new_n1258), .A3(G378), .A4(G375), .ZN(G407));
  OAI21_X1  g1059(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1168), .B1(new_n1260), .B2(new_n749), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1175), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n710), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1181), .B2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n687), .A2(G343), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(G407), .B(G213), .C1(G375), .C2(new_n1266), .ZN(G409));
  INV_X1    g1067(.A(KEYINPUT124), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G384), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1227), .A2(new_n1234), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(new_n710), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1175), .A2(new_n1270), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1272), .B1(new_n1273), .B2(new_n1238), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(G384), .A2(new_n1268), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1275), .A2(new_n1255), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1269), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1276), .A3(new_n1269), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1278), .A2(G2897), .A3(new_n1265), .A4(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1265), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1279), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1281), .B1(new_n1282), .B2(new_n1277), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(G378), .B(new_n1226), .C1(new_n1230), .C2(new_n1236), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1228), .A2(new_n1287), .A3(new_n990), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1264), .B1(new_n1288), .B2(new_n1225), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1286), .A2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1265), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  AOI211_X1 g1093(.A(new_n1293), .B(new_n1265), .C1(new_n1286), .C2(new_n1289), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1285), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1265), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G393), .A2(G396), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1017), .A2(new_n744), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n990), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n750), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n987), .A2(new_n989), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G390), .B(new_n1051), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  AOI21_X1  g1105(.A(G390), .B1(new_n1019), .B2(new_n1051), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1257), .B(new_n1299), .C1(new_n1305), .C2(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1052), .A2(new_n1053), .A3(G390), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(KEYINPUT126), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1257), .A2(new_n1299), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT126), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1019), .A2(new_n1311), .A3(new_n1051), .A4(G390), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1309), .A2(new_n1310), .A3(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1307), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1290), .A2(new_n1297), .A3(new_n1291), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1316), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1295), .A2(new_n1298), .A3(new_n1319), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1317), .A2(KEYINPUT62), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1315), .B1(new_n1296), .B2(new_n1284), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1323), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1321), .A2(new_n1322), .A3(new_n1324), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1320), .B1(new_n1325), .B2(new_n1314), .ZN(G405));
  NAND2_X1  g1126(.A1(G375), .A2(new_n1264), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1314), .A2(new_n1286), .A3(KEYINPUT127), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1314), .B1(KEYINPUT127), .B2(new_n1286), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1297), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1286), .A2(KEYINPUT127), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1314), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1314), .A2(new_n1286), .A3(KEYINPUT127), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(new_n1327), .A3(new_n1336), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1331), .A2(new_n1332), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1332), .B1(new_n1331), .B2(new_n1337), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(G402));
endmodule


