

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n680, n681, n682, n683, n684, n685, n688, n689, n690, n691,
         n692, n694, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781;

  XNOR2_X1 U370 ( .A(n349), .B(n348), .ZN(G51) );
  XNOR2_X1 U371 ( .A(n351), .B(n350), .ZN(G60) );
  AND2_X1 U372 ( .A1(n353), .A2(n352), .ZN(n681) );
  INV_X1 U373 ( .A(n694), .ZN(n348) );
  INV_X1 U374 ( .A(KEYINPUT60), .ZN(n350) );
  INV_X1 U375 ( .A(n710), .ZN(n352) );
  INV_X1 U376 ( .A(n710), .ZN(n355) );
  INV_X1 U377 ( .A(n710), .ZN(n358) );
  AND2_X1 U378 ( .A1(n565), .A2(n507), .ZN(n652) );
  XNOR2_X1 U379 ( .A(n595), .B(n594), .ZN(n608) );
  NOR2_X1 U380 ( .A1(n607), .A2(n725), .ZN(n595) );
  XNOR2_X1 U381 ( .A(n490), .B(KEYINPUT113), .ZN(n565) );
  OR2_X1 U382 ( .A1(n561), .A2(n556), .ZN(n633) );
  AND2_X1 U383 ( .A1(n593), .A2(n592), .ZN(n545) );
  XNOR2_X1 U384 ( .A(n505), .B(KEYINPUT94), .ZN(n735) );
  XNOR2_X1 U385 ( .A(n492), .B(n491), .ZN(n362) );
  XNOR2_X1 U386 ( .A(n516), .B(KEYINPUT16), .ZN(n361) );
  XNOR2_X1 U387 ( .A(KEYINPUT71), .B(n383), .ZN(n517) );
  INV_X2 U388 ( .A(G902), .ZN(n535) );
  NAND2_X1 U389 ( .A1(n551), .A2(n552), .ZN(n553) );
  NAND2_X1 U390 ( .A1(n356), .A2(n355), .ZN(n349) );
  NAND2_X1 U391 ( .A1(n359), .A2(n358), .ZN(n351) );
  XNOR2_X2 U392 ( .A(n603), .B(KEYINPUT109), .ZN(n552) );
  NAND2_X1 U393 ( .A1(n545), .A2(n412), .ZN(n603) );
  XNOR2_X2 U394 ( .A(n487), .B(n375), .ZN(n673) );
  XNOR2_X1 U395 ( .A(n677), .B(n354), .ZN(n353) );
  INV_X1 U396 ( .A(n676), .ZN(n354) );
  XNOR2_X1 U397 ( .A(n692), .B(n357), .ZN(n356) );
  INV_X1 U398 ( .A(n691), .ZN(n357) );
  XNOR2_X1 U399 ( .A(n685), .B(n360), .ZN(n359) );
  INV_X1 U400 ( .A(n684), .ZN(n360) );
  XNOR2_X1 U401 ( .A(n362), .B(n361), .ZN(n371) );
  XNOR2_X2 U402 ( .A(n432), .B(n387), .ZN(n749) );
  NOR2_X2 U403 ( .A1(n650), .A2(n649), .ZN(n651) );
  OR2_X2 U404 ( .A1(n707), .A2(G902), .ZN(n488) );
  XNOR2_X2 U405 ( .A(n653), .B(KEYINPUT47), .ZN(n427) );
  XNOR2_X1 U406 ( .A(n667), .B(KEYINPUT72), .ZN(n365) );
  XNOR2_X1 U407 ( .A(n662), .B(n388), .ZN(n372) );
  AND2_X1 U408 ( .A1(n369), .A2(n437), .ZN(n368) );
  INV_X2 U409 ( .A(G953), .ZN(n773) );
  INV_X1 U410 ( .A(KEYINPUT35), .ZN(n431) );
  NOR2_X1 U411 ( .A1(n712), .A2(n501), .ZN(n363) );
  NAND2_X1 U412 ( .A1(n372), .A2(n434), .ZN(n666) );
  AND2_X1 U413 ( .A1(n400), .A2(n384), .ZN(n615) );
  XNOR2_X1 U414 ( .A(n409), .B(n431), .ZN(n611) );
  NAND2_X1 U415 ( .A1(n403), .A2(n404), .ZN(n409) );
  AND2_X1 U416 ( .A1(n608), .A2(n419), .ZN(n415) );
  NOR2_X1 U417 ( .A1(n640), .A2(n639), .ZN(n642) );
  INV_X1 U418 ( .A(n604), .ZN(n722) );
  NAND2_X1 U419 ( .A1(n367), .A2(n436), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n389), .B(n390), .ZN(n542) );
  XOR2_X1 U421 ( .A(KEYINPUT59), .B(n683), .Z(n684) );
  AND2_X1 U422 ( .A1(n735), .A2(n438), .ZN(n436) );
  INV_X1 U423 ( .A(KEYINPUT31), .ZN(n594) );
  XOR2_X1 U424 ( .A(KEYINPUT112), .B(KEYINPUT28), .Z(n479) );
  XNOR2_X1 U425 ( .A(G110), .B(G119), .ZN(n461) );
  XOR2_X1 U426 ( .A(KEYINPUT110), .B(KEYINPUT30), .Z(n547) );
  NAND2_X1 U427 ( .A1(n364), .A2(n363), .ZN(n672) );
  INV_X1 U428 ( .A(n713), .ZN(n364) );
  NAND2_X1 U429 ( .A1(n365), .A2(n669), .ZN(n380) );
  AND2_X1 U430 ( .A1(n365), .A2(KEYINPUT2), .ZN(n754) );
  NAND2_X2 U431 ( .A1(n368), .A2(n366), .ZN(n636) );
  INV_X1 U432 ( .A(n542), .ZN(n367) );
  NAND2_X1 U433 ( .A1(n542), .A2(KEYINPUT87), .ZN(n369) );
  INV_X1 U434 ( .A(n370), .ZN(n631) );
  OR2_X1 U435 ( .A1(n371), .A2(n630), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n500), .B(n371), .ZN(n688) );
  AND2_X1 U437 ( .A1(n372), .A2(n423), .ZN(n772) );
  NAND2_X1 U438 ( .A1(n373), .A2(n670), .ZN(n667) );
  XNOR2_X1 U439 ( .A(n373), .B(KEYINPUT72), .ZN(n713) );
  XNOR2_X2 U440 ( .A(n666), .B(KEYINPUT81), .ZN(n373) );
  XNOR2_X1 U441 ( .A(n587), .B(G110), .ZN(G12) );
  XNOR2_X2 U442 ( .A(n374), .B(G472), .ZN(n546) );
  OR2_X2 U443 ( .A1(n673), .A2(G902), .ZN(n374) );
  INV_X1 U444 ( .A(n446), .ZN(n375) );
  XNOR2_X2 U445 ( .A(n771), .B(G146), .ZN(n487) );
  XNOR2_X2 U446 ( .A(n377), .B(n376), .ZN(n492) );
  XNOR2_X2 U447 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n376) );
  XNOR2_X2 U448 ( .A(G119), .B(G116), .ZN(n377) );
  XNOR2_X2 U449 ( .A(n378), .B(G107), .ZN(n491) );
  XNOR2_X2 U450 ( .A(G101), .B(G110), .ZN(n378) );
  XNOR2_X2 U451 ( .A(n379), .B(G104), .ZN(n516) );
  XNOR2_X2 U452 ( .A(G113), .B(G122), .ZN(n379) );
  NAND2_X1 U453 ( .A1(n380), .A2(n672), .ZN(n381) );
  NAND2_X1 U454 ( .A1(n380), .A2(n672), .ZN(n696) );
  XNOR2_X2 U455 ( .A(n575), .B(n426), .ZN(n425) );
  BUF_X1 U456 ( .A(n532), .Z(n382) );
  AND2_X1 U457 ( .A1(n736), .A2(n421), .ZN(n419) );
  INV_X1 U458 ( .A(KEYINPUT104), .ZN(n421) );
  NAND2_X1 U459 ( .A1(n418), .A2(n417), .ZN(n416) );
  OR2_X1 U460 ( .A1(n736), .A2(n421), .ZN(n417) );
  XNOR2_X1 U461 ( .A(G143), .B(G140), .ZN(n511) );
  INV_X1 U462 ( .A(KEYINPUT66), .ZN(n401) );
  NOR2_X1 U463 ( .A1(n396), .A2(n405), .ZN(n403) );
  NOR2_X1 U464 ( .A1(n749), .A2(n407), .ZN(n396) );
  INV_X1 U465 ( .A(KEYINPUT22), .ZN(n426) );
  INV_X1 U466 ( .A(KEYINPUT1), .ZN(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT91), .B(KEYINPUT15), .ZN(n447) );
  NAND2_X1 U468 ( .A1(n422), .A2(n420), .ZN(n413) );
  INV_X1 U469 ( .A(KEYINPUT87), .ZN(n438) );
  OR2_X1 U470 ( .A1(n735), .A2(n438), .ZN(n437) );
  INV_X1 U471 ( .A(G237), .ZN(n502) );
  XNOR2_X1 U472 ( .A(G101), .B(G113), .ZN(n442) );
  XNOR2_X1 U473 ( .A(n511), .B(n510), .ZN(n512) );
  INV_X1 U474 ( .A(KEYINPUT12), .ZN(n510) );
  NAND2_X1 U475 ( .A1(G234), .A2(G237), .ZN(n453) );
  INV_X1 U476 ( .A(n665), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n428), .B(n462), .ZN(n465) );
  XNOR2_X1 U478 ( .A(n463), .B(n461), .ZN(n428) );
  XNOR2_X1 U479 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n460) );
  XNOR2_X1 U480 ( .A(G137), .B(G140), .ZN(n483) );
  INV_X1 U481 ( .A(KEYINPUT2), .ZN(n435) );
  INV_X1 U482 ( .A(KEYINPUT39), .ZN(n582) );
  NOR2_X1 U483 ( .A1(n433), .A2(n715), .ZN(n432) );
  NAND2_X1 U484 ( .A1(n599), .A2(n545), .ZN(n433) );
  NAND2_X1 U485 ( .A1(n385), .A2(n643), .ZN(n725) );
  XNOR2_X1 U486 ( .A(n675), .B(n674), .ZN(n676) );
  BUF_X1 U487 ( .A(n696), .Z(n705) );
  XNOR2_X1 U488 ( .A(n689), .B(n690), .ZN(n691) );
  XNOR2_X1 U489 ( .A(n678), .B(KEYINPUT90), .ZN(n710) );
  XOR2_X1 U490 ( .A(KEYINPUT42), .B(n566), .Z(n649) );
  XNOR2_X1 U491 ( .A(n646), .B(n645), .ZN(n656) );
  XNOR2_X1 U492 ( .A(n397), .B(KEYINPUT32), .ZN(n424) );
  OR2_X1 U493 ( .A1(n557), .A2(n560), .ZN(n763) );
  OR2_X1 U494 ( .A1(G953), .A2(G237), .ZN(n383) );
  INV_X1 U495 ( .A(n715), .ZN(n643) );
  AND2_X1 U496 ( .A1(n610), .A2(n609), .ZN(n384) );
  NOR2_X1 U497 ( .A1(n395), .A2(n714), .ZN(n385) );
  AND2_X1 U498 ( .A1(n590), .A2(n589), .ZN(n386) );
  INV_X1 U499 ( .A(KEYINPUT34), .ZN(n410) );
  XNOR2_X1 U500 ( .A(KEYINPUT106), .B(KEYINPUT33), .ZN(n387) );
  XOR2_X1 U501 ( .A(n661), .B(KEYINPUT67), .Z(n388) );
  NOR2_X1 U502 ( .A1(n688), .A2(n671), .ZN(n389) );
  XOR2_X1 U503 ( .A(n503), .B(KEYINPUT78), .Z(n390) );
  XOR2_X1 U504 ( .A(G107), .B(G122), .Z(n525) );
  XNOR2_X1 U505 ( .A(n625), .B(n624), .ZN(n391) );
  XNOR2_X1 U506 ( .A(n625), .B(n624), .ZN(n670) );
  NAND2_X1 U507 ( .A1(n551), .A2(n552), .ZN(n392) );
  XNOR2_X1 U508 ( .A(n392), .B(KEYINPUT73), .ZN(n393) );
  XNOR2_X1 U509 ( .A(n553), .B(KEYINPUT73), .ZN(n581) );
  AND2_X1 U510 ( .A1(n565), .A2(n507), .ZN(n394) );
  BUF_X1 U511 ( .A(n604), .Z(n395) );
  NAND2_X1 U512 ( .A1(n406), .A2(n601), .ZN(n405) );
  NAND2_X1 U513 ( .A1(n425), .A2(n386), .ZN(n397) );
  INV_X1 U514 ( .A(n591), .ZN(n607) );
  BUF_X1 U515 ( .A(n634), .Z(n398) );
  BUF_X1 U516 ( .A(n650), .Z(n399) );
  NAND2_X1 U517 ( .A1(n602), .A2(n424), .ZN(n617) );
  NAND2_X1 U518 ( .A1(n414), .A2(n413), .ZN(n610) );
  NAND2_X1 U519 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U520 ( .A1(n425), .A2(n715), .ZN(n585) );
  NAND2_X1 U521 ( .A1(n660), .A2(n659), .ZN(n662) );
  NAND2_X1 U522 ( .A1(n617), .A2(KEYINPUT44), .ZN(n402) );
  NAND2_X1 U523 ( .A1(n617), .A2(KEYINPUT66), .ZN(n612) );
  NAND2_X1 U524 ( .A1(n607), .A2(KEYINPUT34), .ZN(n406) );
  XNOR2_X1 U525 ( .A(n585), .B(KEYINPUT105), .ZN(n430) );
  NOR2_X2 U526 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U527 ( .A1(n749), .A2(KEYINPUT34), .ZN(n404) );
  NAND2_X1 U528 ( .A1(n408), .A2(n410), .ZN(n407) );
  INV_X1 U529 ( .A(n607), .ZN(n408) );
  XNOR2_X2 U530 ( .A(n412), .B(n411), .ZN(n715) );
  XNOR2_X2 U531 ( .A(n488), .B(G469), .ZN(n412) );
  NAND2_X1 U532 ( .A1(n489), .A2(n412), .ZN(n490) );
  NOR2_X1 U533 ( .A1(n415), .A2(n416), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n757), .A2(n419), .ZN(n418) );
  NOR2_X1 U535 ( .A1(n757), .A2(n421), .ZN(n420) );
  INV_X1 U536 ( .A(n608), .ZN(n422) );
  XNOR2_X1 U537 ( .A(n424), .B(G119), .ZN(G21) );
  XNOR2_X1 U538 ( .A(n487), .B(n486), .ZN(n707) );
  NOR2_X1 U539 ( .A1(n665), .A2(n435), .ZN(n434) );
  NAND2_X1 U540 ( .A1(n581), .A2(n580), .ZN(n583) );
  NOR2_X2 U541 ( .A1(n427), .A2(n654), .ZN(n655) );
  AND2_X2 U542 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X2 U543 ( .A1(n572), .A2(n571), .ZN(n429) );
  XNOR2_X2 U544 ( .A(n429), .B(KEYINPUT0), .ZN(n591) );
  NAND2_X1 U545 ( .A1(n430), .A2(n586), .ZN(n602) );
  XNOR2_X2 U546 ( .A(n498), .B(n440), .ZN(n771) );
  XNOR2_X2 U547 ( .A(n532), .B(KEYINPUT4), .ZN(n498) );
  INV_X1 U548 ( .A(n611), .ZN(n619) );
  NAND2_X1 U549 ( .A1(n546), .A2(n735), .ZN(n548) );
  XNOR2_X2 U550 ( .A(n636), .B(KEYINPUT19), .ZN(n572) );
  XNOR2_X1 U551 ( .A(n513), .B(n512), .ZN(n515) );
  INV_X1 U552 ( .A(KEYINPUT114), .ZN(n645) );
  BUF_X1 U553 ( .A(n602), .Z(n587) );
  XNOR2_X2 U554 ( .A(G143), .B(KEYINPUT65), .ZN(n439) );
  XNOR2_X2 U555 ( .A(n439), .B(G128), .ZN(n532) );
  XNOR2_X1 U556 ( .A(G134), .B(G131), .ZN(n440) );
  XNOR2_X1 U557 ( .A(G137), .B(KEYINPUT5), .ZN(n441) );
  XNOR2_X1 U558 ( .A(n442), .B(n441), .ZN(n444) );
  NAND2_X1 U559 ( .A1(n517), .A2(G210), .ZN(n443) );
  XNOR2_X1 U560 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U561 ( .A(n492), .B(n445), .ZN(n446) );
  INV_X1 U562 ( .A(n546), .ZN(n604) );
  XNOR2_X1 U563 ( .A(n447), .B(n535), .ZN(n501) );
  NAND2_X1 U564 ( .A1(n501), .A2(G234), .ZN(n448) );
  XNOR2_X1 U565 ( .A(n448), .B(KEYINPUT20), .ZN(n471) );
  INV_X1 U566 ( .A(n471), .ZN(n450) );
  INV_X1 U567 ( .A(G221), .ZN(n449) );
  OR2_X1 U568 ( .A1(n450), .A2(n449), .ZN(n452) );
  INV_X1 U569 ( .A(KEYINPUT21), .ZN(n451) );
  XNOR2_X1 U570 ( .A(n452), .B(n451), .ZN(n592) );
  XNOR2_X1 U571 ( .A(n453), .B(KEYINPUT14), .ZN(n457) );
  AND2_X1 U572 ( .A1(G953), .A2(n457), .ZN(n454) );
  NAND2_X1 U573 ( .A1(G902), .A2(n454), .ZN(n567) );
  XOR2_X1 U574 ( .A(n567), .B(KEYINPUT108), .Z(n456) );
  INV_X1 U575 ( .A(G900), .ZN(n455) );
  NAND2_X1 U576 ( .A1(n456), .A2(n455), .ZN(n458) );
  NAND2_X1 U577 ( .A1(G952), .A2(n457), .ZN(n746) );
  OR2_X1 U578 ( .A1(n746), .A2(G953), .ZN(n569) );
  NAND2_X1 U579 ( .A1(n458), .A2(n569), .ZN(n549) );
  NAND2_X1 U580 ( .A1(n592), .A2(n549), .ZN(n459) );
  XNOR2_X1 U581 ( .A(n459), .B(KEYINPUT68), .ZN(n637) );
  XOR2_X1 U582 ( .A(KEYINPUT23), .B(KEYINPUT75), .Z(n463) );
  XNOR2_X1 U583 ( .A(n460), .B(G128), .ZN(n462) );
  XNOR2_X2 U584 ( .A(G146), .B(G125), .ZN(n494) );
  XNOR2_X1 U585 ( .A(n494), .B(KEYINPUT10), .ZN(n514) );
  INV_X1 U586 ( .A(n483), .ZN(n464) );
  XNOR2_X1 U587 ( .A(n514), .B(n464), .ZN(n770) );
  XNOR2_X1 U588 ( .A(n465), .B(n770), .ZN(n470) );
  AND2_X1 U589 ( .A1(G234), .A2(n773), .ZN(n466) );
  XNOR2_X1 U590 ( .A(KEYINPUT8), .B(n466), .ZN(n530) );
  NAND2_X1 U591 ( .A1(n530), .A2(G221), .ZN(n468) );
  XNOR2_X1 U592 ( .A(KEYINPUT97), .B(KEYINPUT79), .ZN(n467) );
  XNOR2_X1 U593 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U594 ( .A(n470), .B(n469), .ZN(n697) );
  NAND2_X1 U595 ( .A1(n697), .A2(n535), .ZN(n477) );
  NAND2_X1 U596 ( .A1(n471), .A2(G217), .ZN(n475) );
  XNOR2_X1 U597 ( .A(KEYINPUT98), .B(KEYINPUT99), .ZN(n473) );
  XNOR2_X1 U598 ( .A(KEYINPUT25), .B(KEYINPUT74), .ZN(n472) );
  XNOR2_X1 U599 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U600 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X2 U601 ( .A(n477), .B(n476), .ZN(n593) );
  NOR2_X1 U602 ( .A1(n637), .A2(n593), .ZN(n478) );
  NAND2_X1 U603 ( .A1(n722), .A2(n478), .ZN(n480) );
  XNOR2_X1 U604 ( .A(n480), .B(n479), .ZN(n489) );
  XNOR2_X1 U605 ( .A(G104), .B(KEYINPUT76), .ZN(n481) );
  XNOR2_X1 U606 ( .A(n491), .B(n481), .ZN(n485) );
  NAND2_X1 U607 ( .A1(G227), .A2(n773), .ZN(n482) );
  XNOR2_X1 U608 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U609 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U610 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n493) );
  XNOR2_X1 U611 ( .A(n494), .B(n493), .ZN(n497) );
  NAND2_X1 U612 ( .A1(n773), .A2(G224), .ZN(n495) );
  XNOR2_X1 U613 ( .A(n495), .B(KEYINPUT93), .ZN(n496) );
  XNOR2_X1 U614 ( .A(n497), .B(n496), .ZN(n499) );
  XNOR2_X1 U615 ( .A(n498), .B(n499), .ZN(n500) );
  INV_X1 U616 ( .A(n501), .ZN(n671) );
  NAND2_X1 U617 ( .A1(n535), .A2(n502), .ZN(n504) );
  NAND2_X1 U618 ( .A1(n504), .A2(G210), .ZN(n503) );
  NAND2_X1 U619 ( .A1(n504), .A2(G214), .ZN(n505) );
  INV_X1 U620 ( .A(n735), .ZN(n731) );
  BUF_X1 U621 ( .A(n572), .Z(n506) );
  INV_X1 U622 ( .A(n506), .ZN(n507) );
  XOR2_X1 U623 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n509) );
  XNOR2_X1 U624 ( .A(G131), .B(KEYINPUT100), .ZN(n508) );
  XNOR2_X1 U625 ( .A(n509), .B(n508), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n515), .B(n514), .ZN(n521) );
  INV_X1 U627 ( .A(n516), .ZN(n519) );
  NAND2_X1 U628 ( .A1(n517), .A2(G214), .ZN(n518) );
  XNOR2_X1 U629 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U630 ( .A(n521), .B(n520), .ZN(n682) );
  NAND2_X1 U631 ( .A1(n682), .A2(n535), .ZN(n523) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(G475), .ZN(n522) );
  XNOR2_X1 U633 ( .A(n523), .B(n522), .ZN(n561) );
  XNOR2_X1 U634 ( .A(G116), .B(G134), .ZN(n524) );
  XNOR2_X1 U635 ( .A(n525), .B(n524), .ZN(n529) );
  XOR2_X1 U636 ( .A(KEYINPUT102), .B(KEYINPUT7), .Z(n527) );
  XNOR2_X1 U637 ( .A(KEYINPUT9), .B(KEYINPUT103), .ZN(n526) );
  XNOR2_X1 U638 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U639 ( .A(n529), .B(n528), .Z(n534) );
  NAND2_X1 U640 ( .A1(n530), .A2(G217), .ZN(n531) );
  XNOR2_X1 U641 ( .A(n382), .B(n531), .ZN(n533) );
  XNOR2_X1 U642 ( .A(n534), .B(n533), .ZN(n701) );
  NAND2_X1 U643 ( .A1(n701), .A2(n535), .ZN(n536) );
  XNOR2_X1 U644 ( .A(n536), .B(G478), .ZN(n556) );
  XNOR2_X2 U645 ( .A(n633), .B(KEYINPUT107), .ZN(n758) );
  NAND2_X1 U646 ( .A1(n394), .A2(n758), .ZN(n537) );
  XNOR2_X1 U647 ( .A(n537), .B(G146), .ZN(G48) );
  INV_X1 U648 ( .A(n593), .ZN(n718) );
  NAND2_X1 U649 ( .A1(n758), .A2(n718), .ZN(n538) );
  XNOR2_X1 U650 ( .A(n546), .B(KEYINPUT6), .ZN(n588) );
  OR2_X1 U651 ( .A1(n538), .A2(n588), .ZN(n640) );
  NOR2_X1 U652 ( .A1(n637), .A2(n731), .ZN(n539) );
  NAND2_X1 U653 ( .A1(n715), .A2(n539), .ZN(n540) );
  NOR2_X1 U654 ( .A1(n640), .A2(n540), .ZN(n541) );
  XOR2_X1 U655 ( .A(KEYINPUT43), .B(n541), .Z(n544) );
  BUF_X1 U656 ( .A(n542), .Z(n543) );
  NAND2_X1 U657 ( .A1(n544), .A2(n543), .ZN(n663) );
  XNOR2_X1 U658 ( .A(n663), .B(G140), .ZN(G42) );
  XNOR2_X1 U659 ( .A(n548), .B(n547), .ZN(n550) );
  INV_X1 U660 ( .A(n561), .ZN(n557) );
  NAND2_X1 U661 ( .A1(n557), .A2(n556), .ZN(n600) );
  NOR2_X1 U662 ( .A1(n600), .A2(n543), .ZN(n554) );
  NAND2_X1 U663 ( .A1(n393), .A2(n554), .ZN(n555) );
  XNOR2_X1 U664 ( .A(n555), .B(KEYINPUT111), .ZN(n654) );
  XOR2_X1 U665 ( .A(G143), .B(n654), .Z(G45) );
  XNOR2_X1 U666 ( .A(G128), .B(KEYINPUT29), .ZN(n559) );
  INV_X1 U667 ( .A(n556), .ZN(n560) );
  INV_X1 U668 ( .A(n763), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n394), .A2(n597), .ZN(n558) );
  XOR2_X1 U670 ( .A(n559), .B(n558), .Z(G30) );
  AND2_X1 U671 ( .A1(n561), .A2(n560), .ZN(n732) );
  NAND2_X1 U672 ( .A1(n732), .A2(n735), .ZN(n563) );
  XNOR2_X1 U673 ( .A(KEYINPUT70), .B(KEYINPUT38), .ZN(n562) );
  XNOR2_X1 U674 ( .A(n543), .B(n562), .ZN(n580) );
  INV_X1 U675 ( .A(n580), .ZN(n737) );
  OR2_X1 U676 ( .A1(n737), .A2(n563), .ZN(n564) );
  XNOR2_X1 U677 ( .A(n564), .B(KEYINPUT41), .ZN(n729) );
  NAND2_X1 U678 ( .A1(n565), .A2(n729), .ZN(n566) );
  XOR2_X1 U679 ( .A(G137), .B(n649), .Z(G39) );
  NOR2_X1 U680 ( .A1(G898), .A2(n567), .ZN(n568) );
  XNOR2_X1 U681 ( .A(n568), .B(KEYINPUT95), .ZN(n570) );
  AND2_X1 U682 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U683 ( .A(n732), .ZN(n573) );
  INV_X1 U684 ( .A(n592), .ZN(n717) );
  NOR2_X1 U685 ( .A1(n573), .A2(n717), .ZN(n574) );
  NAND2_X1 U686 ( .A1(n591), .A2(n574), .ZN(n575) );
  BUF_X1 U687 ( .A(n585), .Z(n576) );
  INV_X1 U688 ( .A(n576), .ZN(n578) );
  INV_X1 U689 ( .A(n588), .ZN(n599) );
  NOR2_X1 U690 ( .A1(n599), .A2(n718), .ZN(n577) );
  NAND2_X1 U691 ( .A1(n578), .A2(n577), .ZN(n609) );
  XOR2_X1 U692 ( .A(G101), .B(KEYINPUT115), .Z(n579) );
  XNOR2_X1 U693 ( .A(n609), .B(n579), .ZN(G3) );
  XNOR2_X2 U694 ( .A(n583), .B(n582), .ZN(n634) );
  INV_X1 U695 ( .A(n398), .ZN(n584) );
  NAND2_X1 U696 ( .A1(n584), .A2(n597), .ZN(n664) );
  XNOR2_X1 U697 ( .A(n664), .B(G134), .ZN(G36) );
  NOR2_X1 U698 ( .A1(n722), .A2(n593), .ZN(n586) );
  XOR2_X1 U699 ( .A(KEYINPUT77), .B(n588), .Z(n590) );
  NOR2_X1 U700 ( .A1(n715), .A2(n593), .ZN(n589) );
  NAND2_X1 U701 ( .A1(n593), .A2(n592), .ZN(n714) );
  NAND2_X1 U702 ( .A1(n608), .A2(n758), .ZN(n596) );
  XNOR2_X1 U703 ( .A(n596), .B(G113), .ZN(G15) );
  NAND2_X1 U704 ( .A1(n608), .A2(n597), .ZN(n598) );
  XNOR2_X1 U705 ( .A(n598), .B(G116), .ZN(G18) );
  INV_X1 U706 ( .A(n600), .ZN(n601) );
  XNOR2_X1 U707 ( .A(n611), .B(G122), .ZN(G24) );
  INV_X1 U708 ( .A(n603), .ZN(n605) );
  NAND2_X1 U709 ( .A1(n605), .A2(n395), .ZN(n606) );
  NOR2_X1 U710 ( .A1(n607), .A2(n606), .ZN(n757) );
  NAND2_X1 U711 ( .A1(n763), .A2(n633), .ZN(n736) );
  NAND2_X1 U712 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U713 ( .A1(n613), .A2(KEYINPUT44), .ZN(n614) );
  NAND2_X1 U714 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U715 ( .A(n616), .B(KEYINPUT85), .ZN(n623) );
  BUF_X1 U716 ( .A(n617), .Z(n618) );
  INV_X1 U717 ( .A(n618), .ZN(n621) );
  NOR2_X1 U718 ( .A1(n619), .A2(KEYINPUT44), .ZN(n620) );
  NAND2_X1 U719 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U720 ( .A1(n623), .A2(n622), .ZN(n625) );
  XNOR2_X1 U721 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n624) );
  NAND2_X1 U722 ( .A1(n391), .A2(n773), .ZN(n629) );
  NAND2_X1 U723 ( .A1(G953), .A2(G224), .ZN(n626) );
  XNOR2_X1 U724 ( .A(KEYINPUT61), .B(n626), .ZN(n627) );
  NAND2_X1 U725 ( .A1(n627), .A2(G898), .ZN(n628) );
  NAND2_X1 U726 ( .A1(n629), .A2(n628), .ZN(n632) );
  NOR2_X1 U727 ( .A1(G898), .A2(n773), .ZN(n630) );
  XNOR2_X1 U728 ( .A(n632), .B(n631), .ZN(G69) );
  XNOR2_X1 U729 ( .A(n635), .B(KEYINPUT40), .ZN(n650) );
  XOR2_X1 U730 ( .A(n399), .B(G131), .Z(G33) );
  INV_X1 U731 ( .A(n637), .ZN(n638) );
  NAND2_X1 U732 ( .A1(n636), .A2(n638), .ZN(n639) );
  XNOR2_X1 U733 ( .A(KEYINPUT86), .B(KEYINPUT36), .ZN(n641) );
  XNOR2_X1 U734 ( .A(n642), .B(n641), .ZN(n644) );
  NAND2_X1 U735 ( .A1(n644), .A2(n643), .ZN(n646) );
  XOR2_X1 U736 ( .A(KEYINPUT120), .B(KEYINPUT37), .Z(n647) );
  XOR2_X1 U737 ( .A(n647), .B(G125), .Z(n648) );
  XNOR2_X1 U738 ( .A(n656), .B(n648), .ZN(G27) );
  XNOR2_X1 U739 ( .A(n651), .B(KEYINPUT46), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n652), .A2(n736), .ZN(n653) );
  XNOR2_X1 U741 ( .A(n655), .B(KEYINPUT69), .ZN(n658) );
  XNOR2_X1 U742 ( .A(n656), .B(KEYINPUT84), .ZN(n657) );
  NOR2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U744 ( .A(KEYINPUT83), .B(KEYINPUT48), .ZN(n661) );
  NAND2_X1 U745 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U746 ( .A(n671), .B(KEYINPUT80), .ZN(n668) );
  AND2_X1 U747 ( .A1(KEYINPUT2), .A2(n668), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n391), .A2(n772), .ZN(n712) );
  NAND2_X1 U749 ( .A1(n696), .A2(G472), .ZN(n677) );
  BUF_X1 U750 ( .A(n673), .Z(n675) );
  XOR2_X1 U751 ( .A(KEYINPUT89), .B(KEYINPUT62), .Z(n674) );
  NOR2_X1 U752 ( .A1(n773), .A2(G952), .ZN(n678) );
  XOR2_X1 U753 ( .A(KEYINPUT88), .B(KEYINPUT63), .Z(n680) );
  XNOR2_X1 U754 ( .A(n681), .B(n680), .ZN(G57) );
  NAND2_X1 U755 ( .A1(n381), .A2(G475), .ZN(n685) );
  INV_X1 U756 ( .A(n682), .ZN(n683) );
  NAND2_X1 U757 ( .A1(n381), .A2(G210), .ZN(n692) );
  BUF_X1 U758 ( .A(n688), .Z(n689) );
  XOR2_X1 U759 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n690) );
  XNOR2_X1 U760 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n705), .A2(G217), .ZN(n699) );
  XNOR2_X1 U762 ( .A(n697), .B(KEYINPUT125), .ZN(n698) );
  XNOR2_X1 U763 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U764 ( .A1(n700), .A2(n710), .ZN(G66) );
  NAND2_X1 U765 ( .A1(n705), .A2(G478), .ZN(n703) );
  XOR2_X1 U766 ( .A(n701), .B(KEYINPUT124), .Z(n702) );
  XNOR2_X1 U767 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U768 ( .A1(n704), .A2(n710), .ZN(G63) );
  NAND2_X1 U769 ( .A1(n705), .A2(G469), .ZN(n709) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  XNOR2_X1 U771 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U772 ( .A(n709), .B(n708), .ZN(n711) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(G54) );
  OR2_X1 U774 ( .A1(n713), .A2(n712), .ZN(n753) );
  NAND2_X1 U775 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U776 ( .A(n716), .B(KEYINPUT50), .ZN(n724) );
  NAND2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n720) );
  XOR2_X1 U778 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n719) );
  XNOR2_X1 U779 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U780 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U781 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U783 ( .A(KEYINPUT51), .B(KEYINPUT122), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n728), .B(n727), .ZN(n730) );
  INV_X1 U785 ( .A(n729), .ZN(n748) );
  NOR2_X1 U786 ( .A1(n730), .A2(n748), .ZN(n743) );
  NAND2_X1 U787 ( .A1(n737), .A2(n731), .ZN(n733) );
  NAND2_X1 U788 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n734), .B(KEYINPUT123), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n736), .A2(n735), .ZN(n738) );
  NOR2_X1 U791 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U792 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n749), .A2(n741), .ZN(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U795 ( .A(n744), .B(KEYINPUT52), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n747) );
  OR2_X1 U797 ( .A1(n747), .A2(G953), .ZN(n751) );
  NOR2_X1 U798 ( .A1(n749), .A2(n748), .ZN(n750) );
  NOR2_X1 U799 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n753), .A2(n752), .ZN(n755) );
  NOR2_X1 U801 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U802 ( .A(n756), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U803 ( .A(n757), .ZN(n764) );
  INV_X1 U804 ( .A(n758), .ZN(n759) );
  NOR2_X1 U805 ( .A1(n764), .A2(n759), .ZN(n761) );
  XNOR2_X1 U806 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n760) );
  XNOR2_X1 U807 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U808 ( .A(G104), .B(n762), .ZN(G6) );
  NOR2_X1 U809 ( .A1(n764), .A2(n763), .ZN(n769) );
  XOR2_X1 U810 ( .A(KEYINPUT27), .B(KEYINPUT119), .Z(n766) );
  XNOR2_X1 U811 ( .A(G107), .B(KEYINPUT26), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n766), .B(n765), .ZN(n767) );
  XNOR2_X1 U813 ( .A(KEYINPUT118), .B(n767), .ZN(n768) );
  XNOR2_X1 U814 ( .A(n769), .B(n768), .ZN(G9) );
  XNOR2_X1 U815 ( .A(n771), .B(n770), .ZN(n775) );
  XNOR2_X1 U816 ( .A(n772), .B(n775), .ZN(n774) );
  NAND2_X1 U817 ( .A1(n774), .A2(n773), .ZN(n781) );
  XOR2_X1 U818 ( .A(G227), .B(n775), .Z(n776) );
  XNOR2_X1 U819 ( .A(n776), .B(KEYINPUT126), .ZN(n777) );
  NAND2_X1 U820 ( .A1(n777), .A2(G900), .ZN(n778) );
  XOR2_X1 U821 ( .A(KEYINPUT127), .B(n778), .Z(n779) );
  NAND2_X1 U822 ( .A1(G953), .A2(n779), .ZN(n780) );
  NAND2_X1 U823 ( .A1(n781), .A2(n780), .ZN(G72) );
endmodule

