//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  XNOR2_X1  g000(.A(KEYINPUT75), .B(G125), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT16), .A2(G140), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G125), .A2(G140), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n187), .B2(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(KEYINPUT16), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  AOI211_X1 g010(.A(new_n196), .B(new_n189), .C1(KEYINPUT16), .C2(new_n193), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G214), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n199), .A2(G237), .A3(G953), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n201), .B1(new_n206), .B2(new_n200), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT17), .A3(G131), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n207), .B(G131), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n198), .B(new_n208), .C1(KEYINPUT17), .C2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G113), .B(G122), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n211), .B(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT18), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  OAI221_X1 g029(.A(new_n201), .B1(new_n214), .B2(new_n215), .C1(new_n206), .C2(new_n200), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G125), .B(G140), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n196), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n220), .B(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n196), .B2(new_n193), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n207), .A2(KEYINPUT18), .A3(G131), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n218), .B(new_n223), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n210), .A2(new_n213), .A3(new_n227), .ZN(new_n228));
  OAI211_X1 g042(.A(KEYINPUT19), .B(new_n191), .C1(new_n187), .C2(new_n192), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT19), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT84), .B1(new_n219), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT84), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(new_n229), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(new_n196), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n194), .A2(G146), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n209), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n213), .B1(new_n227), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n228), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(G475), .A2(G902), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT85), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT20), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n238), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n210), .A2(new_n227), .A3(new_n213), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT20), .ZN(new_n246));
  INV_X1    g060(.A(new_n241), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G902), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n213), .B1(new_n210), .B2(new_n227), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n249), .B1(new_n228), .B2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n242), .A2(new_n248), .B1(G475), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G952), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(G234), .B2(G237), .ZN(new_n255));
  AOI211_X1 g069(.A(new_n249), .B(new_n253), .C1(G234), .C2(G237), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT21), .B(G898), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G122), .ZN(new_n263));
  INV_X1    g077(.A(G122), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G116), .ZN(new_n265));
  NOR3_X1   g079(.A1(new_n263), .A2(new_n265), .A3(G107), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n262), .A2(G122), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT14), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT91), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n268), .A2(new_n269), .A3(new_n263), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT14), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n270), .B1(new_n271), .B2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(G107), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n268), .B2(new_n269), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT87), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n202), .B2(G128), .ZN(new_n277));
  INV_X1    g091(.A(G128), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(KEYINPUT87), .A3(G143), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n203), .A2(new_n205), .A3(G128), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G134), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n281), .A3(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n283), .A2(KEYINPUT90), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT90), .B1(new_n283), .B2(new_n285), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n275), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(KEYINPUT9), .B(G234), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(G217), .A3(new_n253), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n285), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT88), .A4(new_n284), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT86), .A2(KEYINPUT13), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT86), .A2(KEYINPUT13), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n281), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n280), .B1(new_n281), .B2(new_n299), .ZN(new_n301));
  OAI21_X1  g115(.A(G134), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n264), .A2(G116), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n273), .B1(new_n303), .B2(new_n267), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n266), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AND4_X1   g120(.A1(KEYINPUT89), .A2(new_n296), .A3(new_n302), .A4(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n294), .B2(new_n295), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT89), .B1(new_n308), .B2(new_n302), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n288), .B(new_n292), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n288), .B1(new_n307), .B2(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n291), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n296), .A2(new_n302), .A3(new_n306), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n308), .A2(KEYINPUT89), .A3(new_n302), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n319), .A2(KEYINPUT92), .A3(new_n288), .A4(new_n292), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n312), .A2(new_n314), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n249), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT93), .ZN(new_n323));
  INV_X1    g137(.A(G478), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n324), .A2(KEYINPUT15), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT93), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n326), .A3(new_n249), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n322), .A2(new_n325), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n328), .A2(KEYINPUT94), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT94), .B1(new_n328), .B2(new_n330), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n261), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G221), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n290), .B2(new_n249), .ZN(new_n335));
  XNOR2_X1  g149(.A(G110), .B(G140), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n253), .A2(G227), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n284), .B2(G137), .ZN(new_n340));
  INV_X1    g154(.A(G137), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT11), .A3(G134), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n284), .A2(G137), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n340), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(G131), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n348), .A2(new_n273), .A3(G104), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n212), .A2(G107), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(KEYINPUT78), .B(G101), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n273), .A2(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n350), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n351), .A2(new_n352), .B1(G101), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT64), .B(G143), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT1), .B1(new_n356), .B2(G146), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT66), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n202), .B2(G146), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n196), .A2(KEYINPUT66), .A3(G143), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n203), .A2(new_n205), .A3(G146), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n357), .A2(G128), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n278), .A2(KEYINPUT1), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n355), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AND2_X1   g182(.A1(KEYINPUT0), .A2(G128), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n362), .A2(new_n359), .A3(new_n360), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n361), .A2(new_n372), .A3(new_n362), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n375), .B1(new_n202), .B2(G146), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n376), .B1(new_n356), .B2(G146), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n206), .A2(new_n375), .A3(new_n196), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT0), .A2(G128), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n369), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g195(.A1(new_n352), .A2(new_n347), .A3(new_n349), .A4(new_n350), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n383));
  AOI22_X1  g197(.A1(new_n382), .A2(KEYINPUT4), .B1(G101), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n383), .A2(KEYINPUT4), .A3(G101), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n374), .B(new_n381), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n212), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n273), .A2(G104), .ZN(new_n388));
  OAI21_X1  g202(.A(G101), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT78), .B(G101), .Z(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(KEYINPUT10), .C1(new_n383), .C2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G128), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n377), .A2(new_n378), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n361), .A2(new_n362), .A3(new_n364), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n346), .A2(new_n368), .A3(new_n386), .A4(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n396), .B1(new_n366), .B2(new_n367), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n346), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n338), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n346), .A3(new_n386), .ZN(new_n402));
  INV_X1    g216(.A(new_n338), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n382), .A2(new_n389), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n394), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n366), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT12), .B1(new_n406), .B2(new_n345), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT12), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n346), .C1(new_n366), .C2(new_n405), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n402), .B(new_n403), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n401), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n249), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT79), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(G902), .B1(new_n401), .B2(new_n410), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT79), .A3(new_n412), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n398), .A2(new_n338), .ZN(new_n419));
  INV_X1    g233(.A(new_n400), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n402), .B1(new_n407), .B2(new_n409), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n419), .A2(new_n420), .B1(new_n421), .B2(new_n338), .ZN(new_n422));
  OAI21_X1  g236(.A(G469), .B1(new_n422), .B2(G902), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n335), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT75), .B(G125), .Z(new_n427));
  NAND3_X1  g241(.A1(new_n374), .A2(new_n381), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n394), .A2(new_n395), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n187), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n253), .A2(G224), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n428), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n428), .B2(new_n430), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n262), .A2(G119), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT69), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT69), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n437), .A3(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(KEYINPUT2), .B(G113), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n438), .A2(new_n442), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n384), .B2(new_n385), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT5), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n439), .B2(new_n441), .ZN(new_n448));
  OAI21_X1  g262(.A(G113), .B1(new_n436), .B2(KEYINPUT5), .ZN(new_n449));
  OAI211_X1 g263(.A(new_n355), .B(new_n444), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n446), .A2(new_n450), .A3(new_n452), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n452), .B1(new_n446), .B2(new_n450), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT80), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n458), .B1(new_n457), .B2(new_n459), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n434), .B(new_n456), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n428), .A2(new_n430), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n431), .A2(KEYINPUT7), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n428), .A2(KEYINPUT7), .A3(new_n430), .A4(new_n431), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n452), .B(KEYINPUT8), .Z(new_n468));
  NOR2_X1   g282(.A1(new_n438), .A2(new_n447), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n444), .B1(new_n469), .B2(new_n449), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n468), .B1(new_n470), .B2(new_n355), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n444), .B1(new_n448), .B2(new_n449), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n471), .B1(new_n472), .B2(new_n355), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n473), .A2(new_n455), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n462), .A2(new_n477), .A3(new_n475), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n426), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n424), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n333), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n374), .A2(new_n345), .A3(new_n381), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n344), .A2(G131), .ZN(new_n485));
  INV_X1    g299(.A(new_n343), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n284), .A2(G137), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n429), .A2(new_n485), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(new_n489), .A3(KEYINPUT30), .ZN(new_n490));
  INV_X1    g304(.A(new_n489), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT68), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n484), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n374), .A2(KEYINPUT68), .A3(new_n345), .A4(new_n381), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n445), .B(new_n490), .C1(new_n495), .C2(KEYINPUT30), .ZN(new_n496));
  XOR2_X1   g310(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n497));
  INV_X1    g311(.A(G237), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n253), .A3(G210), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n497), .B(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n445), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n484), .A2(new_n489), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n496), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT31), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n496), .A2(KEYINPUT31), .A3(new_n503), .A4(new_n505), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n505), .B(new_n511), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n495), .A2(new_n504), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT32), .ZN(new_n516));
  NOR2_X1   g330(.A1(G472), .A2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n514), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n508), .B2(new_n509), .ZN(new_n520));
  INV_X1    g334(.A(new_n517), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT32), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n496), .A2(new_n505), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n502), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n512), .A2(new_n513), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n503), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n484), .A2(new_n489), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n445), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(KEYINPUT71), .A3(new_n505), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT71), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n532), .A3(new_n445), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n531), .A2(KEYINPUT28), .A3(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT72), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n505), .B2(new_n511), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n531), .A2(new_n535), .A3(KEYINPUT28), .A4(new_n533), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n502), .A2(new_n527), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n528), .A2(new_n541), .A3(new_n249), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n518), .A2(new_n522), .B1(G472), .B2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  INV_X1    g358(.A(G234), .ZN(new_n545));
  NOR3_X1   g359(.A1(new_n334), .A2(new_n545), .A3(G953), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n544), .B(new_n546), .Z(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  XOR2_X1   g362(.A(KEYINPUT24), .B(G110), .Z(new_n549));
  XNOR2_X1  g363(.A(G119), .B(G128), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT23), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n435), .B2(G128), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n278), .A2(KEYINPUT23), .A3(G119), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n554), .B(new_n555), .C1(G119), .C2(new_n278), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G110), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT74), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n559), .A3(G110), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n552), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n195), .B2(new_n197), .ZN(new_n562));
  OAI22_X1  g376(.A1(new_n556), .A2(G110), .B1(new_n550), .B2(new_n549), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n236), .A2(new_n222), .A3(new_n563), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n562), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT77), .B1(new_n562), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n548), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n548), .B1(new_n562), .B2(new_n564), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(G217), .B1(new_n545), .B2(G902), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT73), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(G902), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n249), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT25), .ZN(new_n577));
  AOI21_X1  g391(.A(G902), .B1(new_n567), .B2(new_n569), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n572), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n575), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n543), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n483), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(new_n390), .ZN(G3));
  NAND2_X1  g399(.A1(new_n515), .A2(new_n517), .ZN(new_n586));
  OAI21_X1  g400(.A(G472), .B1(new_n520), .B2(G902), .ZN(new_n587));
  AND2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND4_X1   g402(.A1(KEYINPUT79), .A2(new_n411), .A3(new_n412), .A4(new_n249), .ZN(new_n589));
  AOI21_X1  g403(.A(KEYINPUT79), .B1(new_n416), .B2(new_n412), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n423), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n335), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n581), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n462), .A2(new_n477), .A3(new_n475), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n477), .B1(new_n462), .B2(new_n475), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n425), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT95), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT95), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(new_n425), .C1(new_n596), .C2(new_n597), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n599), .A2(new_n259), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n251), .A2(G475), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n239), .A2(KEYINPUT20), .A3(new_n241), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n246), .B1(new_n245), .B2(new_n247), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT96), .B(KEYINPUT33), .Z(new_n608));
  NAND2_X1  g422(.A1(new_n321), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n314), .A2(KEYINPUT33), .A3(new_n310), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n324), .A2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT97), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n609), .A2(new_n616), .A3(new_n610), .A4(new_n612), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n602), .A2(new_n603), .A3(new_n607), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n607), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n599), .A2(new_n259), .A3(new_n601), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT98), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n595), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT34), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NOR2_X1   g439(.A1(new_n331), .A2(new_n332), .ZN(new_n626));
  INV_X1    g440(.A(new_n604), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n248), .B1(new_n606), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n605), .A2(new_n242), .A3(KEYINPUT99), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n626), .A2(new_n602), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n595), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  INV_X1    g449(.A(KEYINPUT94), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n321), .A2(new_n326), .A3(new_n249), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n326), .B1(new_n321), .B2(new_n249), .ZN(new_n638));
  INV_X1    g452(.A(new_n325), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n636), .B1(new_n640), .B2(new_n329), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n328), .A2(KEYINPUT94), .A3(new_n330), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n260), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n591), .A2(new_n592), .A3(new_n481), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT77), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n556), .A2(new_n559), .A3(G110), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n559), .B1(new_n556), .B2(G110), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n551), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n194), .A2(G146), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n236), .ZN(new_n650));
  INV_X1    g464(.A(new_n564), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n645), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n562), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n653));
  OAI211_X1 g467(.A(new_n652), .B(new_n653), .C1(KEYINPUT36), .C2(new_n548), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n548), .A2(KEYINPUT36), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n565), .B2(new_n566), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n574), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n547), .B1(new_n652), .B2(new_n653), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n579), .B(new_n249), .C1(new_n659), .C2(new_n568), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n573), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n579), .B1(new_n570), .B2(new_n249), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT100), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OAI211_X1 g479(.A(KEYINPUT100), .B(new_n658), .C1(new_n661), .C2(new_n662), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n643), .A2(new_n644), .A3(new_n588), .A4(new_n667), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  INV_X1    g484(.A(new_n255), .ZN(new_n671));
  INV_X1    g485(.A(new_n256), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n671), .B1(new_n672), .B2(G900), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n642), .A2(new_n641), .A3(new_n631), .A4(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n665), .A2(new_n592), .A3(new_n591), .A4(new_n666), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n599), .A2(new_n601), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n542), .A2(G472), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n520), .A2(KEYINPUT32), .A3(new_n521), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n674), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  INV_X1    g497(.A(new_n663), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n626), .A2(new_n607), .A3(new_n425), .A4(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n685), .A2(KEYINPUT102), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(KEYINPUT102), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n479), .A2(new_n480), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(KEYINPUT38), .Z(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n531), .A2(new_n533), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n502), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT101), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n694), .A3(new_n502), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n693), .A2(new_n506), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n696), .B2(G902), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n679), .B2(new_n680), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n690), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n686), .A2(new_n687), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n673), .B(KEYINPUT39), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n424), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(new_n703), .B(KEYINPUT40), .Z(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n700), .A2(KEYINPUT103), .ZN(new_n706));
  OR2_X1    g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n206), .ZN(G45));
  AND3_X1   g522(.A1(new_n618), .A2(new_n607), .A3(new_n673), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n677), .A2(new_n681), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  NAND2_X1  g525(.A1(new_n619), .A2(new_n622), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  OAI221_X1 g527(.A(new_n592), .B1(new_n412), .B2(new_n416), .C1(new_n589), .C2(new_n590), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n543), .A2(new_n582), .A3(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n713), .B1(new_n712), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  INV_X1    g534(.A(new_n632), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n715), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  INV_X1    g537(.A(new_n416), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n415), .A2(new_n417), .B1(G469), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n599), .A3(new_n592), .A4(new_n601), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n665), .A2(new_n666), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n543), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n643), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NOR2_X1   g544(.A1(new_n714), .A2(new_n258), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n510), .B1(new_n503), .B2(new_n539), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n517), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n731), .A2(new_n581), .A3(new_n587), .A4(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(new_n676), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n626), .A2(KEYINPUT105), .A3(new_n607), .A4(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n641), .A2(new_n642), .A3(new_n607), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n737), .B1(new_n738), .B2(new_n676), .ZN(new_n739));
  AOI211_X1 g553(.A(KEYINPUT106), .B(new_n734), .C1(new_n736), .C2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT106), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n739), .ZN(new_n742));
  INV_X1    g556(.A(new_n734), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n264), .ZN(G24));
  NAND2_X1  g560(.A1(new_n733), .A2(new_n587), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n747), .A2(new_n684), .ZN(new_n748));
  INV_X1    g562(.A(new_n726), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n709), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT107), .B(G125), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G27));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n592), .A2(new_n425), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n419), .A2(new_n420), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n421), .A2(new_n338), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n412), .B1(new_n757), .B2(new_n249), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n249), .A3(G469), .ZN(new_n760));
  OAI22_X1  g574(.A1(new_n758), .A2(new_n759), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n688), .B(new_n754), .C1(new_n761), .C2(new_n418), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n709), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n681), .A2(new_n581), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n753), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n583), .A2(KEYINPUT42), .A3(new_n709), .A4(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  AND2_X1   g582(.A1(new_n674), .A2(new_n762), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n583), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  NAND2_X1  g585(.A1(new_n618), .A2(new_n252), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT43), .B1(new_n252), .B2(KEYINPUT109), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n586), .A2(new_n587), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n663), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n422), .A2(KEYINPUT45), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n422), .A2(KEYINPUT45), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(G469), .A2(G902), .ZN(new_n783));
  AOI21_X1  g597(.A(KEYINPUT46), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n784), .B1(new_n415), .B2(new_n417), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n783), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n335), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n702), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n688), .A2(new_n426), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n778), .A2(new_n779), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  XNOR2_X1  g607(.A(new_n787), .B(KEYINPUT47), .ZN(new_n794));
  AND4_X1   g608(.A1(new_n543), .A2(new_n709), .A3(new_n582), .A4(new_n789), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  XOR2_X1   g613(.A(KEYINPUT111), .B(G140), .Z(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G42));
  AND2_X1   g615(.A1(new_n774), .A2(new_n255), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n714), .A2(new_n790), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n583), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT48), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n747), .A2(new_n582), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n749), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n254), .B(KEYINPUT119), .Z(new_n810));
  NAND3_X1  g624(.A1(new_n803), .A2(new_n581), .A3(new_n255), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n698), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n813));
  INV_X1    g627(.A(new_n620), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n805), .A2(new_n809), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT50), .ZN(new_n818));
  INV_X1    g632(.A(new_n714), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n689), .A2(new_n819), .A3(new_n426), .ZN(new_n820));
  OR3_X1    g634(.A1(new_n807), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n818), .B1(new_n807), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n618), .A2(new_n607), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n813), .A2(new_n815), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n802), .A2(new_n748), .A3(new_n803), .ZN(new_n826));
  INV_X1    g640(.A(new_n725), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n592), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n808), .B(new_n789), .C1(new_n794), .C2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n823), .A2(new_n825), .A3(new_n826), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n817), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n831), .B2(new_n830), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT120), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n721), .A2(new_n715), .B1(new_n728), .B2(new_n643), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n716), .B2(new_n717), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n745), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n586), .A2(new_n587), .A3(new_n665), .A4(new_n666), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n333), .A2(new_n839), .A3(new_n482), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n252), .B1(new_n640), .B2(new_n329), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n481), .A2(new_n259), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n775), .A2(new_n593), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n838), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n842), .ZN(new_n845));
  INV_X1    g659(.A(new_n841), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n588), .A2(new_n594), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n668), .A2(KEYINPUT113), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n775), .A2(new_n593), .A3(new_n842), .ZN(new_n849));
  AOI22_X1  g663(.A1(new_n483), .A2(new_n583), .B1(new_n849), .B2(new_n814), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT114), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n844), .A2(new_n850), .A3(KEYINPUT114), .A4(new_n848), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n673), .A2(new_n592), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n856), .B(new_n663), .C1(new_n761), .C2(new_n418), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n698), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n742), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n681), .B(new_n677), .C1(new_n674), .C2(new_n709), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n750), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n682), .A2(new_n710), .A3(new_n750), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n858), .B1(new_n736), .B2(new_n739), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT52), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n748), .A2(new_n709), .A3(new_n762), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n631), .A2(new_n673), .A3(new_n789), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n869), .A2(new_n675), .A3(new_n329), .A4(new_n640), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n681), .ZN(new_n871));
  AND4_X1   g685(.A1(new_n767), .A2(new_n770), .A3(new_n868), .A4(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n837), .A2(new_n855), .A3(new_n867), .A4(new_n872), .ZN(new_n873));
  XOR2_X1   g687(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n874));
  OR2_X1    g688(.A1(new_n740), .A2(new_n744), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n722), .A2(new_n729), .ZN(new_n876));
  INV_X1    g690(.A(new_n717), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT113), .B1(new_n668), .B2(new_n847), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n814), .A2(new_n588), .A3(new_n594), .A4(new_n845), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n643), .A2(new_n644), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n764), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT114), .B1(new_n884), .B2(new_n848), .ZN(new_n885));
  AND4_X1   g699(.A1(KEYINPUT114), .A2(new_n844), .A3(new_n848), .A4(new_n850), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n875), .B(new_n879), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n770), .A2(new_n868), .A3(new_n871), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n889), .B1(new_n765), .B2(new_n766), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n888), .A2(new_n863), .A3(new_n866), .A4(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT117), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n866), .A2(new_n888), .A3(new_n890), .A4(new_n863), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT117), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(new_n894), .A3(new_n855), .A4(new_n837), .ZN(new_n895));
  AOI221_X4 g709(.A(KEYINPUT54), .B1(new_n873), .B2(new_n874), .C1(new_n892), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n837), .A2(new_n855), .A3(new_n872), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT115), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n837), .A2(new_n855), .A3(new_n900), .A4(new_n872), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n867), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n889), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n873), .A2(new_n874), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n897), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI22_X1  g721(.A1(new_n834), .A2(new_n907), .B1(G952), .B2(G953), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n581), .A2(new_n592), .A3(new_n425), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n910), .A2(KEYINPUT112), .B1(KEYINPUT49), .B2(new_n827), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(KEYINPUT49), .B2(new_n827), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n689), .B1(new_n910), .B2(KEYINPUT112), .ZN(new_n913));
  OR4_X1    g727(.A1(new_n698), .A2(new_n912), .A3(new_n772), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n908), .A2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n253), .A2(G952), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT121), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n892), .A2(new_n895), .B1(new_n873), .B2(new_n874), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n249), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n919), .A2(new_n478), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n434), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT55), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n917), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n919), .A2(G210), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n923), .B1(new_n927), .B2(new_n924), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n926), .A2(new_n928), .ZN(G51));
  XOR2_X1   g743(.A(new_n783), .B(KEYINPUT57), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n892), .A2(new_n895), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n873), .A2(new_n874), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n906), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n896), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n411), .ZN(new_n935));
  OR3_X1    g749(.A1(new_n918), .A2(new_n249), .A3(new_n782), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n916), .B1(new_n935), .B2(new_n936), .ZN(G54));
  AND2_X1   g751(.A1(KEYINPUT58), .A2(G475), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n919), .A2(new_n245), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n245), .B1(new_n919), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n916), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT59), .Z(new_n943));
  NOR2_X1   g757(.A1(new_n611), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n896), .B2(new_n933), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT122), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT122), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n944), .C1(new_n896), .C2(new_n933), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n903), .A2(new_n904), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n896), .B1(new_n950), .B2(KEYINPUT54), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n611), .B1(new_n951), .B2(new_n943), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n949), .A2(new_n952), .A3(new_n917), .ZN(G63));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n955));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n918), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n955), .B1(new_n958), .B2(new_n657), .ZN(new_n959));
  INV_X1    g773(.A(new_n657), .ZN(new_n960));
  NOR4_X1   g774(.A1(new_n918), .A2(KEYINPUT123), .A3(new_n960), .A4(new_n957), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n917), .B1(new_n958), .B2(new_n570), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n954), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n963), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(KEYINPUT61), .C1(new_n959), .C2(new_n961), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(G66));
  INV_X1    g781(.A(G224), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n257), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n887), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(G953), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n921), .B1(G898), .B2(new_n253), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n971), .B(new_n973), .ZN(G69));
  OAI21_X1  g788(.A(new_n490), .B1(new_n495), .B2(KEYINPUT30), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(new_n234), .Z(new_n976));
  INV_X1    g790(.A(new_n707), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT62), .B1(new_n977), .B2(new_n864), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n707), .A2(new_n979), .A3(new_n750), .A4(new_n862), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n792), .A2(new_n799), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n703), .A2(new_n790), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n583), .B(new_n982), .C1(new_n814), .C2(new_n846), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT125), .Z(new_n984));
  NAND4_X1  g798(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n976), .B1(new_n985), .B2(new_n253), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n253), .B1(G227), .B2(G900), .ZN(new_n987));
  NAND2_X1  g801(.A1(G900), .A2(G953), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n976), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n788), .B1(new_n739), .B2(new_n736), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n583), .B1(new_n990), .B2(new_n769), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n864), .B1(new_n766), .B2(new_n765), .ZN(new_n992));
  AND4_X1   g806(.A1(new_n792), .A2(new_n991), .A3(new_n799), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n989), .B1(new_n993), .B2(new_n253), .ZN(new_n994));
  OR3_X1    g808(.A1(new_n986), .A2(new_n987), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n987), .B1(new_n986), .B2(new_n994), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G72));
  NAND2_X1  g811(.A1(G472), .A2(G902), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT63), .Z(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n985), .B2(new_n887), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n502), .B1(new_n496), .B2(new_n505), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n993), .A2(new_n970), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n503), .B(new_n523), .C1(new_n1003), .C2(new_n999), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1004), .A2(new_n916), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1005), .A2(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1007));
  NOR3_X1   g821(.A1(new_n1004), .A2(new_n1007), .A3(new_n916), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1002), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n524), .A2(new_n506), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n999), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT127), .Z(new_n1012));
  NOR2_X1   g826(.A1(new_n905), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1009), .A2(new_n1013), .ZN(G57));
endmodule


