//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1248,
    new_n1249, new_n1251, new_n1252, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT0), .ZN(new_n206));
  OAI21_X1  g0006(.A(G50), .B1(G58), .B2(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n206), .B(new_n212), .C1(KEYINPUT1), .C2(new_n222), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n223), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XNOR2_X1  g0024(.A(G238), .B(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(KEYINPUT2), .B(G226), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(G169), .ZN(new_n241));
  NAND2_X1  g0041(.A1(G33), .A2(G41), .ZN(new_n242));
  NAND3_X1  g0042(.A1(new_n242), .A2(G1), .A3(G13), .ZN(new_n243));
  OR2_X1    g0043(.A1(KEYINPUT3), .A2(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(KEYINPUT3), .A2(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n246), .A2(G232), .A3(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT68), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g0050(.A1(new_n246), .A2(KEYINPUT68), .A3(G232), .A4(new_n247), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(new_n247), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n256), .A2(G238), .B1(G107), .B2(new_n255), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n243), .B1(new_n252), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n243), .A3(G274), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n243), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n263), .B1(G244), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n241), .B1(new_n258), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n271), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n272));
  AOI21_X1  g0072(.A(KEYINPUT65), .B1(new_n271), .B2(new_n209), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT15), .B(G87), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n210), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G77), .ZN(new_n277));
  OAI22_X1  g0077(.A1(new_n275), .A2(new_n276), .B1(new_n210), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n274), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n271), .A2(new_n209), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT65), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n271), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n277), .B1(new_n264), .B2(G20), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n277), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n283), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT69), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n283), .A2(new_n291), .A3(KEYINPUT69), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n246), .A2(G1698), .ZN(new_n300));
  INV_X1    g0100(.A(G107), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n300), .A2(new_n217), .B1(new_n301), .B2(new_n246), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n250), .B2(new_n251), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n299), .B(new_n268), .C1(new_n303), .C2(new_n243), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n270), .A2(new_n298), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n296), .A2(KEYINPUT70), .A3(new_n297), .ZN(new_n306));
  OAI211_X1 g0106(.A(G190), .B(new_n268), .C1(new_n303), .C2(new_n243), .ZN(new_n307));
  OAI21_X1  g0107(.A(G200), .B1(new_n258), .B2(new_n269), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT70), .B1(new_n296), .B2(new_n297), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n210), .A2(G33), .A3(G77), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n312), .B1(new_n210), .B2(G68), .C1(new_n281), .C2(new_n214), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n274), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT11), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n264), .A2(G20), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n288), .A2(G68), .A3(new_n289), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n292), .A2(new_n216), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT12), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n274), .A2(new_n313), .A3(KEYINPUT11), .ZN(new_n321));
  AND4_X1   g0121(.A1(new_n316), .A2(new_n318), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT71), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT71), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n325), .A2(G33), .A3(G97), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n215), .A2(new_n247), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n226), .A2(G1698), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n328), .B(new_n329), .C1(new_n253), .C2(new_n254), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n243), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n267), .A2(G238), .ZN(new_n335));
  NAND4_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n262), .A4(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n243), .B1(new_n327), .B2(new_n330), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n262), .B1(new_n217), .B2(new_n266), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT13), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n336), .A2(G190), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n322), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G200), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n336), .B2(new_n339), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT72), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n343), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(new_n340), .A4(new_n322), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n322), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n336), .A2(new_n339), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT14), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT73), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n350), .A2(G169), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT14), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT73), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n350), .A2(new_n356), .A3(new_n351), .A4(G169), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n336), .A2(G179), .A3(new_n339), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n353), .A2(new_n355), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n311), .B(new_n348), .C1(new_n349), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT17), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT8), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT67), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT67), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT8), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G58), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n367), .A2(KEYINPUT66), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n363), .A3(new_n365), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n317), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n274), .A2(new_n292), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n370), .A2(new_n371), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n373), .A2(new_n374), .B1(new_n292), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n246), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n255), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n216), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n367), .A2(new_n216), .ZN(new_n381));
  NOR2_X1   g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n280), .A2(G159), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n274), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n255), .B2(new_n210), .ZN(new_n388));
  NOR4_X1   g0188(.A1(new_n253), .A2(new_n254), .A3(new_n377), .A4(G20), .ZN(new_n389));
  OAI21_X1  g0189(.A(G68), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n383), .A2(new_n384), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n387), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n376), .B1(new_n386), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  OR2_X1    g0195(.A1(G223), .A2(G1698), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n215), .A2(G1698), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n396), .B(new_n397), .C1(new_n253), .C2(new_n254), .ZN(new_n398));
  NAND2_X1  g0198(.A1(G33), .A2(G87), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n395), .B1(new_n400), .B2(new_n332), .ZN(new_n401));
  AOI211_X1 g0201(.A(KEYINPUT75), .B(new_n243), .C1(new_n398), .C2(new_n399), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n243), .A2(G232), .A3(new_n265), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n262), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G190), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n400), .A2(new_n332), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n405), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n403), .A2(new_n407), .B1(new_n342), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n361), .B1(new_n394), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n375), .A2(new_n292), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n288), .A2(new_n289), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n372), .ZN(new_n414));
  INV_X1    g0214(.A(new_n387), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n380), .B2(new_n391), .ZN(new_n416));
  INV_X1    g0216(.A(new_n385), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n288), .B1(new_n390), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n414), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g0219(.A1(G223), .A2(G1698), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n215), .B2(G1698), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n421), .A2(new_n246), .B1(G33), .B2(G87), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT75), .B1(new_n422), .B2(new_n243), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n400), .A2(new_n395), .A3(new_n332), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(new_n406), .A3(new_n405), .A4(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n409), .A2(new_n342), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n419), .A2(new_n427), .A3(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n411), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(G169), .B1(new_n408), .B2(new_n405), .ZN(new_n430));
  AND3_X1   g0230(.A1(new_n262), .A2(new_n404), .A3(new_n299), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n430), .B1(new_n403), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT18), .B1(new_n394), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n394), .A2(KEYINPUT18), .A3(new_n432), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(KEYINPUT76), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT76), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n394), .A2(new_n432), .A3(new_n436), .A4(KEYINPUT18), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n429), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n214), .A2(new_n367), .A3(new_n216), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(G20), .B1(G150), .B2(new_n280), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n375), .B2(new_n276), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n441), .A2(new_n274), .B1(new_n214), .B2(new_n292), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n374), .A2(G50), .A3(new_n317), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n246), .A2(G222), .A3(new_n247), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n246), .A2(G223), .A3(G1698), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n255), .A2(G77), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT64), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT64), .A4(new_n448), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n332), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n263), .B1(G226), .B2(new_n267), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n445), .B1(new_n241), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n299), .A3(new_n454), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT9), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n444), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n455), .A2(G200), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n453), .A2(G190), .A3(new_n454), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n442), .A2(KEYINPUT9), .A3(new_n443), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n460), .A2(new_n461), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT10), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n464), .A2(KEYINPUT10), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n458), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n360), .A2(new_n438), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT24), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT23), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n210), .B2(G107), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n301), .A2(KEYINPUT23), .A3(G20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G33), .ZN(new_n474));
  INV_X1    g0274(.A(G116), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n210), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n210), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n478));
  XNOR2_X1  g0278(.A(KEYINPUT79), .B(KEYINPUT22), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n473), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n469), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n479), .ZN(new_n483));
  AOI21_X1  g0283(.A(G20), .B1(new_n244), .B2(new_n245), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n483), .A2(new_n484), .A3(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n478), .A2(new_n479), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n471), .A2(new_n472), .B1(new_n476), .B2(new_n210), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT24), .A4(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n482), .A2(new_n274), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n264), .A2(new_n301), .A3(G13), .A4(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT25), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n264), .A2(G33), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n289), .B(new_n494), .C1(new_n272), .C2(new_n273), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n490), .B(new_n493), .C1(new_n495), .C2(new_n301), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n288), .A2(G107), .A3(new_n289), .A4(new_n494), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n490), .B1(new_n498), .B2(new_n493), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n489), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT5), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G41), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n264), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(KEYINPUT77), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n501), .A2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT77), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n264), .A4(G45), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n332), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(G257), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(new_n247), .C1(new_n253), .C2(new_n254), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n508), .A2(G264), .B1(new_n332), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G274), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n332), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n504), .A3(new_n507), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n299), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n516), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n241), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n500), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n493), .B1(new_n495), .B2(new_n301), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT80), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n496), .ZN(new_n524));
  AOI21_X1  g0324(.A(G200), .B1(new_n513), .B2(new_n516), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n264), .A2(G45), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT77), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n502), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n507), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(G264), .A3(new_n243), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n512), .A2(new_n332), .ZN(new_n532));
  AND4_X1   g0332(.A1(new_n406), .A2(new_n531), .A3(new_n516), .A4(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n524), .B(new_n489), .C1(new_n525), .C2(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n520), .A2(new_n521), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n521), .B1(new_n520), .B2(new_n534), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n530), .A2(G270), .A3(new_n243), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT78), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n528), .A2(new_n507), .A3(new_n529), .ZN(new_n540));
  OAI211_X1 g0340(.A(G264), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(new_n247), .C1(new_n253), .C2(new_n254), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n244), .A2(G303), .A3(new_n245), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n540), .A2(new_n515), .B1(new_n544), .B2(new_n332), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n508), .A2(new_n546), .A3(G270), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n539), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  INV_X1    g0350(.A(G97), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n210), .C1(G33), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n475), .A2(G20), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n284), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n284), .A3(KEYINPUT20), .A4(new_n553), .ZN(new_n557));
  INV_X1    g0357(.A(G13), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(G1), .ZN(new_n559));
  INV_X1    g0359(.A(new_n553), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n556), .A2(new_n557), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n288), .A2(G116), .A3(new_n289), .A4(new_n494), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n539), .A2(new_n545), .A3(G190), .A4(new_n547), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n549), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g0366(.A1(new_n539), .A2(new_n545), .A3(new_n547), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(G179), .A3(new_n563), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n241), .B1(new_n561), .B2(new_n562), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n548), .B2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n548), .A2(new_n569), .A3(new_n570), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n566), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(G97), .A2(G107), .ZN(new_n574));
  INV_X1    g0374(.A(G87), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n324), .B2(new_n326), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n578), .B2(G20), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n484), .A2(G68), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n288), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n495), .A2(new_n275), .ZN(new_n583));
  INV_X1    g0383(.A(new_n275), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(new_n289), .ZN(new_n585));
  OR3_X1    g0385(.A1(new_n582), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G250), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n260), .B2(G1), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n264), .A2(new_n514), .A3(G45), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n243), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n591));
  OAI211_X1 g0391(.A(G238), .B(new_n247), .C1(new_n253), .C2(new_n254), .ZN(new_n592));
  INV_X1    g0392(.A(new_n476), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n590), .B1(new_n594), .B2(new_n332), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G179), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n241), .B2(new_n595), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n406), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(G200), .B2(new_n595), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n495), .A2(new_n575), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n582), .A2(new_n600), .A3(new_n585), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n586), .A2(new_n597), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g0402(.A1(KEYINPUT4), .A2(G244), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n247), .B(new_n603), .C1(new_n253), .C2(new_n254), .ZN(new_n604));
  INV_X1    g0404(.A(G244), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n244), .B2(new_n245), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n604), .B(new_n550), .C1(new_n606), .C2(KEYINPUT4), .ZN(new_n607));
  OAI21_X1  g0407(.A(G250), .B1(new_n253), .B2(new_n254), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n247), .B1(new_n608), .B2(KEYINPUT4), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n332), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n508), .A2(G257), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n516), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n241), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT6), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n614), .A2(new_n551), .A3(G107), .ZN(new_n615));
  XNOR2_X1  g0415(.A(G97), .B(G107), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n615), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI22_X1  g0417(.A1(new_n617), .A2(new_n210), .B1(new_n277), .B2(new_n281), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n301), .B1(new_n378), .B2(new_n379), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n274), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n289), .A2(G97), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n622), .B1(new_n495), .B2(new_n551), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n613), .B(new_n625), .C1(G179), .C2(new_n612), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n612), .A2(G200), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n551), .A2(new_n301), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n614), .B1(new_n628), .B2(new_n574), .ZN(new_n629));
  INV_X1    g0429(.A(new_n615), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n631), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n632));
  OAI21_X1  g0432(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n623), .B1(new_n634), .B2(new_n274), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n627), .B(new_n635), .C1(new_n406), .C2(new_n612), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n602), .A2(new_n626), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n573), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n468), .A2(new_n537), .A3(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n586), .A2(new_n597), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n599), .A2(new_n601), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NOR3_X1   g0444(.A1(new_n643), .A2(new_n626), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n641), .B1(new_n645), .B2(KEYINPUT82), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n520), .B(new_n568), .C1(new_n571), .C2(new_n572), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n626), .A2(new_n636), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n647), .A2(new_n648), .A3(new_n534), .A4(new_n602), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n643), .B2(new_n626), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n610), .A2(new_n611), .A3(new_n516), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n635), .B1(new_n299), .B2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n602), .A2(new_n652), .A3(KEYINPUT26), .A4(new_n613), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT82), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n650), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n646), .A2(new_n649), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n468), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT18), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n423), .A2(new_n424), .A3(new_n431), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n409), .A2(new_n241), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n419), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n434), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n344), .A2(new_n347), .ZN(new_n664));
  INV_X1    g0464(.A(new_n305), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n359), .B2(new_n349), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n429), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n464), .B(KEYINPUT10), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n458), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n657), .A2(new_n669), .ZN(G369));
  OAI21_X1  g0470(.A(new_n568), .B1(new_n572), .B2(new_n571), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n559), .A2(new_n210), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(G213), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n564), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n671), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n573), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n500), .A2(new_n677), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n537), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n520), .A2(new_n678), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n677), .B(KEYINPUT83), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n520), .A2(new_n690), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n671), .A2(new_n678), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n537), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n688), .A2(new_n693), .ZN(G399));
  NOR2_X1   g0494(.A1(new_n576), .A2(G116), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n204), .A2(new_n259), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n207), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n647), .A2(new_n648), .A3(new_n534), .A4(new_n642), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n641), .B1(new_n650), .B2(new_n653), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n677), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n656), .A2(new_n689), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(KEYINPUT29), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n689), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n595), .A2(G179), .A3(new_n531), .A4(new_n532), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n567), .A2(new_n709), .A3(KEYINPUT30), .A4(new_n651), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT85), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n548), .A2(new_n612), .A3(new_n708), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT85), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  AOI22_X1  g0516(.A1(G257), .A2(new_n508), .B1(new_n540), .B2(new_n515), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n299), .B(new_n590), .C1(new_n594), .C2(new_n332), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n717), .A2(new_n718), .A3(new_n513), .A4(new_n610), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n716), .B1(new_n719), .B2(new_n548), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n595), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n548), .A2(new_n518), .A3(new_n612), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT84), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n723), .A2(KEYINPUT84), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n707), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n537), .A2(new_n638), .A3(new_n689), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n723), .B1(new_n714), .B2(new_n711), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n706), .B1(new_n729), .B2(new_n678), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G330), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n705), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n699), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(new_n558), .A2(G20), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n264), .B1(new_n736), .B2(G45), .ZN(new_n737));
  AND2_X1   g0537(.A1(new_n737), .A2(new_n696), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT86), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n209), .B1(G20), .B2(new_n241), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n299), .A2(new_n342), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT89), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n210), .A2(G190), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G159), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT32), .Z(new_n749));
  OAI21_X1  g0549(.A(G20), .B1(new_n744), .B2(new_n406), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G97), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n210), .A2(new_n406), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n299), .A2(G200), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XOR2_X1   g0554(.A(new_n754), .B(KEYINPUT88), .Z(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G58), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n210), .A2(new_n299), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n758), .A2(new_n406), .A3(G200), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n759), .A2(new_n216), .B1(new_n760), .B2(new_n214), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n342), .A2(G179), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n745), .A2(new_n762), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n575), .B1(new_n764), .B2(new_n301), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n745), .A2(new_n753), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n246), .B1(new_n766), .B2(new_n277), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n761), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n749), .A2(new_n751), .A3(new_n757), .A4(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n763), .ZN(new_n770));
  INV_X1    g0570(.A(new_n754), .ZN(new_n771));
  AOI22_X1  g0571(.A1(G303), .A2(new_n770), .B1(new_n771), .B2(G322), .ZN(new_n772));
  INV_X1    g0572(.A(G283), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n764), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G329), .B2(new_n747), .ZN(new_n775));
  INV_X1    g0575(.A(new_n759), .ZN(new_n776));
  NOR2_X1   g0576(.A1(KEYINPUT33), .A2(G317), .ZN(new_n777));
  AND2_X1   g0577(.A1(KEYINPUT33), .A2(G317), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n766), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n246), .B1(new_n780), .B2(G311), .ZN(new_n781));
  INV_X1    g0581(.A(new_n760), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G326), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G294), .ZN(new_n785));
  INV_X1    g0585(.A(new_n750), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n775), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n742), .B1(new_n769), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT87), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(G20), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n741), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n255), .A2(new_n204), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n260), .B2(new_n208), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n236), .B2(new_n260), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n246), .A2(new_n204), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n795), .B1(G116), .B2(new_n204), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  AOI211_X1 g0598(.A(new_n740), .B(new_n788), .C1(new_n792), .C2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT90), .ZN(new_n800));
  INV_X1    g0600(.A(new_n791), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n681), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n683), .A2(new_n739), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(G330), .B2(new_n681), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G396));
  NAND2_X1  g0606(.A1(new_n298), .A2(new_n677), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n309), .B2(new_n310), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n305), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n305), .A2(new_n677), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n704), .B(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n739), .B1(new_n814), .B2(new_n732), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n732), .B2(new_n814), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n782), .A2(G137), .B1(new_n780), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  INV_X1    g0618(.A(G143), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n759), .C1(new_n755), .C2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT34), .Z(new_n821));
  OAI221_X1 g0621(.A(new_n246), .B1(new_n764), .B2(new_n216), .C1(new_n214), .C2(new_n763), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G132), .B2(new_n747), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n367), .B2(new_n786), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n751), .B1(new_n785), .B2(new_n754), .ZN(new_n825));
  XOR2_X1   g0625(.A(new_n825), .B(KEYINPUT94), .Z(new_n826));
  AOI22_X1  g0626(.A1(new_n776), .A2(G283), .B1(new_n780), .B2(G116), .ZN(new_n827));
  INV_X1    g0627(.A(G303), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n760), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(KEYINPUT92), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n255), .B1(new_n763), .B2(new_n301), .ZN(new_n831));
  XOR2_X1   g0631(.A(new_n831), .B(KEYINPUT93), .Z(new_n832));
  INV_X1    g0632(.A(new_n764), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n747), .A2(G311), .B1(G87), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n830), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n821), .A2(new_n824), .B1(new_n826), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n742), .B1(new_n836), .B2(KEYINPUT95), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(KEYINPUT95), .B2(new_n836), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n741), .A2(new_n789), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT91), .Z(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n740), .B1(new_n277), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n838), .B(new_n842), .C1(new_n790), .C2(new_n813), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n816), .A2(new_n843), .ZN(G384));
  AOI22_X1  g0644(.A1(new_n419), .A2(new_n427), .B1(KEYINPUT97), .B2(KEYINPUT37), .ZN(new_n845));
  INV_X1    g0645(.A(new_n675), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n394), .B1(new_n432), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(KEYINPUT97), .A2(KEYINPUT37), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n845), .B2(new_n847), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n419), .A2(new_n675), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n438), .B2(new_n855), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n411), .A2(new_n428), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(new_n663), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n845), .A2(new_n847), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n848), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n856), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n434), .A2(KEYINPUT76), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(new_n437), .A3(new_n662), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n857), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n854), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(KEYINPUT98), .A3(new_n853), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT98), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n855), .B1(new_n867), .B2(new_n857), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n850), .A2(new_n851), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n438), .B2(new_n855), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n870), .A2(new_n874), .B1(new_n876), .B2(new_n852), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n865), .B1(new_n877), .B2(new_n864), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n359), .A2(new_n349), .A3(new_n678), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT99), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n663), .A2(new_n846), .ZN(new_n883));
  OAI211_X1 g0683(.A(new_n349), .B(new_n677), .C1(new_n348), .C2(new_n359), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n359), .A2(new_n349), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n322), .A2(new_n678), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n664), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n656), .A2(new_n689), .A3(new_n813), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n810), .B(KEYINPUT96), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n876), .A2(new_n852), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT98), .B1(new_n869), .B2(new_n853), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n872), .A2(new_n873), .A3(new_n871), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n883), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n881), .A2(new_n882), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n882), .B1(new_n881), .B2(new_n899), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n468), .B(new_n703), .C1(new_n704), .C2(KEYINPUT29), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n669), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n902), .B(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n711), .A2(new_n714), .ZN(new_n906));
  OAI211_X1 g0706(.A(KEYINPUT31), .B(new_n677), .C1(new_n906), .C2(new_n723), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n728), .A2(new_n730), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n812), .B1(new_n884), .B2(new_n888), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n898), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT100), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n908), .A2(new_n909), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n872), .A2(new_n873), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n419), .A2(new_n661), .A3(new_n658), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(new_n433), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n854), .B1(new_n916), .B2(new_n429), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT38), .B1(new_n875), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT40), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n912), .B1(new_n913), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n911), .B1(new_n856), .B2(new_n863), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(KEYINPUT100), .A3(new_n908), .A4(new_n909), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n910), .A2(new_n911), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(new_n468), .A3(new_n908), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(G330), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n923), .B1(new_n468), .B2(new_n908), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n905), .A2(new_n927), .B1(new_n264), .B2(new_n736), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT101), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n905), .A2(new_n927), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n631), .A2(KEYINPUT35), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n631), .A2(KEYINPUT35), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n934), .A2(G116), .A3(new_n211), .A4(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n381), .A2(new_n207), .A3(new_n277), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n216), .A2(G50), .ZN(new_n939));
  OAI211_X1 g0739(.A(G1), .B(new_n558), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n933), .A2(new_n937), .A3(new_n940), .ZN(G367));
  OAI21_X1  g0741(.A(new_n636), .B1(new_n635), .B2(new_n689), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n626), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n537), .A2(new_n692), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n652), .A2(new_n613), .A3(new_n689), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n691), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n945), .B(new_n946), .C1(new_n693), .C2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n601), .A2(new_n678), .ZN(new_n953));
  MUX2_X1   g0753(.A(new_n602), .B(new_n641), .S(new_n953), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT104), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(KEYINPUT102), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n954), .A2(KEYINPUT102), .ZN(new_n960));
  XOR2_X1   g0760(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  OR3_X1    g0762(.A1(new_n959), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n956), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(KEYINPUT104), .B2(new_n963), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n688), .A2(new_n947), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n956), .A2(new_n957), .A3(new_n964), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n966), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n967), .B1(new_n966), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n696), .B(KEYINPUT41), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n687), .A2(new_n692), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n537), .A2(new_n692), .ZN(new_n974));
  AND3_X1   g0774(.A1(new_n973), .A2(new_n682), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n682), .B1(new_n973), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n977), .A2(new_n733), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n693), .A2(new_n948), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT45), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n974), .A2(new_n949), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT105), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(new_n947), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT105), .B1(new_n693), .B2(new_n948), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT44), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n983), .A2(KEYINPUT44), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n980), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n688), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n980), .A2(new_n987), .A3(new_n688), .A4(new_n988), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n978), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n972), .B1(new_n993), .B2(new_n734), .ZN(new_n994));
  INV_X1    g0794(.A(new_n737), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n971), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n792), .B1(new_n204), .B2(new_n275), .C1(new_n232), .C2(new_n793), .ZN(new_n997));
  AND2_X1   g0797(.A1(new_n997), .A2(new_n739), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n246), .B1(new_n766), .B2(new_n214), .C1(new_n760), .C2(new_n819), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G159), .B2(new_n776), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n750), .A2(G68), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(KEYINPUT106), .B(G137), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n747), .A2(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n367), .A2(new_n763), .B1(new_n754), .B2(new_n818), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G77), .B2(new_n833), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n764), .A2(new_n551), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n246), .B(new_n1007), .C1(G283), .C2(new_n780), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n747), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1008), .B1(new_n828), .B2(new_n755), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n763), .A2(new_n475), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1012), .A2(KEYINPUT46), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G294), .B2(new_n776), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n1012), .A2(KEYINPUT46), .B1(new_n782), .B2(G311), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n786), .C2(new_n301), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1006), .B1(new_n1011), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT47), .Z(new_n1018));
  OAI221_X1 g0818(.A(new_n998), .B1(new_n801), .B2(new_n954), .C1(new_n1018), .C2(new_n742), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n996), .A2(new_n1019), .ZN(G387));
  XNOR2_X1  g0820(.A(new_n696), .B(KEYINPUT112), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT113), .B1(new_n978), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n734), .B1(new_n976), .B2(new_n975), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT113), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n1025), .A3(new_n1021), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n977), .A2(new_n733), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OR3_X1    g0828(.A1(new_n977), .A2(KEYINPUT107), .A3(new_n737), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT107), .B1(new_n977), .B2(new_n737), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n685), .A2(new_n686), .A3(new_n791), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n782), .A2(G322), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n776), .A2(G311), .B1(new_n780), .B2(G303), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n755), .C2(new_n1009), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT48), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n750), .A2(G283), .B1(G294), .B2(new_n770), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n255), .B1(new_n764), .B2(new_n475), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n747), .B2(G326), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n750), .A2(new_n584), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n214), .B2(new_n754), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT110), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n375), .A2(new_n759), .B1(new_n216), .B2(new_n766), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT111), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n255), .B(new_n1007), .C1(G77), .C2(new_n770), .ZN(new_n1051));
  INV_X1    g0851(.A(G159), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1051), .B1(new_n1052), .B2(new_n760), .C1(new_n818), .C2(new_n1010), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n1048), .A2(new_n1050), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n742), .B1(new_n1045), .B2(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n797), .A2(new_n695), .B1(G107), .B2(new_n204), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n229), .A2(new_n260), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT108), .Z(new_n1058));
  INV_X1    g0858(.A(new_n695), .ZN(new_n1059));
  AOI211_X1 g0859(.A(G45), .B(new_n1059), .C1(G68), .C2(G77), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n279), .A2(G50), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1061), .B(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n793), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1056), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n792), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n739), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1055), .A2(new_n1067), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n1029), .A2(new_n1030), .B1(new_n1031), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1028), .A2(new_n1069), .ZN(G393));
  NAND3_X1  g0870(.A1(new_n991), .A2(new_n995), .A3(new_n992), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n792), .B1(new_n551), .B2(new_n204), .C1(new_n239), .C2(new_n793), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n739), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n747), .A2(G322), .B1(G283), .B2(new_n770), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT116), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n782), .A2(G317), .B1(new_n771), .B2(G311), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n255), .B1(new_n766), .B2(new_n785), .C1(new_n301), .C2(new_n764), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G303), .B2(new_n776), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1078), .B(new_n1080), .C1(new_n475), .C2(new_n786), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n763), .A2(new_n216), .B1(new_n766), .B2(new_n279), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n255), .B(new_n1082), .C1(G87), .C2(new_n833), .ZN(new_n1083));
  OAI221_X1 g0883(.A(new_n1083), .B1(new_n214), .B2(new_n759), .C1(new_n819), .C2(new_n1010), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n760), .A2(new_n818), .B1(new_n754), .B2(new_n1052), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n750), .A2(G77), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n1075), .A2(new_n1081), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1073), .B1(new_n1090), .B2(new_n741), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n948), .B2(new_n801), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1071), .A2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n993), .A2(new_n1021), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n991), .A2(new_n992), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1024), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(G390));
  AOI21_X1  g0898(.A(new_n892), .B1(new_n702), .B2(new_n813), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n879), .B1(new_n914), .B2(new_n918), .C1(new_n1099), .C2(new_n890), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n891), .A2(new_n893), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n880), .B1(new_n1101), .B2(new_n889), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1102), .B2(new_n878), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n908), .A2(G330), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1104), .A2(new_n812), .A3(new_n890), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1105), .A2(KEYINPUT117), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n731), .A2(G330), .A3(new_n813), .A4(new_n889), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n908), .A2(new_n909), .A3(new_n1110), .A4(G330), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1112), .B(new_n1100), .C1(new_n878), .C2(new_n1102), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1107), .A2(new_n995), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n740), .B1(new_n375), .B2(new_n841), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n255), .B1(new_n763), .B2(new_n575), .C1(new_n773), .C2(new_n760), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G107), .B2(new_n776), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n747), .A2(G294), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n754), .A2(new_n475), .B1(new_n764), .B2(new_n216), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G97), .B2(new_n780), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1088), .A3(new_n1118), .A4(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n770), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT53), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n763), .B2(new_n818), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n747), .A2(G125), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n255), .B1(new_n833), .B2(G50), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n766), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G132), .B2(new_n771), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1002), .A2(new_n776), .B1(new_n782), .B2(G128), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1125), .A2(new_n1126), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n786), .A2(new_n1052), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1121), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1133), .A2(KEYINPUT118), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(KEYINPUT118), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n741), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n1115), .B1(new_n1134), .B2(new_n1136), .C1(new_n878), .C2(new_n790), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1104), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n468), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n903), .A2(new_n1139), .A3(new_n669), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n890), .B1(new_n1104), .B2(new_n812), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n1099), .A3(new_n1108), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n731), .A2(G330), .A3(new_n813), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1138), .A2(new_n909), .B1(new_n1144), .B2(new_n890), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1101), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1107), .A2(new_n1113), .A3(new_n1141), .A4(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n1021), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1144), .A2(new_n890), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1101), .B1(new_n1150), .B2(new_n1105), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1140), .B1(new_n1151), .B2(new_n1143), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n1113), .B2(new_n1107), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1114), .B(new_n1137), .C1(new_n1149), .C2(new_n1153), .ZN(G378));
  NAND3_X1  g0954(.A1(new_n881), .A2(new_n882), .A3(new_n899), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n920), .A2(new_n922), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n911), .B1(new_n877), .B2(new_n913), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(G330), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n458), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n668), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n444), .A2(new_n846), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT120), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n467), .A2(new_n1162), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g0966(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1158), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n879), .B1(new_n1174), .B2(new_n865), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n898), .A2(new_n1101), .A3(new_n889), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n883), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT99), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1156), .A2(new_n1171), .A3(G330), .A4(new_n1157), .ZN(new_n1180));
  AND4_X1   g0980(.A1(new_n1155), .A2(new_n1173), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1180), .A2(new_n1173), .B1(new_n1179), .B2(new_n1155), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n995), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n739), .B1(new_n840), .B2(G50), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(G33), .A2(G41), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT119), .ZN(new_n1186));
  AOI211_X1 g0986(.A(G50), .B(new_n1186), .C1(new_n259), .C2(new_n255), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G41), .B(new_n246), .C1(new_n770), .C2(G77), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n475), .B2(new_n760), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(G97), .B2(new_n776), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n584), .A2(new_n780), .B1(new_n833), .B2(G58), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n301), .B2(new_n754), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G283), .B2(new_n747), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1001), .A3(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT58), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1187), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(G137), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n763), .A2(new_n1127), .B1(new_n766), .B2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G128), .B2(new_n771), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n776), .A2(G132), .B1(new_n782), .B2(G125), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1199), .B(new_n1200), .C1(new_n786), .C2(new_n818), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1186), .B1(new_n1052), .B2(new_n764), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n747), .B2(G124), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1196), .B1(new_n1195), .B2(new_n1194), .C1(new_n1202), .C2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1184), .B1(new_n1207), .B2(new_n741), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n1172), .B2(new_n790), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1183), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1171), .B1(new_n923), .B2(G330), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1180), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1211), .A2(new_n1212), .B1(new_n900), .B2(new_n901), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1173), .A2(new_n1179), .A3(new_n1155), .A4(new_n1180), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1148), .A2(new_n1141), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT57), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1148), .B2(new_n1141), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1022), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1210), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(G375));
  NOR2_X1   g1023(.A1(new_n1147), .A2(new_n1141), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1224), .A2(new_n1152), .A3(new_n972), .ZN(new_n1225));
  XNOR2_X1  g1025(.A(new_n1225), .B(KEYINPUT121), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n255), .B1(new_n764), .B2(new_n277), .C1(new_n759), .C2(new_n475), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G294), .B2(new_n782), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n747), .A2(G303), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n763), .A2(new_n551), .B1(new_n766), .B2(new_n301), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G283), .B2(new_n771), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1228), .A2(new_n1046), .A3(new_n1229), .A4(new_n1231), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n756), .A2(new_n1002), .B1(G128), .B2(new_n747), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n763), .A2(new_n1052), .B1(new_n766), .B2(new_n818), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n255), .B(new_n1234), .C1(G58), .C2(new_n833), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1233), .B(new_n1235), .C1(new_n759), .C2(new_n1127), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n782), .A2(G132), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1237), .B(KEYINPUT123), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n214), .B2(new_n786), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1232), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(new_n741), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1241), .B(new_n739), .C1(G68), .C2(new_n840), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n890), .B2(new_n789), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n737), .B(KEYINPUT122), .Z(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1243), .B1(new_n1147), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1226), .A2(new_n1246), .ZN(G381));
  OR4_X1    g1047(.A1(G396), .A2(G378), .A3(G393), .A4(G384), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1097), .A2(new_n996), .A3(new_n1019), .ZN(new_n1249));
  OR4_X1    g1049(.A1(G375), .A2(new_n1248), .A3(G381), .A4(new_n1249), .ZN(G407));
  INV_X1    g1050(.A(G378), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1222), .A2(new_n676), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(G407), .A2(G213), .A3(new_n1252), .ZN(G409));
  INV_X1    g1053(.A(new_n1209), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n1215), .B2(new_n995), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1215), .A2(new_n1220), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1021), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT57), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G378), .B(new_n1255), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n972), .B1(new_n1148), .B2(new_n1141), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1215), .B1(new_n1260), .B2(new_n1245), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1209), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1251), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n676), .A2(G213), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT60), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n1147), .B2(new_n1141), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1268), .B2(new_n1224), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1151), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1270));
  OAI211_X1 g1070(.A(KEYINPUT124), .B(new_n1270), .C1(new_n1152), .C2(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1022), .B1(new_n1224), .B2(KEYINPUT60), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1269), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1273), .A2(G384), .A3(new_n1246), .ZN(new_n1274));
  AOI21_X1  g1074(.A(G384), .B1(new_n1273), .B2(new_n1246), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1264), .A2(new_n1265), .A3(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(KEYINPUT127), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1273), .A2(new_n1246), .ZN(new_n1281));
  INV_X1    g1081(.A(G384), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1273), .A2(G384), .A3(new_n1246), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1265), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(KEYINPUT126), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(G2897), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1276), .A2(new_n1288), .A3(new_n1286), .ZN(new_n1291));
  AOI21_X1  g1091(.A(G378), .B1(new_n1261), .B2(new_n1209), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1222), .B2(G378), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1290), .B(new_n1291), .C1(new_n1293), .C2(new_n1285), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1264), .A2(new_n1265), .A3(new_n1276), .A4(new_n1296), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1280), .A2(new_n1294), .A3(new_n1295), .A4(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(G393), .B(new_n805), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1249), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1097), .B1(new_n996), .B2(new_n1019), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(G393), .B(G396), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(G390), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1249), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1298), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1286), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1274), .A2(new_n1275), .A3(new_n1308), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(new_n1264), .A2(new_n1265), .B1(new_n1309), .B2(new_n1288), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1310), .B2(new_n1290), .ZN(new_n1311));
  AND2_X1   g1111(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1312));
  XOR2_X1   g1112(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n1313));
  NAND2_X1  g1113(.A1(new_n1277), .A2(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1264), .A2(KEYINPUT63), .A3(new_n1265), .A4(new_n1276), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1311), .A2(new_n1312), .A3(new_n1314), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1307), .A2(new_n1316), .ZN(G405));
  NAND2_X1  g1117(.A1(G375), .A2(new_n1251), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1259), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1312), .A2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1306), .A2(new_n1318), .A3(new_n1259), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1276), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1320), .A2(new_n1276), .A3(new_n1321), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(G402));
endmodule


