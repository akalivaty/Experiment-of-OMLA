//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  NAND2_X1  g000(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n187));
  XNOR2_X1  g001(.A(G125), .B(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(G146), .A3(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT23), .B1(new_n198), .B2(G119), .ZN(new_n199));
  AOI21_X1  g013(.A(KEYINPUT72), .B1(new_n198), .B2(G119), .ZN(new_n200));
  XNOR2_X1  g014(.A(new_n199), .B(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G110), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT24), .B(G110), .Z(new_n203));
  XNOR2_X1  g017(.A(G119), .B(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n197), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n201), .A2(G110), .B1(new_n204), .B2(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n188), .A2(new_n194), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n196), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G137), .ZN(new_n211));
  INV_X1    g025(.A(G221), .ZN(new_n212));
  INV_X1    g026(.A(G234), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n212), .A2(new_n213), .A3(G953), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n211), .B(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n210), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G902), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n187), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n210), .A2(new_n216), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n215), .B1(new_n206), .B2(new_n209), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n218), .B(new_n187), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n219), .A2(new_n223), .B1(KEYINPUT73), .B2(KEYINPUT25), .ZN(new_n224));
  OAI21_X1  g038(.A(G217), .B1(new_n213), .B2(G902), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT71), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G902), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n224), .A2(new_n226), .B1(new_n217), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G472), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n194), .A2(KEYINPUT65), .A3(G143), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G146), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n233), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT1), .B1(new_n232), .B2(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n240), .B(KEYINPUT1), .C1(new_n232), .C2(G146), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n198), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G143), .B(G146), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n237), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G134), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G137), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(G137), .ZN(new_n248));
  OAI21_X1  g062(.A(G131), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n250), .B1(new_n245), .B2(G137), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  INV_X1    g067(.A(G131), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .A4(new_n246), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n244), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G119), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT67), .B(G116), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n260), .B1(new_n261), .B2(G119), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT2), .B(G113), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n251), .A2(new_n253), .A3(new_n246), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G131), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n255), .ZN(new_n267));
  AND2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT0), .B(G128), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT64), .B1(new_n243), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n194), .A2(G143), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n236), .ZN(new_n273));
  NOR2_X1   g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT64), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n267), .A2(new_n269), .A3(new_n271), .A4(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n258), .A2(new_n264), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n283));
  AOI211_X1 g097(.A(new_n283), .B(new_n264), .C1(new_n258), .C2(new_n278), .ZN(new_n284));
  INV_X1    g098(.A(new_n237), .ZN(new_n285));
  INV_X1    g099(.A(new_n241), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n240), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n287));
  OAI21_X1  g101(.A(G128), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n288), .B2(new_n273), .ZN(new_n289));
  AND2_X1   g103(.A1(new_n266), .A2(new_n255), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n271), .A2(new_n269), .A3(new_n277), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n289), .A2(new_n256), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G116), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n295), .A3(G119), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n296), .B1(new_n259), .B2(G119), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n263), .ZN(new_n298));
  INV_X1    g112(.A(new_n263), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n262), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT69), .B1(new_n292), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n279), .B1(new_n284), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n282), .B1(new_n303), .B2(KEYINPUT28), .ZN(new_n304));
  NOR2_X1   g118(.A1(G237), .A2(G953), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G210), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT27), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT26), .B(G101), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT29), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n304), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT68), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n279), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n264), .B1(new_n258), .B2(new_n278), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT28), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n291), .ZN(new_n318));
  AOI22_X1  g132(.A1(new_n318), .A2(new_n267), .B1(new_n244), .B2(new_n257), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n319), .A2(new_n314), .A3(new_n264), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n309), .B(new_n281), .C1(new_n317), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n258), .A2(new_n322), .A3(new_n278), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n322), .B1(new_n258), .B2(new_n278), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n301), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n279), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n310), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n327), .A3(new_n311), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n230), .B1(new_n313), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n329), .B(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n325), .A2(new_n309), .A3(new_n279), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT31), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n325), .A2(KEYINPUT31), .A3(new_n309), .A4(new_n279), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n281), .B1(new_n317), .B2(new_n320), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n310), .ZN(new_n338));
  AOI21_X1  g152(.A(G902), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n230), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT32), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT32), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n342), .A3(new_n230), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n229), .B1(new_n331), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G214), .B1(G237), .B2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G110), .B(G122), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(G107), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT4), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G101), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(G101), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n350), .A2(new_n353), .A3(new_n359), .A4(new_n354), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(KEYINPUT4), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n301), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n260), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(G113), .B(new_n364), .C1(new_n297), .C2(new_n363), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n352), .A2(G104), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n349), .A2(G107), .ZN(new_n367));
  OAI21_X1  g181(.A(G101), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n365), .A2(new_n300), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n362), .A2(KEYINPUT76), .A3(new_n371), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n348), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n348), .A3(new_n371), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT6), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT77), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n348), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n362), .A2(KEYINPUT76), .A3(new_n371), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT76), .B1(new_n362), .B2(new_n371), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT77), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT6), .A4(new_n377), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n318), .A2(G125), .ZN(new_n386));
  INV_X1    g200(.A(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n244), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G224), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G953), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n389), .B(new_n391), .Z(new_n392));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n376), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n379), .A2(new_n385), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n389), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n391), .ZN(new_n397));
  AND2_X1   g211(.A1(KEYINPUT78), .A2(KEYINPUT7), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n389), .B1(KEYINPUT78), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n397), .A2(new_n398), .B1(new_n400), .B2(new_n391), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n399), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n348), .B(KEYINPUT8), .ZN(new_n403));
  INV_X1    g217(.A(new_n371), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n370), .B1(new_n365), .B2(new_n300), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n402), .A2(new_n406), .A3(new_n377), .ZN(new_n407));
  AOI21_X1  g221(.A(G902), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n395), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(new_n410), .A3(new_n408), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n347), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT15), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n198), .A2(G143), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n232), .A2(G128), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n245), .ZN(new_n420));
  OAI21_X1  g234(.A(G134), .B1(new_n417), .B2(new_n418), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n293), .A2(new_n295), .A3(G122), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n259), .A2(G122), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n352), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  OR2_X1    g240(.A1(new_n423), .A2(KEYINPUT14), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n423), .A2(KEYINPUT14), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n429), .B2(G107), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n232), .A2(KEYINPUT13), .A3(G128), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n198), .B2(G143), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n432), .B1(new_n434), .B2(new_n417), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n435), .A2(KEYINPUT82), .A3(G134), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT82), .B1(new_n435), .B2(G134), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n425), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n352), .B1(new_n423), .B2(new_n424), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n420), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n438), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n440), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n444), .A2(new_n425), .B1(new_n245), .B2(new_n419), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n435), .A2(G134), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n435), .A2(KEYINPUT82), .A3(G134), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT83), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n431), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT9), .B(G234), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G953), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n454), .A2(G217), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n442), .B1(new_n438), .B2(new_n441), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n445), .A2(new_n450), .A3(KEYINPUT83), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n430), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n456), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n416), .B1(new_n463), .B2(new_n218), .ZN(new_n464));
  INV_X1    g278(.A(new_n416), .ZN(new_n465));
  AOI211_X1 g279(.A(G902), .B(new_n465), .C1(new_n457), .C2(new_n462), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(G475), .A2(G902), .ZN(new_n468));
  XNOR2_X1  g282(.A(G113), .B(G122), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n469), .B(new_n349), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n471));
  AOI21_X1  g285(.A(G143), .B1(new_n305), .B2(G214), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n305), .A2(G214), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n232), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n305), .A2(G143), .A3(G214), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n254), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT17), .B(G131), .C1(new_n471), .C2(new_n472), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n195), .A4(new_n196), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n471), .A2(new_n472), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n387), .A2(G140), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n191), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G146), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n482), .A2(new_n483), .B1(new_n208), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT18), .B(G131), .C1(new_n471), .C2(new_n472), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT79), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n208), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n475), .A2(new_n476), .A3(new_n483), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT79), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n470), .B(new_n481), .C1(new_n489), .C2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n487), .A2(KEYINPUT79), .A3(new_n488), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n493), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n473), .A2(new_n477), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT80), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT80), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n473), .A2(new_n477), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT81), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n191), .A2(new_n484), .A3(new_n504), .A4(KEYINPUT19), .ZN(new_n505));
  XOR2_X1   g319(.A(KEYINPUT81), .B(KEYINPUT19), .Z(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n506), .B2(new_n188), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n194), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n501), .A2(new_n196), .A3(new_n503), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n470), .B1(new_n499), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n468), .B1(new_n496), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT20), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n503), .A2(new_n508), .A3(new_n196), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n513), .A2(new_n501), .B1(new_n497), .B2(new_n498), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n495), .B1(new_n514), .B2(new_n470), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n468), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n470), .B1(new_n499), .B2(new_n481), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n218), .B1(new_n496), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n512), .A2(new_n517), .B1(G475), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(G234), .A2(G237), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(G952), .A3(new_n455), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT21), .B(G898), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(KEYINPUT84), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n521), .A2(G902), .A3(G953), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n467), .A2(KEYINPUT85), .A3(new_n520), .A4(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT85), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n460), .A2(new_n461), .ZN(new_n529));
  AOI211_X1 g343(.A(new_n456), .B(new_n430), .C1(new_n458), .C2(new_n459), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n218), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n465), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n463), .A2(new_n218), .A3(new_n416), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n519), .A2(G475), .ZN(new_n535));
  INV_X1    g349(.A(new_n517), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n516), .B1(new_n515), .B2(new_n468), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n535), .B(new_n526), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n528), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n527), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n290), .A2(KEYINPUT74), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n233), .A2(new_n234), .A3(new_n236), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n198), .B1(new_n272), .B2(KEYINPUT1), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n237), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n370), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n369), .B(new_n237), .C1(new_n242), .C2(new_n243), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT75), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT75), .B1(new_n289), .B2(new_n369), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n318), .A2(new_n361), .A3(new_n357), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT10), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n244), .A2(KEYINPUT10), .A3(new_n370), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n552), .A2(new_n554), .A3(new_n555), .A4(new_n290), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G140), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n455), .A2(G227), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n558), .B(new_n559), .Z(new_n560));
  NAND3_X1  g374(.A1(new_n289), .A2(KEYINPUT75), .A3(new_n369), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n546), .A2(new_n547), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n545), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT74), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT12), .A4(new_n267), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n557), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n554), .A2(new_n555), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n318), .A2(new_n357), .A3(new_n361), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n267), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n560), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n556), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n566), .A2(new_n567), .A3(new_n218), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(G469), .A2(G902), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n557), .A2(new_n571), .A3(new_n565), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n570), .A2(new_n560), .A3(new_n556), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n573), .B(new_n574), .C1(new_n567), .C2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n212), .B1(new_n454), .B2(new_n218), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n414), .A2(new_n540), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n345), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  AOI22_X1  g399(.A1(new_n334), .A2(new_n335), .B1(new_n337), .B2(new_n310), .ZN(new_n586));
  OAI21_X1  g400(.A(G472), .B1(new_n586), .B2(G902), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n340), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(new_n229), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n582), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(KEYINPUT86), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n395), .A2(new_n410), .A3(new_n408), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n410), .B1(new_n395), .B2(new_n408), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n526), .B(new_n346), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT87), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n452), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n457), .A2(new_n596), .A3(KEYINPUT33), .A4(new_n462), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT33), .B1(new_n460), .B2(KEYINPUT87), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(new_n529), .B2(new_n530), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n597), .A2(new_n599), .A3(G478), .A4(new_n218), .ZN(new_n600));
  NOR2_X1   g414(.A1(KEYINPUT88), .A2(G478), .ZN(new_n601));
  AND2_X1   g415(.A1(KEYINPUT88), .A2(G478), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n531), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n520), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n594), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n591), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NAND2_X1  g424(.A1(new_n534), .A2(new_n520), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n594), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n591), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT89), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  INV_X1    g430(.A(new_n588), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n215), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n210), .B(new_n618), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n224), .A2(new_n226), .B1(new_n227), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n583), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT91), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT90), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G12));
  AND3_X1   g440(.A1(new_n321), .A2(new_n311), .A3(new_n327), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n283), .B1(new_n319), .B2(new_n264), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n316), .A2(KEYINPUT69), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n628), .A2(new_n629), .B1(new_n264), .B2(new_n319), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n281), .B(new_n312), .C1(new_n630), .C2(new_n280), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n218), .ZN(new_n632));
  OAI21_X1  g446(.A(G472), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n330), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n329), .A2(KEYINPUT70), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n342), .B1(new_n339), .B2(new_n230), .ZN(new_n636));
  NOR4_X1   g450(.A1(new_n586), .A2(KEYINPUT32), .A3(G472), .A4(G902), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n634), .B(new_n635), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n522), .B(KEYINPUT92), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n639), .B1(G900), .B2(new_n525), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT93), .Z(new_n641));
  NOR3_X1   g455(.A1(new_n581), .A2(new_n611), .A3(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n638), .A2(new_n414), .A3(new_n621), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  NAND2_X1  g458(.A1(new_n412), .A2(new_n413), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT38), .Z(new_n646));
  XOR2_X1   g460(.A(new_n641), .B(KEYINPUT39), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n582), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(G472), .A2(G902), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n332), .A2(G472), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n630), .A2(new_n309), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT94), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n344), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n648), .A2(KEYINPUT40), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n520), .B1(new_n532), .B2(new_n533), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n620), .A2(new_n658), .A3(new_n346), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n656), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n650), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT95), .B(G143), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G45));
  INV_X1    g477(.A(new_n641), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n604), .A2(new_n605), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n581), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n638), .A2(new_n666), .A3(new_n414), .A4(new_n621), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT96), .B(G146), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G48));
  NAND3_X1  g483(.A1(new_n566), .A2(new_n218), .A3(new_n572), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(G469), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n580), .A3(new_n573), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT97), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n607), .A2(new_n638), .A3(new_n228), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND4_X1  g491(.A1(new_n612), .A2(new_n638), .A3(new_n228), .A4(new_n674), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  AND2_X1   g493(.A1(new_n414), .A2(new_n540), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(new_n638), .A3(new_n621), .A4(new_n674), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G119), .ZN(G21));
  OAI211_X1 g496(.A(new_n658), .B(new_n346), .C1(new_n592), .C2(new_n593), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT100), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n645), .A2(new_n685), .A3(new_n346), .A4(new_n658), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(G472), .A2(G902), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n689), .B(KEYINPUT98), .Z(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n303), .A2(KEYINPUT28), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT99), .B1(new_n692), .B2(new_n281), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT99), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n694), .B(new_n282), .C1(new_n303), .C2(KEYINPUT28), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n310), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n691), .B1(new_n696), .B2(new_n336), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n339), .A2(new_n230), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n674), .A2(new_n699), .A3(new_n228), .A4(new_n526), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT101), .B1(new_n688), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n700), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n687), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NOR3_X1   g520(.A1(new_n697), .A2(new_n698), .A3(new_n620), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n512), .A2(new_n517), .ZN(new_n708));
  AOI221_X4 g522(.A(new_n641), .B1(new_n708), .B2(new_n535), .C1(new_n600), .C2(new_n603), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n707), .A2(new_n674), .A3(new_n414), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NAND3_X1  g525(.A1(new_n412), .A2(new_n346), .A3(new_n413), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n576), .A2(KEYINPUT102), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT102), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n570), .A2(new_n714), .A3(new_n560), .A4(new_n556), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n716), .A2(G469), .A3(new_n575), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n573), .A2(new_n574), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n580), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT103), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n716), .A2(G469), .A3(new_n575), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n573), .A3(new_n574), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n723), .A3(new_n580), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n712), .B1(new_n720), .B2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n228), .A3(new_n638), .A4(new_n709), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT42), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n345), .A2(KEYINPUT42), .A3(new_n709), .A4(new_n725), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G131), .ZN(G33));
  NOR2_X1   g545(.A1(new_n611), .A2(new_n641), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n725), .A2(new_n228), .A3(new_n638), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT104), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n345), .A2(new_n735), .A3(new_n732), .A4(new_n725), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT105), .B(G134), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G36));
  NAND3_X1  g553(.A1(new_n716), .A2(KEYINPUT45), .A3(new_n575), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n577), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(G469), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT46), .A3(new_n574), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n573), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT46), .B1(new_n743), .B2(new_n574), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n580), .A3(new_n647), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n604), .A2(new_n520), .ZN(new_n750));
  XOR2_X1   g564(.A(new_n750), .B(KEYINPUT43), .Z(new_n751));
  NOR2_X1   g565(.A1(new_n617), .A2(new_n620), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT44), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n712), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n752), .A3(KEYINPUT44), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT106), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n749), .B(new_n754), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  INV_X1    g574(.A(KEYINPUT47), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT107), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n747), .A2(new_n580), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n745), .A2(new_n746), .ZN(new_n765));
  OAI211_X1 g579(.A(KEYINPUT107), .B(new_n761), .C1(new_n765), .C2(new_n579), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n638), .A2(new_n228), .A3(new_n665), .A4(new_n712), .ZN(new_n768));
  AND3_X1   g582(.A1(new_n767), .A2(KEYINPUT108), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT108), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n190), .ZN(G42));
  NOR3_X1   g586(.A1(new_n592), .A2(new_n593), .A3(new_n347), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n674), .A2(new_n773), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n774), .A2(new_n656), .A3(new_n229), .A4(new_n522), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n604), .A2(new_n605), .ZN(new_n778));
  INV_X1    g592(.A(new_n639), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n779), .A2(new_n751), .A3(new_n674), .A4(new_n773), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n777), .A2(new_n778), .B1(new_n707), .B2(new_n780), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n228), .A2(new_n751), .A3(new_n779), .A4(new_n699), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n783));
  INV_X1    g597(.A(new_n674), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n783), .B1(new_n784), .B2(new_n346), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n674), .A2(KEYINPUT116), .A3(new_n347), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n782), .A2(new_n646), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n782), .A2(new_n773), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n671), .A2(new_n579), .A3(new_n573), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n764), .A2(new_n766), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n781), .A2(new_n789), .A3(KEYINPUT51), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n777), .A2(new_n605), .A3(new_n604), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n780), .A2(new_n345), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT48), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n455), .A2(G952), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n674), .A2(new_n414), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n798), .B1(new_n782), .B2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n794), .A2(new_n795), .A3(new_n797), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n789), .A2(KEYINPUT117), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n791), .B(KEYINPUT115), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n790), .B1(new_n767), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n789), .A2(KEYINPUT117), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n803), .A2(new_n805), .A3(new_n781), .A4(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n534), .B(KEYINPUT110), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n605), .A2(new_n641), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n582), .A2(new_n773), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n620), .B1(new_n331), .B2(new_n344), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n724), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n723), .B1(new_n722), .B2(new_n580), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n773), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n281), .B1(new_n630), .B2(new_n280), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(new_n694), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n304), .A2(KEYINPUT99), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n309), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n336), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n690), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n709), .A2(new_n621), .A3(new_n824), .A4(new_n587), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  INV_X1    g641(.A(new_n825), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n828), .B2(new_n725), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n815), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n606), .B1(new_n811), .B2(new_n605), .ZN(new_n831));
  INV_X1    g645(.A(new_n594), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n589), .A4(new_n582), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n584), .A2(new_n622), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n830), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n681), .A2(new_n675), .A3(new_n678), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n704), .B2(new_n701), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n728), .A2(new_n729), .B1(new_n734), .B2(new_n736), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n620), .A2(new_n580), .A3(new_n664), .A4(new_n722), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n344), .B2(new_n655), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n687), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n643), .A3(new_n667), .A4(new_n710), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT52), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n810), .B1(new_n839), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n584), .A2(new_n622), .A3(new_n833), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT111), .B1(new_n818), .B2(new_n825), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n828), .A2(new_n725), .A3(new_n827), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(new_n848), .B1(new_n814), .B2(new_n813), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n730), .A2(new_n846), .A3(new_n737), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n687), .B2(new_n841), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n643), .A2(new_n710), .A3(KEYINPUT112), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT112), .B1(new_n643), .B2(new_n710), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n667), .B(new_n852), .C1(new_n853), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n843), .A2(new_n851), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n850), .A2(new_n857), .A3(KEYINPUT53), .A4(new_n837), .ZN(new_n858));
  XNOR2_X1  g672(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n845), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n839), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT53), .B1(new_n861), .B2(new_n857), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n839), .A2(new_n844), .A3(new_n810), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n863), .A2(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(KEYINPUT113), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n809), .B(new_n860), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n868), .B1(G952), .B2(G953), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n228), .A2(new_n580), .A3(new_n346), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n671), .A2(new_n573), .ZN(new_n871));
  AOI211_X1 g685(.A(new_n750), .B(new_n870), .C1(new_n871), .C2(KEYINPUT49), .ZN(new_n872));
  INV_X1    g686(.A(new_n656), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n871), .A2(KEYINPUT49), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n874), .B(KEYINPUT109), .Z(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n646), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(G75));
  AOI21_X1  g691(.A(new_n218), .B1(new_n845), .B2(new_n858), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(G210), .ZN(new_n879));
  NOR2_X1   g693(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT55), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT55), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n879), .A2(new_n883), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n379), .A2(new_n385), .A3(new_n394), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(new_n392), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n887), .B1(new_n882), .B2(new_n884), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n455), .A2(G952), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(G51));
  NAND2_X1  g706(.A1(new_n845), .A2(new_n858), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(new_n859), .Z(new_n894));
  XOR2_X1   g708(.A(new_n574), .B(KEYINPUT57), .Z(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n566), .A3(new_n572), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n743), .B(KEYINPUT120), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n878), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n891), .B1(new_n897), .B2(new_n899), .ZN(G54));
  NAND3_X1  g714(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n901));
  INV_X1    g715(.A(new_n515), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n891), .ZN(G60));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT59), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n894), .A2(new_n599), .A3(new_n597), .A4(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(new_n891), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n907), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n597), .A2(new_n599), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G63));
  NAND2_X1  g728(.A1(G217), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT60), .Z(new_n916));
  NAND2_X1  g730(.A1(new_n893), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT122), .ZN(new_n918));
  INV_X1    g732(.A(new_n217), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n893), .A2(new_n920), .A3(new_n916), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n893), .B2(new_n916), .ZN(new_n923));
  INV_X1    g737(.A(new_n916), .ZN(new_n924));
  AOI211_X1 g738(.A(KEYINPUT122), .B(new_n924), .C1(new_n845), .C2(new_n858), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n619), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n922), .A2(new_n926), .A3(new_n909), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n927), .A2(KEYINPUT121), .A3(KEYINPUT61), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT61), .B1(new_n927), .B2(KEYINPUT121), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  INV_X1    g744(.A(new_n524), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n931), .B2(new_n390), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n837), .A2(new_n846), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n934), .B2(G953), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n886), .B1(G898), .B2(new_n455), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT123), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n935), .B(new_n937), .ZN(G69));
  AOI21_X1  g752(.A(new_n455), .B1(G227), .B2(G900), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n323), .A2(new_n324), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(new_n507), .Z(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n648), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n345), .A2(new_n948), .A3(new_n773), .A4(new_n831), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n759), .B(new_n949), .C1(new_n769), .C2(new_n770), .ZN(new_n950));
  INV_X1    g764(.A(new_n661), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n643), .A2(new_n710), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT112), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n643), .A2(new_n710), .A3(KEYINPUT112), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n957), .B2(new_n667), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n952), .B(new_n667), .C1(new_n853), .C2(new_n854), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n951), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n667), .B1(new_n853), .B2(new_n854), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n959), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(KEYINPUT62), .A3(new_n951), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n950), .B1(new_n963), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n947), .B1(new_n968), .B2(G953), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n749), .A2(new_n345), .A3(new_n687), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n759), .A2(new_n730), .A3(new_n737), .A4(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n771), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n972), .A2(new_n455), .A3(new_n966), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n947), .B1(G900), .B2(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n940), .A2(KEYINPUT126), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n943), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  AOI211_X1 g793(.A(KEYINPUT127), .B(new_n979), .C1(new_n969), .C2(new_n975), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n942), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n950), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT62), .B1(new_n966), .B2(new_n951), .ZN(new_n983));
  AOI211_X1 g797(.A(new_n962), .B(new_n661), .C1(new_n965), .C2(new_n959), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n946), .B1(new_n985), .B2(new_n455), .ZN(new_n986));
  INV_X1    g800(.A(new_n975), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n977), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT127), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n976), .A2(new_n943), .A3(new_n977), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n990), .A3(new_n941), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n981), .A2(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(new_n327), .A2(new_n332), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n651), .B(KEYINPUT63), .Z(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n866), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n326), .A2(new_n309), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n968), .A2(new_n934), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n998), .B2(new_n994), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n972), .A2(new_n934), .A3(new_n966), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n309), .B(new_n326), .C1(new_n1000), .C2(new_n994), .ZN(new_n1001));
  NOR4_X1   g815(.A1(new_n996), .A2(new_n999), .A3(new_n891), .A4(new_n1001), .ZN(G57));
endmodule


