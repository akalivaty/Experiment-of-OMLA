

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(G2104), .A2(G2105), .ZN(n904) );
  INV_X2 U553 ( .A(n747), .ZN(n731) );
  XNOR2_X2 U554 ( .A(KEYINPUT15), .B(n587), .ZN(n1003) );
  AND2_X2 U555 ( .A1(n530), .A2(G2104), .ZN(n908) );
  XNOR2_X1 U556 ( .A(n746), .B(n745), .ZN(n762) );
  NOR2_X1 U557 ( .A1(n690), .A2(n689), .ZN(n692) );
  AND2_X1 U558 ( .A1(n813), .A2(n812), .ZN(n517) );
  AND2_X1 U559 ( .A1(n810), .A2(n839), .ZN(n518) );
  AND2_X1 U560 ( .A1(n731), .A2(G1996), .ZN(n705) );
  INV_X1 U561 ( .A(KEYINPUT31), .ZN(n744) );
  NOR2_X1 U562 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U563 ( .A(n744), .B(KEYINPUT106), .ZN(n745) );
  INV_X1 U564 ( .A(KEYINPUT100), .ZN(n736) );
  XNOR2_X1 U565 ( .A(n759), .B(KEYINPUT32), .ZN(n768) );
  OR2_X1 U566 ( .A1(G1384), .A2(n695), .ZN(n696) );
  XOR2_X1 U567 ( .A(G2443), .B(G2446), .Z(n520) );
  XNOR2_X1 U568 ( .A(G2427), .B(G2451), .ZN(n519) );
  XNOR2_X1 U569 ( .A(n520), .B(n519), .ZN(n526) );
  XOR2_X1 U570 ( .A(G2430), .B(G2454), .Z(n522) );
  XNOR2_X1 U571 ( .A(G1341), .B(G1348), .ZN(n521) );
  XNOR2_X1 U572 ( .A(n522), .B(n521), .ZN(n524) );
  XOR2_X1 U573 ( .A(G2435), .B(G2438), .Z(n523) );
  XNOR2_X1 U574 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U575 ( .A(n526), .B(n525), .Z(n527) );
  AND2_X1 U576 ( .A1(G14), .A2(n527), .ZN(G401) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n528) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n528), .Z(n907) );
  NAND2_X1 U579 ( .A1(n907), .A2(G138), .ZN(n535) );
  INV_X1 U580 ( .A(G2105), .ZN(n530) );
  NOR2_X1 U581 ( .A1(G2104), .A2(n530), .ZN(n607) );
  NAND2_X1 U582 ( .A1(G126), .A2(n607), .ZN(n529) );
  XNOR2_X1 U583 ( .A(KEYINPUT91), .B(n529), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G102), .A2(n908), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G114), .A2(n904), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n695) );
  AND2_X1 U588 ( .A1(n535), .A2(n695), .ZN(G164) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G57), .ZN(G237) );
  INV_X1 U591 ( .A(G82), .ZN(G220) );
  NAND2_X1 U592 ( .A1(n907), .A2(G137), .ZN(n691) );
  NAND2_X1 U593 ( .A1(G101), .A2(n908), .ZN(n536) );
  XNOR2_X1 U594 ( .A(KEYINPUT23), .B(n536), .ZN(n689) );
  NAND2_X1 U595 ( .A1(G125), .A2(n607), .ZN(n538) );
  NAND2_X1 U596 ( .A1(G113), .A2(n904), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n687) );
  NOR2_X1 U598 ( .A1(n689), .A2(n687), .ZN(n539) );
  AND2_X1 U599 ( .A1(n691), .A2(n539), .ZN(G160) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n648) );
  NAND2_X1 U601 ( .A1(n648), .A2(G89), .ZN(n540) );
  XNOR2_X1 U602 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  XOR2_X1 U603 ( .A(G543), .B(KEYINPUT0), .Z(n637) );
  INV_X1 U604 ( .A(G651), .ZN(n545) );
  NOR2_X1 U605 ( .A1(n637), .A2(n545), .ZN(n656) );
  NAND2_X1 U606 ( .A1(G76), .A2(n656), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(KEYINPUT5), .B(n543), .ZN(n554) );
  NOR2_X1 U609 ( .A1(G651), .A2(n637), .ZN(n544) );
  XOR2_X1 U610 ( .A(KEYINPUT65), .B(n544), .Z(n652) );
  NAND2_X1 U611 ( .A1(G51), .A2(n652), .ZN(n549) );
  NOR2_X1 U612 ( .A1(G543), .A2(n545), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT1), .B(n546), .Z(n581) );
  BUF_X1 U614 ( .A(n581), .Z(n647) );
  NAND2_X1 U615 ( .A1(n647), .A2(G63), .ZN(n547) );
  XOR2_X1 U616 ( .A(KEYINPUT77), .B(n547), .Z(n548) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n550), .B(KEYINPUT6), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT7), .B(n555), .ZN(G168) );
  XOR2_X1 U623 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U624 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT72), .B(KEYINPUT10), .Z(n557) );
  NAND2_X1 U626 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U627 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U628 ( .A(KEYINPUT71), .B(n558), .Z(n844) );
  NAND2_X1 U629 ( .A1(n844), .A2(G567), .ZN(n559) );
  XNOR2_X1 U630 ( .A(n560), .B(n559), .ZN(n561) );
  XOR2_X1 U631 ( .A(KEYINPUT73), .B(n561), .Z(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n647), .ZN(n562) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n562), .Z(n568) );
  NAND2_X1 U634 ( .A1(n648), .A2(G81), .ZN(n563) );
  XNOR2_X1 U635 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U636 ( .A1(G68), .A2(n656), .ZN(n564) );
  NAND2_X1 U637 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NOR2_X1 U639 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U640 ( .A1(n652), .A2(G43), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n1006) );
  XNOR2_X1 U642 ( .A(G860), .B(KEYINPUT75), .ZN(n601) );
  OR2_X1 U643 ( .A1(n1006), .A2(n601), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G52), .A2(n652), .ZN(n571) );
  XNOR2_X1 U645 ( .A(n571), .B(KEYINPUT67), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G90), .A2(n648), .ZN(n573) );
  NAND2_X1 U647 ( .A1(G77), .A2(n656), .ZN(n572) );
  NAND2_X1 U648 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U649 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  NOR2_X1 U650 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n647), .A2(G64), .ZN(n577) );
  NAND2_X1 U652 ( .A1(n578), .A2(n577), .ZN(G301) );
  NAND2_X1 U653 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n652), .A2(G54), .ZN(n586) );
  NAND2_X1 U655 ( .A1(G92), .A2(n648), .ZN(n580) );
  NAND2_X1 U656 ( .A1(G79), .A2(n656), .ZN(n579) );
  NAND2_X1 U657 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n581), .A2(G66), .ZN(n582) );
  XOR2_X1 U659 ( .A(KEYINPUT76), .B(n582), .Z(n583) );
  NOR2_X1 U660 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U662 ( .A(n1003), .ZN(n714) );
  INV_X1 U663 ( .A(G868), .ZN(n671) );
  NAND2_X1 U664 ( .A1(n714), .A2(n671), .ZN(n588) );
  NAND2_X1 U665 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U666 ( .A1(G91), .A2(n648), .ZN(n590) );
  XOR2_X1 U667 ( .A(KEYINPUT68), .B(n590), .Z(n595) );
  NAND2_X1 U668 ( .A1(G65), .A2(n647), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G53), .A2(n652), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U671 ( .A(KEYINPUT69), .B(n593), .Z(n594) );
  NOR2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n656), .A2(G78), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U675 ( .A1(G868), .A2(G299), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT80), .ZN(n600) );
  NOR2_X1 U677 ( .A1(n671), .A2(G286), .ZN(n599) );
  NOR2_X1 U678 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U679 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U680 ( .A1(n602), .A2(n1003), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U682 ( .A1(G868), .A2(n1006), .ZN(n606) );
  NAND2_X1 U683 ( .A1(G868), .A2(n1003), .ZN(n604) );
  NOR2_X1 U684 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U685 ( .A1(n606), .A2(n605), .ZN(G282) );
  XNOR2_X1 U686 ( .A(G2100), .B(KEYINPUT81), .ZN(n616) );
  BUF_X1 U687 ( .A(n607), .Z(n903) );
  NAND2_X1 U688 ( .A1(n903), .A2(G123), .ZN(n608) );
  XNOR2_X1 U689 ( .A(n608), .B(KEYINPUT18), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G111), .A2(n904), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U692 ( .A1(G135), .A2(n907), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G99), .A2(n908), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n934) );
  XNOR2_X1 U696 ( .A(n934), .B(G2096), .ZN(n615) );
  NAND2_X1 U697 ( .A1(n616), .A2(n615), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G80), .A2(n656), .ZN(n617) );
  XNOR2_X1 U699 ( .A(n617), .B(KEYINPUT82), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G67), .A2(n647), .ZN(n619) );
  NAND2_X1 U701 ( .A1(G93), .A2(n648), .ZN(n618) );
  NAND2_X1 U702 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G55), .A2(n652), .ZN(n620) );
  XNOR2_X1 U704 ( .A(KEYINPUT83), .B(n620), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n670) );
  NAND2_X1 U707 ( .A1(G559), .A2(n1003), .ZN(n625) );
  XNOR2_X1 U708 ( .A(n1006), .B(n625), .ZN(n668) );
  NOR2_X1 U709 ( .A1(G860), .A2(n668), .ZN(n626) );
  XOR2_X1 U710 ( .A(n670), .B(n626), .Z(G145) );
  NAND2_X1 U711 ( .A1(n652), .A2(G47), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n647), .A2(G60), .ZN(n627) );
  NAND2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U714 ( .A(KEYINPUT66), .B(n629), .Z(n633) );
  NAND2_X1 U715 ( .A1(G85), .A2(n648), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G72), .A2(n656), .ZN(n630) );
  AND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U719 ( .A1(G49), .A2(n652), .ZN(n635) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n634) );
  NAND2_X1 U721 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U722 ( .A1(n647), .A2(n636), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U724 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U725 ( .A1(G62), .A2(n647), .ZN(n641) );
  NAND2_X1 U726 ( .A1(G75), .A2(n656), .ZN(n640) );
  NAND2_X1 U727 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U728 ( .A1(n648), .A2(G88), .ZN(n642) );
  XOR2_X1 U729 ( .A(KEYINPUT88), .B(n642), .Z(n643) );
  NOR2_X1 U730 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n652), .A2(G50), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(G303) );
  NAND2_X1 U733 ( .A1(G61), .A2(n647), .ZN(n650) );
  NAND2_X1 U734 ( .A1(G86), .A2(n648), .ZN(n649) );
  NAND2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U736 ( .A(KEYINPUT84), .B(n651), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n652), .A2(G48), .ZN(n653) );
  XOR2_X1 U738 ( .A(KEYINPUT86), .B(n653), .Z(n654) );
  NOR2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n660) );
  XOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT2), .Z(n658) );
  NAND2_X1 U741 ( .A1(G73), .A2(n656), .ZN(n657) );
  XNOR2_X1 U742 ( .A(n658), .B(n657), .ZN(n659) );
  NAND2_X1 U743 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U744 ( .A(KEYINPUT87), .B(n661), .Z(G305) );
  XNOR2_X1 U745 ( .A(KEYINPUT89), .B(G290), .ZN(n662) );
  XNOR2_X1 U746 ( .A(n662), .B(G288), .ZN(n665) );
  XOR2_X1 U747 ( .A(G303), .B(G305), .Z(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(n670), .ZN(n664) );
  XNOR2_X1 U749 ( .A(n665), .B(n664), .ZN(n667) );
  XNOR2_X1 U750 ( .A(G299), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n667), .B(n666), .ZN(n851) );
  XOR2_X1 U752 ( .A(n668), .B(n851), .Z(n669) );
  NAND2_X1 U753 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2084), .A2(G2078), .ZN(n674) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n674), .Z(n675) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n675), .ZN(n676) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n676), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U762 ( .A(KEYINPUT70), .B(G132), .Z(G219) );
  NOR2_X1 U763 ( .A1(G219), .A2(G220), .ZN(n678) );
  XOR2_X1 U764 ( .A(KEYINPUT22), .B(n678), .Z(n679) );
  XNOR2_X1 U765 ( .A(n679), .B(KEYINPUT90), .ZN(n680) );
  NOR2_X1 U766 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G96), .A2(n681), .ZN(n849) );
  NAND2_X1 U768 ( .A1(n849), .A2(G2106), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G120), .A2(G108), .ZN(n682) );
  NOR2_X1 U770 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U771 ( .A1(G69), .A2(n683), .ZN(n850) );
  NAND2_X1 U772 ( .A1(n850), .A2(G567), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n925) );
  NAND2_X1 U774 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n925), .A2(n686), .ZN(n848) );
  NAND2_X1 U776 ( .A1(n848), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G303), .ZN(G166) );
  INV_X1 U778 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U779 ( .A(KEYINPUT112), .B(KEYINPUT40), .ZN(n843) );
  XOR2_X1 U780 ( .A(G1981), .B(G305), .Z(n1021) );
  INV_X1 U781 ( .A(n687), .ZN(n688) );
  NAND2_X1 U782 ( .A1(G40), .A2(n688), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n791) );
  INV_X1 U784 ( .A(n791), .ZN(n698) );
  INV_X1 U785 ( .A(G1384), .ZN(n693) );
  AND2_X1 U786 ( .A1(G138), .A2(n693), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n907), .A2(n694), .ZN(n697) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n790) );
  NAND2_X2 U789 ( .A1(n698), .A2(n790), .ZN(n747) );
  NAND2_X1 U790 ( .A1(G8), .A2(n747), .ZN(n787) );
  NOR2_X1 U791 ( .A1(G288), .A2(G1976), .ZN(n699) );
  XOR2_X1 U792 ( .A(n699), .B(KEYINPUT107), .Z(n770) );
  INV_X1 U793 ( .A(n770), .ZN(n700) );
  NOR2_X1 U794 ( .A1(n787), .A2(n700), .ZN(n701) );
  NAND2_X1 U795 ( .A1(KEYINPUT33), .A2(n701), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n1021), .A2(n702), .ZN(n776) );
  XOR2_X1 U797 ( .A(KEYINPUT26), .B(KEYINPUT102), .Z(n703) );
  XNOR2_X1 U798 ( .A(KEYINPUT64), .B(n703), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n747), .A2(G1341), .ZN(n706) );
  NAND2_X1 U801 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X2 U802 ( .A1(n1006), .A2(n708), .ZN(n715) );
  NOR2_X2 U803 ( .A1(n715), .A2(n714), .ZN(n709) );
  XNOR2_X1 U804 ( .A(n709), .B(KEYINPUT103), .ZN(n713) );
  NOR2_X1 U805 ( .A1(n731), .A2(G1348), .ZN(n711) );
  NOR2_X1 U806 ( .A1(G2067), .A2(n747), .ZN(n710) );
  NOR2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U811 ( .A(KEYINPUT104), .B(n718), .Z(n724) );
  NAND2_X1 U812 ( .A1(n731), .A2(G2072), .ZN(n719) );
  XOR2_X1 U813 ( .A(KEYINPUT27), .B(n719), .Z(n721) );
  NAND2_X1 U814 ( .A1(G1956), .A2(n747), .ZN(n720) );
  NAND2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G299), .A2(n725), .ZN(n722) );
  XOR2_X1 U817 ( .A(KEYINPUT105), .B(n722), .Z(n723) );
  NOR2_X1 U818 ( .A1(n724), .A2(n723), .ZN(n728) );
  NAND2_X1 U819 ( .A1(G299), .A2(n725), .ZN(n726) );
  XOR2_X1 U820 ( .A(KEYINPUT28), .B(n726), .Z(n727) );
  XNOR2_X1 U821 ( .A(n729), .B(KEYINPUT29), .ZN(n735) );
  INV_X1 U822 ( .A(G1961), .ZN(n867) );
  NAND2_X1 U823 ( .A1(n747), .A2(n867), .ZN(n733) );
  XOR2_X1 U824 ( .A(G2078), .B(KEYINPUT25), .Z(n730) );
  XNOR2_X1 U825 ( .A(KEYINPUT101), .B(n730), .ZN(n951) );
  NAND2_X1 U826 ( .A1(n731), .A2(n951), .ZN(n732) );
  NAND2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n741) );
  NAND2_X1 U828 ( .A1(G171), .A2(n741), .ZN(n734) );
  NAND2_X1 U829 ( .A1(n735), .A2(n734), .ZN(n761) );
  NOR2_X1 U830 ( .A1(G2084), .A2(n747), .ZN(n760) );
  NOR2_X1 U831 ( .A1(G1966), .A2(n787), .ZN(n737) );
  XNOR2_X1 U832 ( .A(n737), .B(n736), .ZN(n763) );
  NAND2_X1 U833 ( .A1(n763), .A2(G8), .ZN(n738) );
  NOR2_X1 U834 ( .A1(n760), .A2(n738), .ZN(n739) );
  XOR2_X1 U835 ( .A(KEYINPUT30), .B(n739), .Z(n740) );
  NOR2_X1 U836 ( .A1(G168), .A2(n740), .ZN(n743) );
  NOR2_X1 U837 ( .A1(G171), .A2(n741), .ZN(n742) );
  NOR2_X1 U838 ( .A1(n743), .A2(n742), .ZN(n746) );
  INV_X1 U839 ( .A(G8), .ZN(n752) );
  NOR2_X1 U840 ( .A1(G1971), .A2(n787), .ZN(n749) );
  NOR2_X1 U841 ( .A1(G2090), .A2(n747), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n750), .A2(G303), .ZN(n751) );
  OR2_X1 U844 ( .A1(n752), .A2(n751), .ZN(n754) );
  AND2_X1 U845 ( .A1(n762), .A2(n754), .ZN(n753) );
  NAND2_X1 U846 ( .A1(n761), .A2(n753), .ZN(n758) );
  INV_X1 U847 ( .A(n754), .ZN(n756) );
  AND2_X1 U848 ( .A1(G286), .A2(G8), .ZN(n755) );
  OR2_X1 U849 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U851 ( .A1(G8), .A2(n760), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n762), .A2(n761), .ZN(n764) );
  AND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n784) );
  NOR2_X1 U856 ( .A1(G1971), .A2(G303), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n1012) );
  NAND2_X1 U858 ( .A1(n784), .A2(n1012), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n1011) );
  NAND2_X1 U860 ( .A1(n771), .A2(n1011), .ZN(n772) );
  XNOR2_X1 U861 ( .A(n772), .B(KEYINPUT108), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n773), .A2(n787), .ZN(n774) );
  NOR2_X1 U863 ( .A1(KEYINPUT33), .A2(n774), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n781) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n777) );
  XNOR2_X1 U866 ( .A(n777), .B(KEYINPUT99), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT24), .ZN(n779) );
  NOR2_X1 U868 ( .A1(n779), .A2(n787), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n789) );
  NAND2_X1 U870 ( .A1(G8), .A2(G166), .ZN(n782) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n782), .ZN(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT109), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U874 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n813) );
  XNOR2_X1 U876 ( .A(G1986), .B(G290), .ZN(n1008) );
  NOR2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n839) );
  NAND2_X1 U878 ( .A1(n1008), .A2(n839), .ZN(n792) );
  XOR2_X1 U879 ( .A(KEYINPUT92), .B(n792), .Z(n811) );
  NAND2_X1 U880 ( .A1(G129), .A2(n903), .ZN(n794) );
  NAND2_X1 U881 ( .A1(G141), .A2(n907), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n794), .A2(n793), .ZN(n797) );
  NAND2_X1 U883 ( .A1(n908), .A2(G105), .ZN(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT38), .B(n795), .Z(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n904), .A2(G117), .ZN(n798) );
  NAND2_X1 U887 ( .A1(n799), .A2(n798), .ZN(n896) );
  NAND2_X1 U888 ( .A1(G1996), .A2(n896), .ZN(n800) );
  XOR2_X1 U889 ( .A(KEYINPUT98), .B(n800), .Z(n809) );
  NAND2_X1 U890 ( .A1(G119), .A2(n903), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G107), .A2(n904), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n807) );
  NAND2_X1 U893 ( .A1(G131), .A2(n907), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G95), .A2(n908), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT97), .B(n805), .Z(n806) );
  OR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n914) );
  AND2_X1 U898 ( .A1(n914), .A2(G1991), .ZN(n808) );
  NOR2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n936) );
  INV_X1 U900 ( .A(n936), .ZN(n810) );
  NOR2_X1 U901 ( .A1(n811), .A2(n518), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G140), .A2(n907), .ZN(n815) );
  NAND2_X1 U903 ( .A1(G104), .A2(n908), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U905 ( .A(KEYINPUT34), .B(n816), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G128), .A2(n903), .ZN(n818) );
  NAND2_X1 U907 ( .A1(G116), .A2(n904), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U909 ( .A(KEYINPUT93), .B(n819), .ZN(n820) );
  XNOR2_X1 U910 ( .A(KEYINPUT35), .B(n820), .ZN(n821) );
  NOR2_X1 U911 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U912 ( .A(n823), .B(KEYINPUT36), .ZN(n824) );
  XOR2_X1 U913 ( .A(n824), .B(KEYINPUT94), .Z(n893) );
  XOR2_X1 U914 ( .A(G2067), .B(KEYINPUT37), .Z(n835) );
  NAND2_X1 U915 ( .A1(n893), .A2(n835), .ZN(n825) );
  XNOR2_X1 U916 ( .A(n825), .B(KEYINPUT95), .ZN(n946) );
  NAND2_X1 U917 ( .A1(n946), .A2(n839), .ZN(n826) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT96), .ZN(n833) );
  NAND2_X1 U919 ( .A1(n517), .A2(n833), .ZN(n841) );
  NOR2_X1 U920 ( .A1(G1996), .A2(n896), .ZN(n929) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U922 ( .A1(n914), .A2(G1991), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n827), .B(KEYINPUT110), .ZN(n926) );
  NOR2_X1 U924 ( .A1(n828), .A2(n926), .ZN(n829) );
  NOR2_X1 U925 ( .A1(n518), .A2(n829), .ZN(n830) );
  XOR2_X1 U926 ( .A(KEYINPUT111), .B(n830), .Z(n831) );
  NOR2_X1 U927 ( .A1(n929), .A2(n831), .ZN(n832) );
  XNOR2_X1 U928 ( .A(KEYINPUT39), .B(n832), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n834), .A2(n833), .ZN(n837) );
  NOR2_X1 U930 ( .A1(n893), .A2(n835), .ZN(n927) );
  INV_X1 U931 ( .A(n927), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U933 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U934 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U935 ( .A(n843), .B(n842), .ZN(G329) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n844), .ZN(G217) );
  INV_X1 U937 ( .A(n844), .ZN(G223) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G661), .A2(n845), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n846) );
  XOR2_X1 U941 ( .A(KEYINPUT113), .B(n846), .Z(n847) );
  NAND2_X1 U942 ( .A1(n848), .A2(n847), .ZN(G188) );
  XNOR2_X1 U943 ( .A(G108), .B(KEYINPUT121), .ZN(G238) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U948 ( .A(n1006), .B(n851), .ZN(n853) );
  XOR2_X1 U949 ( .A(G301), .B(n1003), .Z(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U951 ( .A(G286), .B(n854), .ZN(n855) );
  NOR2_X1 U952 ( .A1(G37), .A2(n855), .ZN(G397) );
  XOR2_X1 U953 ( .A(G2678), .B(KEYINPUT115), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT114), .B(G2100), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n858), .B(KEYINPUT42), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(G2096), .B(G2090), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2084), .B(G2078), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U963 ( .A(KEYINPUT43), .B(KEYINPUT116), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G227) );
  INV_X1 U965 ( .A(G1971), .ZN(n1013) );
  XNOR2_X1 U966 ( .A(G1976), .B(n1013), .ZN(n869) );
  XOR2_X1 U967 ( .A(G1986), .B(n867), .Z(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(n870), .B(G2474), .Z(n872) );
  XNOR2_X1 U970 ( .A(G1966), .B(G1981), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT41), .B(G1956), .Z(n874) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1991), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U976 ( .A1(G124), .A2(n903), .ZN(n877) );
  XOR2_X1 U977 ( .A(KEYINPUT117), .B(n877), .Z(n878) );
  XNOR2_X1 U978 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G112), .A2(n904), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G136), .A2(n907), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G100), .A2(n908), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U984 ( .A1(n884), .A2(n883), .ZN(G162) );
  NAND2_X1 U985 ( .A1(G139), .A2(n907), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G103), .A2(n908), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n891) );
  NAND2_X1 U988 ( .A1(G127), .A2(n903), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G115), .A2(n904), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(KEYINPUT118), .B(n892), .Z(n937) );
  XOR2_X1 U994 ( .A(G162), .B(n937), .Z(n895) );
  XOR2_X1 U995 ( .A(G160), .B(n893), .Z(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n900) );
  XNOR2_X1 U997 ( .A(KEYINPUT119), .B(KEYINPUT48), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n896), .B(KEYINPUT46), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U1001 ( .A(G164), .B(n934), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n917) );
  NAND2_X1 U1003 ( .A1(G130), .A2(n903), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(G118), .A2(n904), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n913) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n907), .ZN(n910) );
  NAND2_X1 U1007 ( .A1(G106), .A2(n908), .ZN(n909) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(n911), .B(KEYINPUT45), .Z(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n915), .B(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n918), .ZN(G395) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n919), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n920), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(n925), .A2(G401), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT120), .B(n921), .Z(n922) );
  NOR2_X1 U1019 ( .A1(G395), .A2(n922), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n925), .ZN(G319) );
  INV_X1 U1023 ( .A(G96), .ZN(G221) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(KEYINPUT55), .ZN(n949) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n944) );
  XNOR2_X1 U1027 ( .A(G160), .B(G2084), .ZN(n932) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n930), .Z(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n939) );
  XNOR2_X1 U1035 ( .A(G2072), .B(n937), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n950), .A2(G29), .ZN(n1002) );
  XNOR2_X1 U1044 ( .A(G27), .B(n951), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G2072), .B(G33), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1049 ( .A(G32), .B(G1996), .ZN(n956) );
  NOR2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1051 ( .A(KEYINPUT122), .B(n958), .Z(n960) );
  XNOR2_X1 U1052 ( .A(G1991), .B(G25), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(G28), .A2(n961), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n994) );
  NAND2_X1 U1061 ( .A1(KEYINPUT55), .A2(n994), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n968), .ZN(n1000) );
  XOR2_X1 U1063 ( .A(G1986), .B(G24), .Z(n971) );
  XNOR2_X1 U1064 ( .A(G22), .B(KEYINPUT127), .ZN(n969) );
  XOR2_X1 U1065 ( .A(n969), .B(n1013), .Z(n970) );
  NAND2_X1 U1066 ( .A1(n971), .A2(n970), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(G23), .B(G1976), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1069 ( .A(KEYINPUT58), .B(n974), .Z(n991) );
  XOR2_X1 U1070 ( .A(G1966), .B(G21), .Z(n976) );
  XOR2_X1 U1071 ( .A(G1961), .B(G5), .Z(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n988) );
  XNOR2_X1 U1073 ( .A(G1348), .B(KEYINPUT59), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n977), .B(G4), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(G1956), .B(G20), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(G6), .B(G1981), .ZN(n978) );
  NOR2_X1 U1077 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT124), .B(G1341), .ZN(n982) );
  XNOR2_X1 U1080 ( .A(G19), .B(n982), .ZN(n983) );
  NOR2_X1 U1081 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1082 ( .A(KEYINPUT60), .B(n985), .ZN(n986) );
  XNOR2_X1 U1083 ( .A(KEYINPUT125), .B(n986), .ZN(n987) );
  NOR2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1085 ( .A(KEYINPUT126), .B(n989), .Z(n990) );
  NOR2_X1 U1086 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1087 ( .A(n992), .B(KEYINPUT61), .ZN(n993) );
  INV_X1 U1088 ( .A(G16), .ZN(n1026) );
  NAND2_X1 U1089 ( .A1(n993), .A2(n1026), .ZN(n998) );
  INV_X1 U1090 ( .A(n994), .ZN(n996) );
  NOR2_X1 U1091 ( .A1(G29), .A2(KEYINPUT55), .ZN(n995) );
  NAND2_X1 U1092 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1093 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1094 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1030) );
  XNOR2_X1 U1096 ( .A(G299), .B(G1956), .ZN(n1005) );
  XOR2_X1 U1097 ( .A(n1003), .B(G1348), .Z(n1004) );
  NOR2_X1 U1098 ( .A1(n1005), .A2(n1004), .ZN(n1020) );
  XOR2_X1 U1099 ( .A(G301), .B(G1961), .Z(n1010) );
  XNOR2_X1 U1100 ( .A(G1341), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1101 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  NOR2_X1 U1104 ( .A1(G166), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(n1016), .B(KEYINPUT123), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1108 ( .A1(n1020), .A2(n1019), .ZN(n1025) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G168), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(KEYINPUT57), .B(n1023), .Z(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(KEYINPUT56), .B(n1026), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(n1031), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1117 ( .A(G150), .ZN(G311) );
endmodule

