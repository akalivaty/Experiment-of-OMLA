//key=1010101010101010101010101010101010101010101010101010101010101010

module locked_c3540 ( G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, 
        G97, G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, 
        G179, G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, 
        G264, G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, 
        G343, G1698, G2897, G353, G355, G361, G358, G351, G372, G369, G399, 
        G364, G396, G384, G367, G387, G393, G390, G378, G375, G381, G407, G409, 
        G405, G402, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, 
        KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, 
        KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, 
        KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, 
        KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, 
        KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, 
        KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, 
        KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, 
        KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, 
        KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, 
        KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0 );
  input G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97, G107, G116,
         G124, G125, G128, G132, G137, G143, G150, G159, G169, G179, G190,
         G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
         G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330,
         G343, G1698, G2897, KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60,
         KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55,
         KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50,
         KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45,
         KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40,
         KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35,
         KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30,
         KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25,
         KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20,
         KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15,
         KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9,
         KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3,
         KEYINPUT2, KEYINPUT1, KEYINPUT0;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
         G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire   n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1815, n1816, n1817, n1818, n1819, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905;

  NOR2_X1 U976 ( .A1(n972), .A2(n971), .ZN(n976) );
  INV_X1 U977 ( .A(n1345), .ZN(n1402) );
  INV_X2 U978 ( .A(G20), .ZN(n1827) );
  NAND2_X1 U979 ( .A1(n976), .A2(n975), .ZN(n1122) );
  NOR2_X1 U980 ( .A1(n1122), .A2(G179), .ZN(n993) );
  OR2_X1 U981 ( .A1(G1698), .A2(n986), .ZN(n958) );
  NOR2_X2 U982 ( .A1(n1620), .A2(n1449), .ZN(n1467) );
  AND2_X2 U983 ( .A1(n1448), .A2(n1447), .ZN(n1449) );
  INV_X1 U984 ( .A(n958), .ZN(n959) );
  INV_X2 U985 ( .A(n958), .ZN(n960) );
  NOR2_X2 U986 ( .A1(n1402), .A2(n1015), .ZN(n1305) );
  XNOR2_X2 U987 ( .A(n989), .B(n1092), .ZN(n1015) );
  NOR2_X1 U988 ( .A1(n1826), .A2(G33), .ZN(n968) );
  NAND2_X1 U989 ( .A1(n1006), .A2(G294), .ZN(n967) );
  AND2_X1 U990 ( .A1(n966), .A2(G33), .ZN(n1006) );
  NAND2_X1 U991 ( .A1(G1), .A2(G13), .ZN(n964) );
  AND2_X1 U992 ( .A1(G1), .A2(G20), .ZN(n1850) );
  XNOR2_X2 U993 ( .A(G375), .B(G378), .ZN(n1904) );
  NAND2_X2 U994 ( .A1(n1512), .A2(n1511), .ZN(G375) );
  NOR2_X1 U995 ( .A1(n1340), .A2(n1339), .ZN(n1341) );
  XNOR2_X1 U996 ( .A(n1821), .B(G381), .ZN(n1824) );
  XNOR2_X1 U997 ( .A(G390), .B(G396), .ZN(n1821) );
  XNOR2_X1 U998 ( .A(n1334), .B(n1333), .ZN(n1560) );
  NOR2_X1 U999 ( .A1(n1025), .A2(n1024), .ZN(n1067) );
  NOR2_X1 U1000 ( .A1(n1427), .A2(n1426), .ZN(n1428) );
  OR2_X1 U1001 ( .A1(G375), .A2(G378), .ZN(n1811) );
  XNOR2_X1 U1002 ( .A(n1534), .B(KEYINPUT40), .ZN(n1384) );
  XOR2_X1 U1003 ( .A(KEYINPUT1), .B(n1192), .Z(n1672) );
  AND2_X1 U1004 ( .A1(n1114), .A2(n1113), .ZN(n1853) );
  AND2_X1 U1005 ( .A1(n963), .A2(n1112), .ZN(n1113) );
  INV_X1 U1006 ( .A(n1144), .ZN(n1112) );
  XNOR2_X1 U1007 ( .A(n1746), .B(KEYINPUT55), .ZN(G387) );
  NOR2_X1 U1008 ( .A1(n1745), .A2(n1744), .ZN(n1746) );
  XOR2_X1 U1009 ( .A(n1562), .B(n1561), .Z(n961) );
  NOR2_X2 U1010 ( .A1(n1366), .A2(n1163), .ZN(n1775) );
  NOR2_X2 U1011 ( .A1(G200), .A2(n1154), .ZN(n1778) );
  NOR2_X2 U1012 ( .A1(G200), .A2(n1163), .ZN(n1783) );
  NOR2_X2 U1013 ( .A1(n1066), .A2(n1000), .ZN(n1001) );
  NAND2_X1 U1014 ( .A1(n1563), .A2(n1557), .ZN(n1387) );
  NAND2_X1 U1015 ( .A1(n1826), .A2(n980), .ZN(n1279) );
  XOR2_X1 U1016 ( .A(KEYINPUT8), .B(n1087), .Z(n962) );
  AND2_X1 U1017 ( .A1(n1106), .A2(n1682), .ZN(n963) );
  NOR2_X1 U1018 ( .A1(n974), .A2(n1269), .ZN(n1046) );
  BUF_X1 U1019 ( .A(n1006), .Z(n1389) );
  INV_X1 U1020 ( .A(n1115), .ZN(n1125) );
  OR2_X1 U1021 ( .A1(n1431), .A2(n1870), .ZN(n1445) );
  NOR2_X1 U1022 ( .A1(n1374), .A2(n1372), .ZN(n1373) );
  NOR2_X1 U1023 ( .A1(n1365), .A2(n1364), .ZN(n1371) );
  INV_X1 U1024 ( .A(KEYINPUT41), .ZN(n1386) );
  INV_X1 U1025 ( .A(n1598), .ZN(n1333) );
  NAND2_X1 U1026 ( .A1(n1133), .A2(n1132), .ZN(n1430) );
  XNOR2_X1 U1027 ( .A(n1560), .B(KEYINPUT46), .ZN(n1562) );
  NAND2_X1 U1028 ( .A1(n1689), .A2(n1686), .ZN(n1106) );
  INV_X1 U1029 ( .A(G13), .ZN(n1866) );
  XNOR2_X1 U1030 ( .A(G384), .B(G393), .ZN(n1822) );
  XNOR2_X1 U1031 ( .A(G387), .B(n1822), .ZN(n1823) );
  NOR2_X1 U1032 ( .A1(n1828), .A2(G41), .ZN(n1863) );
  XNOR2_X1 U1033 ( .A(n1824), .B(n1823), .ZN(n1905) );
  NAND2_X1 U1034 ( .A1(n1866), .A2(n1850), .ZN(n1828) );
  XNOR2_X2 U1035 ( .A(n964), .B(KEYINPUT2), .ZN(n1826) );
  INV_X1 U1036 ( .A(n968), .ZN(n986) );
  NAND2_X1 U1037 ( .A1(n959), .A2(G250), .ZN(n965) );
  INV_X1 U1038 ( .A(G45), .ZN(n1650) );
  NOR2_X1 U1039 ( .A1(n1650), .A2(G1), .ZN(n1078) );
  INV_X1 U1040 ( .A(n1078), .ZN(n1081) );
  NOR2_X1 U1041 ( .A1(G41), .A2(n1081), .ZN(n974) );
  NAND2_X1 U1042 ( .A1(G274), .A2(n974), .ZN(n1042) );
  NAND2_X1 U1043 ( .A1(n965), .A2(n1042), .ZN(n972) );
  NOR2_X1 U1044 ( .A1(n1826), .A2(G41), .ZN(n966) );
  XNOR2_X1 U1045 ( .A(n967), .B(KEYINPUT14), .ZN(n970) );
  AND2_X2 U1046 ( .A1(n968), .A2(G1698), .ZN(n1393) );
  NAND2_X1 U1047 ( .A1(G257), .A2(n1393), .ZN(n969) );
  NAND2_X1 U1048 ( .A1(n970), .A2(n969), .ZN(n971) );
  AND2_X1 U1049 ( .A1(G41), .A2(G33), .ZN(n973) );
  NOR2_X1 U1050 ( .A1(n1826), .A2(n973), .ZN(n1269) );
  NAND2_X1 U1051 ( .A1(n1046), .A2(G264), .ZN(n975) );
  INV_X1 U1052 ( .A(G169), .ZN(n1400) );
  AND2_X1 U1053 ( .A1(n1122), .A2(n1400), .ZN(n992) );
  NOR2_X1 U1054 ( .A1(n1826), .A2(G20), .ZN(n977) );
  AND2_X2 U1055 ( .A1(G33), .A2(n977), .ZN(n1401) );
  NAND2_X1 U1056 ( .A1(G116), .A2(n1401), .ZN(n978) );
  XNOR2_X1 U1057 ( .A(n978), .B(KEYINPUT16), .ZN(n984) );
  NAND2_X1 U1058 ( .A1(n1850), .A2(G33), .ZN(n979) );
  XOR2_X1 U1059 ( .A(n979), .B(KEYINPUT3), .Z(n980) );
  NOR2_X1 U1060 ( .A1(G1), .A2(n1827), .ZN(n1278) );
  NAND2_X1 U1061 ( .A1(G13), .A2(n1278), .ZN(n1345) );
  NOR2_X1 U1062 ( .A1(n1279), .A2(n1402), .ZN(n982) );
  INV_X1 U1063 ( .A(G33), .ZN(n1498) );
  OR2_X1 U1064 ( .A1(G1), .A2(n1498), .ZN(n1013) );
  AND2_X1 U1065 ( .A1(G107), .A2(n1013), .ZN(n981) );
  NAND2_X1 U1066 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1067 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1068 ( .A(n985), .B(KEYINPUT17), .ZN(n988) );
  NOR2_X1 U1069 ( .A1(G20), .A2(n986), .ZN(n1405) );
  NAND2_X1 U1070 ( .A1(n1405), .A2(G87), .ZN(n987) );
  NAND2_X1 U1071 ( .A1(n988), .A2(n987), .ZN(n991) );
  INV_X1 U1072 ( .A(KEYINPUT4), .ZN(n989) );
  NAND2_X1 U1073 ( .A1(n1279), .A2(G20), .ZN(n1092) );
  NOR2_X1 U1074 ( .A1(G107), .A2(n1305), .ZN(n990) );
  NOR2_X2 U1075 ( .A1(n991), .A2(n990), .ZN(n1003) );
  NOR2_X1 U1076 ( .A1(n992), .A2(n1003), .ZN(n995) );
  XNOR2_X1 U1077 ( .A(n993), .B(KEYINPUT15), .ZN(n994) );
  AND2_X2 U1078 ( .A1(n995), .A2(n994), .ZN(n1066) );
  INV_X1 U1079 ( .A(n1003), .ZN(n999) );
  NAND2_X1 U1080 ( .A1(G200), .A2(n1122), .ZN(n997) );
  INV_X1 U1081 ( .A(n1122), .ZN(n1117) );
  NAND2_X1 U1082 ( .A1(G190), .A2(n1117), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  NOR2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X2 U1085 ( .A(n1001), .B(KEYINPUT0), .ZN(n1111) );
  NOR2_X1 U1086 ( .A1(G20), .A2(n1866), .ZN(n1190) );
  NAND2_X1 U1087 ( .A1(n1190), .A2(G213), .ZN(n1002) );
  NOR2_X1 U1088 ( .A1(G1), .A2(n1002), .ZN(n1458) );
  NAND2_X1 U1089 ( .A1(n1458), .A2(G343), .ZN(n1292) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1292), .ZN(n1070) );
  NAND2_X1 U1091 ( .A1(n1393), .A2(G264), .ZN(n1004) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1042), .ZN(n1010) );
  NAND2_X1 U1093 ( .A1(n1046), .A2(G270), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(KEYINPUT10), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1389), .A2(G303), .ZN(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n960), .A2(G257), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1119) );
  NAND2_X1 U1100 ( .A1(n1119), .A2(n1400), .ZN(n1023) );
  NAND2_X1 U1101 ( .A1(n1345), .A2(n1013), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(n1279), .A2(n1014), .ZN(n1091) );
  BUF_X1 U1103 ( .A(n1015), .Z(n1344) );
  OR2_X1 U1104 ( .A1(n1091), .A2(n1344), .ZN(n1016) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(G116), .ZN(n1022) );
  NAND2_X1 U1106 ( .A1(G283), .A2(n1401), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1405), .A2(G97), .ZN(n1017) );
  NAND2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(G116), .A2(n1345), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1031) );
  NAND2_X1 U1112 ( .A1(n1023), .A2(n1031), .ZN(n1025) );
  NOR2_X1 U1113 ( .A1(G179), .A2(n1119), .ZN(n1024) );
  AND2_X1 U1114 ( .A1(n1292), .A2(n1067), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1070), .A2(n1026), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(n1111), .B(n1027), .ZN(n1038) );
  INV_X1 U1117 ( .A(n1292), .ZN(n1687) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1687), .ZN(n1035) );
  INV_X1 U1119 ( .A(KEYINPUT11), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(G200), .A2(n1119), .ZN(n1029) );
  INV_X1 U1121 ( .A(n1119), .ZN(n1126) );
  NAND2_X1 U1122 ( .A1(G190), .A2(n1126), .ZN(n1028) );
  NAND2_X1 U1123 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1124 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1125 ( .A1(n1067), .A2(n1032), .ZN(n1033) );
  XNOR2_X1 U1126 ( .A(n1034), .B(n1033), .ZN(n1110) );
  NAND2_X1 U1127 ( .A1(n1035), .A2(n1110), .ZN(n1037) );
  NAND2_X1 U1128 ( .A1(n1067), .A2(n1687), .ZN(n1036) );
  NAND2_X1 U1129 ( .A1(n1037), .A2(n1036), .ZN(n1256) );
  AND2_X1 U1130 ( .A1(G330), .A2(n1256), .ZN(n1074) );
  XOR2_X1 U1131 ( .A(n1038), .B(n1074), .Z(n1669) );
  NAND2_X1 U1132 ( .A1(n960), .A2(G244), .ZN(n1040) );
  NAND2_X1 U1133 ( .A1(n1393), .A2(G250), .ZN(n1039) );
  NAND2_X1 U1134 ( .A1(n1040), .A2(n1039), .ZN(n1044) );
  NAND2_X1 U1135 ( .A1(n1389), .A2(G283), .ZN(n1041) );
  NAND2_X1 U1136 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  NOR2_X1 U1137 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  XNOR2_X1 U1138 ( .A(n1045), .B(KEYINPUT12), .ZN(n1048) );
  NAND2_X1 U1139 ( .A1(n1046), .A2(G257), .ZN(n1047) );
  NAND2_X1 U1140 ( .A1(n1048), .A2(n1047), .ZN(n1123) );
  NOR2_X1 U1141 ( .A1(G179), .A2(n1123), .ZN(n1050) );
  AND2_X1 U1142 ( .A1(n1400), .A2(n1123), .ZN(n1049) );
  NOR2_X1 U1143 ( .A1(n1050), .A2(n1049), .ZN(n1060) );
  NAND2_X1 U1144 ( .A1(G77), .A2(n1405), .ZN(n1052) );
  INV_X1 U1145 ( .A(G107), .ZN(n1762) );
  XOR2_X1 U1146 ( .A(n1762), .B(G97), .Z(n1888) );
  NAND2_X1 U1147 ( .A1(n1888), .A2(n1344), .ZN(n1051) );
  NAND2_X1 U1148 ( .A1(n1052), .A2(n1051), .ZN(n1057) );
  INV_X1 U1149 ( .A(n1401), .ZN(n1273) );
  NOR2_X1 U1150 ( .A1(n1762), .A2(n1273), .ZN(n1054) );
  NOR2_X1 U1151 ( .A1(G97), .A2(n1345), .ZN(n1053) );
  NOR2_X1 U1152 ( .A1(n1054), .A2(n1053), .ZN(n1055) );
  XNOR2_X1 U1153 ( .A(n1055), .B(KEYINPUT13), .ZN(n1056) );
  NOR2_X1 U1154 ( .A1(n1057), .A2(n1056), .ZN(n1059) );
  NAND2_X1 U1155 ( .A1(n1091), .A2(G97), .ZN(n1058) );
  NAND2_X1 U1156 ( .A1(n1059), .A2(n1058), .ZN(n1065) );
  NAND2_X1 U1157 ( .A1(n1060), .A2(n1065), .ZN(n1679) );
  INV_X1 U1158 ( .A(G190), .ZN(n1420) );
  NOR2_X1 U1159 ( .A1(n1420), .A2(n1123), .ZN(n1061) );
  NOR2_X1 U1160 ( .A1(n1065), .A2(n1061), .ZN(n1063) );
  NAND2_X1 U1161 ( .A1(G200), .A2(n1123), .ZN(n1062) );
  NAND2_X1 U1162 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  NAND2_X1 U1163 ( .A1(n1679), .A2(n1064), .ZN(n1144) );
  AND2_X1 U1164 ( .A1(n1065), .A2(n1687), .ZN(n1145) );
  AND2_X2 U1165 ( .A1(n1067), .A2(n1111), .ZN(n1068) );
  NOR2_X1 U1166 ( .A1(n1066), .A2(n1068), .ZN(n1077) );
  NOR2_X1 U1167 ( .A1(n1687), .A2(n1077), .ZN(n1854) );
  NOR2_X1 U1168 ( .A1(n1145), .A2(n1854), .ZN(n1069) );
  XOR2_X1 U1169 ( .A(n1144), .B(n1069), .Z(n1075) );
  NAND2_X1 U1170 ( .A1(n1687), .A2(n1066), .ZN(n1073) );
  INV_X1 U1171 ( .A(n1070), .ZN(n1071) );
  NAND2_X1 U1172 ( .A1(n1071), .A2(n1111), .ZN(n1072) );
  NAND2_X1 U1173 ( .A1(n1073), .A2(n1072), .ZN(n1662) );
  NAND2_X1 U1174 ( .A1(n1074), .A2(n1662), .ZN(n1855) );
  XNOR2_X1 U1175 ( .A(n1075), .B(n1855), .ZN(n1202) );
  NAND2_X1 U1176 ( .A1(n1669), .A2(n1202), .ZN(n1076) );
  XNOR2_X1 U1177 ( .A(KEYINPUT52), .B(n1076), .ZN(n1675) );
  NAND2_X1 U1178 ( .A1(n1863), .A2(n1675), .ZN(n1136) );
  OR2_X1 U1179 ( .A1(n1144), .A2(n1077), .ZN(n1678) );
  NAND2_X1 U1180 ( .A1(G274), .A2(n1078), .ZN(n1080) );
  NAND2_X1 U1181 ( .A1(G116), .A2(n1389), .ZN(n1079) );
  NAND2_X1 U1182 ( .A1(n1080), .A2(n1079), .ZN(n1084) );
  NAND2_X1 U1183 ( .A1(G250), .A2(n1081), .ZN(n1082) );
  NOR2_X1 U1184 ( .A1(n1269), .A2(n1082), .ZN(n1083) );
  NOR2_X1 U1185 ( .A1(n1084), .A2(n1083), .ZN(n1088) );
  NAND2_X1 U1186 ( .A1(G244), .A2(n1393), .ZN(n1086) );
  NAND2_X1 U1187 ( .A1(G238), .A2(n960), .ZN(n1085) );
  NAND2_X1 U1188 ( .A1(n1086), .A2(n1085), .ZN(n1087) );
  NAND2_X1 U1189 ( .A1(n1088), .A2(n962), .ZN(n1115) );
  INV_X1 U1190 ( .A(G179), .ZN(n1372) );
  NOR2_X1 U1191 ( .A1(n1115), .A2(n1372), .ZN(n1090) );
  NOR2_X1 U1192 ( .A1(n1125), .A2(n1400), .ZN(n1089) );
  OR2_X1 U1193 ( .A1(n1090), .A2(n1089), .ZN(n1689) );
  NAND2_X1 U1194 ( .A1(G87), .A2(n1091), .ZN(n1093) );
  XNOR2_X1 U1195 ( .A(KEYINPUT4), .B(n1092), .ZN(n1409) );
  NAND2_X1 U1196 ( .A1(n1093), .A2(n1409), .ZN(n1094) );
  NOR2_X1 U1197 ( .A1(G107), .A2(G97), .ZN(n1205) );
  INV_X1 U1198 ( .A(G87), .ZN(n1272) );
  NAND2_X1 U1199 ( .A1(n1205), .A2(n1272), .ZN(n1642) );
  NAND2_X1 U1200 ( .A1(n1094), .A2(n1642), .ZN(n1095) );
  XNOR2_X1 U1201 ( .A(n1095), .B(KEYINPUT9), .ZN(n1097) );
  NOR2_X1 U1202 ( .A1(n1345), .A2(G87), .ZN(n1096) );
  NOR2_X1 U1203 ( .A1(n1097), .A2(n1096), .ZN(n1099) );
  NAND2_X1 U1204 ( .A1(G97), .A2(n1401), .ZN(n1098) );
  NAND2_X1 U1205 ( .A1(n1099), .A2(n1098), .ZN(n1101) );
  AND2_X1 U1206 ( .A1(n1405), .A2(G68), .ZN(n1100) );
  OR2_X1 U1207 ( .A1(n1101), .A2(n1100), .ZN(n1686) );
  AND2_X1 U1208 ( .A1(n1679), .A2(n1106), .ZN(n1102) );
  NAND2_X1 U1209 ( .A1(n1678), .A2(n1102), .ZN(n1109) );
  INV_X1 U1210 ( .A(n1106), .ZN(n1107) );
  NAND2_X1 U1211 ( .A1(G200), .A2(n1115), .ZN(n1104) );
  NAND2_X1 U1212 ( .A1(n1125), .A2(G190), .ZN(n1103) );
  NAND2_X1 U1213 ( .A1(n1104), .A2(n1103), .ZN(n1105) );
  OR2_X1 U1214 ( .A1(n1686), .A2(n1105), .ZN(n1682) );
  OR2_X1 U1215 ( .A1(n1107), .A2(n963), .ZN(n1108) );
  AND2_X2 U1216 ( .A1(n1109), .A2(n1108), .ZN(n1286) );
  NAND2_X1 U1217 ( .A1(n1292), .A2(n1286), .ZN(n1442) );
  AND2_X1 U1218 ( .A1(n1111), .A2(n1110), .ZN(n1114) );
  NAND2_X1 U1219 ( .A1(n1853), .A2(n1292), .ZN(n1133) );
  NOR2_X1 U1220 ( .A1(n1115), .A2(n1123), .ZN(n1116) );
  XNOR2_X1 U1221 ( .A(KEYINPUT18), .B(n1116), .ZN(n1121) );
  NAND2_X1 U1222 ( .A1(G179), .A2(n1117), .ZN(n1118) );
  NOR2_X1 U1223 ( .A1(n1119), .A2(n1118), .ZN(n1120) );
  NAND2_X1 U1224 ( .A1(n1121), .A2(n1120), .ZN(n1130) );
  NAND2_X1 U1225 ( .A1(n1123), .A2(n1122), .ZN(n1124) );
  NOR2_X1 U1226 ( .A1(n1125), .A2(n1124), .ZN(n1128) );
  NOR2_X1 U1227 ( .A1(n1126), .A2(G179), .ZN(n1127) );
  NAND2_X1 U1228 ( .A1(n1128), .A2(n1127), .ZN(n1129) );
  NAND2_X1 U1229 ( .A1(n1130), .A2(n1129), .ZN(n1131) );
  NAND2_X1 U1230 ( .A1(n1687), .A2(n1131), .ZN(n1132) );
  NAND2_X1 U1231 ( .A1(G330), .A2(n1430), .ZN(n1340) );
  NAND2_X1 U1232 ( .A1(n1442), .A2(n1340), .ZN(n1673) );
  INV_X1 U1233 ( .A(n1673), .ZN(n1857) );
  AND2_X1 U1234 ( .A1(n1669), .A2(n1857), .ZN(n1134) );
  NOR2_X1 U1235 ( .A1(n1202), .A2(n1134), .ZN(n1135) );
  NOR2_X1 U1236 ( .A1(n1136), .A2(n1135), .ZN(n1199) );
  INV_X1 U1237 ( .A(n1828), .ZN(n1206) );
  NAND2_X1 U1238 ( .A1(G33), .A2(n1206), .ZN(n1137) );
  XNOR2_X1 U1239 ( .A(n1137), .B(KEYINPUT24), .ZN(n1700) );
  XNOR2_X1 U1240 ( .A(n1888), .B(KEYINPUT51), .ZN(n1139) );
  INV_X1 U1241 ( .A(G116), .ZN(n1889) );
  XOR2_X1 U1242 ( .A(n1889), .B(G87), .Z(n1138) );
  XNOR2_X1 U1243 ( .A(n1139), .B(n1138), .ZN(n1903) );
  NOR2_X1 U1244 ( .A1(n1700), .A2(n1903), .ZN(n1143) );
  NAND2_X1 U1245 ( .A1(n1866), .A2(n1498), .ZN(n1654) );
  NOR2_X1 U1246 ( .A1(n1654), .A2(G20), .ZN(n1233) );
  NOR2_X1 U1247 ( .A1(G169), .A2(n1827), .ZN(n1140) );
  NOR2_X1 U1248 ( .A1(n1826), .A2(n1140), .ZN(n1239) );
  NOR2_X1 U1249 ( .A1(n1233), .A2(n1239), .ZN(n1697) );
  NAND2_X1 U1250 ( .A1(G97), .A2(n1828), .ZN(n1141) );
  NAND2_X1 U1251 ( .A1(n1697), .A2(n1141), .ZN(n1142) );
  NOR2_X1 U1252 ( .A1(n1143), .A2(n1142), .ZN(n1197) );
  NOR2_X1 U1253 ( .A1(n1145), .A2(n1144), .ZN(n1147) );
  NOR2_X1 U1254 ( .A1(n1679), .A2(n1292), .ZN(n1146) );
  NOR2_X1 U1255 ( .A1(n1147), .A2(n1146), .ZN(n1677) );
  NAND2_X1 U1256 ( .A1(n1677), .A2(n1233), .ZN(n1195) );
  INV_X1 U1257 ( .A(n1239), .ZN(n1753) );
  NOR2_X1 U1258 ( .A1(n1827), .A2(n1372), .ZN(n1156) );
  INV_X1 U1259 ( .A(G200), .ZN(n1366) );
  NOR2_X1 U1260 ( .A1(n1366), .A2(n1420), .ZN(n1148) );
  AND2_X1 U1261 ( .A1(n1156), .A2(n1148), .ZN(n1782) );
  NAND2_X1 U1262 ( .A1(n1782), .A2(G317), .ZN(n1150) );
  NOR2_X1 U1263 ( .A1(n1827), .A2(G179), .ZN(n1153) );
  NAND2_X1 U1264 ( .A1(n1153), .A2(n1148), .ZN(n1761) );
  INV_X1 U1265 ( .A(n1761), .ZN(n1786) );
  NAND2_X1 U1266 ( .A1(n1786), .A2(G283), .ZN(n1149) );
  NAND2_X1 U1267 ( .A1(n1150), .A2(n1149), .ZN(n1151) );
  XOR2_X1 U1268 ( .A(KEYINPUT59), .B(n1151), .Z(n1170) );
  NOR2_X1 U1269 ( .A1(G200), .A2(n1420), .ZN(n1157) );
  AND2_X1 U1270 ( .A1(n1156), .A2(n1157), .ZN(n1772) );
  NAND2_X1 U1271 ( .A1(G311), .A2(n1772), .ZN(n1152) );
  NAND2_X1 U1272 ( .A1(G33), .A2(n1152), .ZN(n1167) );
  NAND2_X1 U1273 ( .A1(n1153), .A2(n1420), .ZN(n1154) );
  NOR2_X1 U1274 ( .A1(n1366), .A2(n1154), .ZN(n1626) );
  NAND2_X1 U1275 ( .A1(G107), .A2(n1626), .ZN(n1218) );
  NAND2_X1 U1276 ( .A1(n1778), .A2(G322), .ZN(n1155) );
  NAND2_X1 U1277 ( .A1(n1218), .A2(n1155), .ZN(n1162) );
  NAND2_X1 U1278 ( .A1(n1156), .A2(n1420), .ZN(n1163) );
  NAND2_X1 U1279 ( .A1(G294), .A2(n1783), .ZN(n1160) );
  NAND2_X1 U1280 ( .A1(n1157), .A2(n1372), .ZN(n1158) );
  NAND2_X1 U1281 ( .A1(G20), .A2(n1158), .ZN(n1787) );
  NAND2_X1 U1282 ( .A1(G116), .A2(n1787), .ZN(n1159) );
  NAND2_X1 U1283 ( .A1(n1160), .A2(n1159), .ZN(n1161) );
  NOR2_X1 U1284 ( .A1(n1162), .A2(n1161), .ZN(n1165) );
  NAND2_X1 U1285 ( .A1(G303), .A2(n1775), .ZN(n1164) );
  NAND2_X1 U1286 ( .A1(n1165), .A2(n1164), .ZN(n1166) );
  NOR2_X1 U1287 ( .A1(n1167), .A2(n1166), .ZN(n1168) );
  XOR2_X1 U1288 ( .A(KEYINPUT58), .B(n1168), .Z(n1169) );
  NOR2_X1 U1289 ( .A1(n1170), .A2(n1169), .ZN(n1188) );
  NAND2_X1 U1290 ( .A1(G159), .A2(n1772), .ZN(n1172) );
  NAND2_X1 U1291 ( .A1(G58), .A2(n1783), .ZN(n1171) );
  NAND2_X1 U1292 ( .A1(n1172), .A2(n1171), .ZN(n1174) );
  NAND2_X1 U1293 ( .A1(G77), .A2(n1787), .ZN(n1536) );
  NAND2_X1 U1294 ( .A1(n1498), .A2(n1536), .ZN(n1173) );
  NOR2_X1 U1295 ( .A1(n1174), .A2(n1173), .ZN(n1184) );
  NAND2_X1 U1296 ( .A1(G143), .A2(n1778), .ZN(n1176) );
  NAND2_X1 U1297 ( .A1(G50), .A2(n1775), .ZN(n1175) );
  NAND2_X1 U1298 ( .A1(n1176), .A2(n1175), .ZN(n1182) );
  NAND2_X1 U1299 ( .A1(n1782), .A2(G150), .ZN(n1177) );
  XNOR2_X1 U1300 ( .A(n1177), .B(KEYINPUT56), .ZN(n1179) );
  NAND2_X1 U1301 ( .A1(n1786), .A2(G68), .ZN(n1178) );
  NAND2_X1 U1302 ( .A1(n1179), .A2(n1178), .ZN(n1180) );
  XOR2_X1 U1303 ( .A(KEYINPUT57), .B(n1180), .Z(n1181) );
  NOR2_X1 U1304 ( .A1(n1182), .A2(n1181), .ZN(n1183) );
  NAND2_X1 U1305 ( .A1(n1184), .A2(n1183), .ZN(n1186) );
  NAND2_X1 U1306 ( .A1(n1626), .A2(G87), .ZN(n1185) );
  XOR2_X1 U1307 ( .A(KEYINPUT22), .B(n1185), .Z(n1767) );
  NOR2_X1 U1308 ( .A1(n1186), .A2(n1767), .ZN(n1187) );
  NOR2_X1 U1309 ( .A1(n1188), .A2(n1187), .ZN(n1189) );
  NOR2_X1 U1310 ( .A1(n1753), .A2(n1189), .ZN(n1193) );
  NAND2_X1 U1311 ( .A1(G45), .A2(n1190), .ZN(n1191) );
  NAND2_X1 U1312 ( .A1(G1), .A2(n1191), .ZN(n1192) );
  NOR2_X1 U1313 ( .A1(n1672), .A2(n1863), .ZN(n1620) );
  INV_X1 U1314 ( .A(n1620), .ZN(n1802) );
  NOR2_X1 U1315 ( .A1(n1193), .A2(n1802), .ZN(n1194) );
  NAND2_X1 U1316 ( .A1(n1195), .A2(n1194), .ZN(n1196) );
  NOR2_X1 U1317 ( .A1(n1197), .A2(n1196), .ZN(n1198) );
  NOR2_X1 U1318 ( .A1(n1199), .A2(n1198), .ZN(n1204) );
  INV_X1 U1319 ( .A(n1672), .ZN(n1201) );
  NAND2_X1 U1320 ( .A1(n1863), .A2(n1673), .ZN(n1200) );
  NAND2_X1 U1321 ( .A1(n1201), .A2(n1200), .ZN(n1668) );
  NAND2_X1 U1322 ( .A1(n1202), .A2(n1668), .ZN(n1203) );
  NAND2_X1 U1323 ( .A1(n1204), .A2(n1203), .ZN(G390) );
  OR2_X1 U1324 ( .A1(n1272), .A2(n1205), .ZN(G355) );
  INV_X1 U1325 ( .A(n1654), .ZN(n1747) );
  NAND2_X1 U1326 ( .A1(G355), .A2(n1747), .ZN(n1215) );
  NOR2_X1 U1327 ( .A1(n1206), .A2(G116), .ZN(n1207) );
  XNOR2_X1 U1328 ( .A(n1207), .B(KEYINPUT60), .ZN(n1213) );
  INV_X1 U1329 ( .A(G77), .ZN(n1881) );
  XOR2_X1 U1330 ( .A(n1881), .B(G50), .Z(n1208) );
  XNOR2_X1 U1331 ( .A(G68), .B(G58), .ZN(n1343) );
  XNOR2_X1 U1332 ( .A(n1208), .B(n1343), .ZN(n1902) );
  NAND2_X1 U1333 ( .A1(G45), .A2(n1902), .ZN(n1210) );
  NOR2_X1 U1334 ( .A1(G68), .A2(G58), .ZN(n1895) );
  INV_X1 U1335 ( .A(G50), .ZN(n1894) );
  NOR2_X1 U1336 ( .A1(n1895), .A2(n1894), .ZN(n1862) );
  NAND2_X1 U1337 ( .A1(n1862), .A2(n1650), .ZN(n1209) );
  NAND2_X1 U1338 ( .A1(n1210), .A2(n1209), .ZN(n1211) );
  NOR2_X1 U1339 ( .A1(n1211), .A2(n1700), .ZN(n1212) );
  NOR2_X1 U1340 ( .A1(n1213), .A2(n1212), .ZN(n1214) );
  NAND2_X1 U1341 ( .A1(n1215), .A2(n1214), .ZN(n1216) );
  NAND2_X1 U1342 ( .A1(n1216), .A2(n1697), .ZN(n1232) );
  NAND2_X1 U1343 ( .A1(n1772), .A2(G58), .ZN(n1217) );
  NAND2_X1 U1344 ( .A1(n1218), .A2(n1217), .ZN(n1226) );
  NAND2_X1 U1345 ( .A1(G159), .A2(n1778), .ZN(n1220) );
  NAND2_X1 U1346 ( .A1(n1775), .A2(G68), .ZN(n1219) );
  NAND2_X1 U1347 ( .A1(n1220), .A2(n1219), .ZN(n1223) );
  NAND2_X1 U1348 ( .A1(G97), .A2(n1787), .ZN(n1754) );
  NAND2_X1 U1349 ( .A1(G77), .A2(n1783), .ZN(n1221) );
  NAND2_X1 U1350 ( .A1(n1754), .A2(n1221), .ZN(n1222) );
  NOR2_X1 U1351 ( .A1(n1223), .A2(n1222), .ZN(n1224) );
  XNOR2_X1 U1352 ( .A(KEYINPUT61), .B(n1224), .ZN(n1225) );
  NOR2_X1 U1353 ( .A1(n1226), .A2(n1225), .ZN(n1230) );
  NOR2_X1 U1354 ( .A1(n1753), .A2(G33), .ZN(n1777) );
  INV_X1 U1355 ( .A(n1777), .ZN(n1709) );
  NAND2_X1 U1356 ( .A1(G87), .A2(n1786), .ZN(n1539) );
  NAND2_X1 U1357 ( .A1(n1782), .A2(G50), .ZN(n1227) );
  NAND2_X1 U1358 ( .A1(n1539), .A2(n1227), .ZN(n1228) );
  NOR2_X1 U1359 ( .A1(n1709), .A2(n1228), .ZN(n1229) );
  NAND2_X1 U1360 ( .A1(n1230), .A2(n1229), .ZN(n1231) );
  NAND2_X1 U1361 ( .A1(n1232), .A2(n1231), .ZN(n1236) );
  INV_X1 U1362 ( .A(n1233), .ZN(n1741) );
  NOR2_X1 U1363 ( .A1(n1741), .A2(n1256), .ZN(n1234) );
  XNOR2_X1 U1364 ( .A(KEYINPUT62), .B(n1234), .ZN(n1235) );
  NOR2_X1 U1365 ( .A1(n1236), .A2(n1235), .ZN(n1255) );
  NAND2_X1 U1366 ( .A1(G311), .A2(n1783), .ZN(n1238) );
  NAND2_X1 U1367 ( .A1(n1786), .A2(G303), .ZN(n1237) );
  NAND2_X1 U1368 ( .A1(n1238), .A2(n1237), .ZN(n1252) );
  NAND2_X1 U1369 ( .A1(G33), .A2(n1239), .ZN(n1624) );
  NAND2_X1 U1370 ( .A1(G322), .A2(n1772), .ZN(n1241) );
  NAND2_X1 U1371 ( .A1(G326), .A2(n1782), .ZN(n1240) );
  NAND2_X1 U1372 ( .A1(n1241), .A2(n1240), .ZN(n1242) );
  NOR2_X1 U1373 ( .A1(n1624), .A2(n1242), .ZN(n1250) );
  NAND2_X1 U1374 ( .A1(n1778), .A2(G329), .ZN(n1244) );
  NAND2_X1 U1375 ( .A1(G294), .A2(n1787), .ZN(n1243) );
  NAND2_X1 U1376 ( .A1(n1244), .A2(n1243), .ZN(n1248) );
  NAND2_X1 U1377 ( .A1(G317), .A2(n1775), .ZN(n1246) );
  NAND2_X1 U1378 ( .A1(n1626), .A2(G283), .ZN(n1245) );
  NAND2_X1 U1379 ( .A1(n1246), .A2(n1245), .ZN(n1247) );
  NOR2_X1 U1380 ( .A1(n1248), .A2(n1247), .ZN(n1249) );
  NAND2_X1 U1381 ( .A1(n1250), .A2(n1249), .ZN(n1251) );
  NOR2_X1 U1382 ( .A1(n1252), .A2(n1251), .ZN(n1253) );
  NOR2_X1 U1383 ( .A1(n1802), .A2(n1253), .ZN(n1254) );
  NAND2_X1 U1384 ( .A1(n1255), .A2(n1254), .ZN(n1259) );
  XOR2_X1 U1385 ( .A(G330), .B(n1256), .Z(n1257) );
  NAND2_X1 U1386 ( .A1(n1257), .A2(n1802), .ZN(n1258) );
  NAND2_X1 U1387 ( .A1(n1259), .A2(n1258), .ZN(G396) );
  NAND2_X1 U1388 ( .A1(n1389), .A2(G107), .ZN(n1261) );
  NAND2_X1 U1389 ( .A1(G232), .A2(n960), .ZN(n1260) );
  NAND2_X1 U1390 ( .A1(n1261), .A2(n1260), .ZN(n1264) );
  NAND2_X1 U1391 ( .A1(G238), .A2(n1393), .ZN(n1262) );
  XOR2_X1 U1392 ( .A(KEYINPUT6), .B(n1262), .Z(n1263) );
  NOR2_X1 U1393 ( .A1(n1264), .A2(n1263), .ZN(n1266) );
  NOR2_X1 U1394 ( .A1(G45), .A2(G41), .ZN(n1265) );
  NOR2_X1 U1395 ( .A1(G1), .A2(n1265), .ZN(n1268) );
  NAND2_X1 U1396 ( .A1(G274), .A2(n1268), .ZN(n1391) );
  NAND2_X1 U1397 ( .A1(n1266), .A2(n1391), .ZN(n1267) );
  XNOR2_X1 U1398 ( .A(n1267), .B(KEYINPUT7), .ZN(n1271) );
  NOR2_X1 U1399 ( .A1(n1269), .A2(n1268), .ZN(n1392) );
  NAND2_X1 U1400 ( .A1(n1392), .A2(G244), .ZN(n1270) );
  NAND2_X1 U1401 ( .A1(n1271), .A2(n1270), .ZN(n1287) );
  NOR2_X1 U1402 ( .A1(n1420), .A2(n1287), .ZN(n1283) );
  NOR2_X1 U1403 ( .A1(G77), .A2(n1345), .ZN(n1275) );
  NOR2_X1 U1404 ( .A1(n1273), .A2(n1272), .ZN(n1274) );
  NOR2_X1 U1405 ( .A1(n1275), .A2(n1274), .ZN(n1277) );
  NAND2_X1 U1406 ( .A1(n1405), .A2(G58), .ZN(n1276) );
  NAND2_X1 U1407 ( .A1(n1277), .A2(n1276), .ZN(n1281) );
  NOR2_X1 U1408 ( .A1(n1279), .A2(n1278), .ZN(n1348) );
  NOR2_X1 U1409 ( .A1(n1348), .A2(n1344), .ZN(n1408) );
  NOR2_X1 U1410 ( .A1(n1408), .A2(n1881), .ZN(n1280) );
  NOR2_X1 U1411 ( .A1(n1281), .A2(n1280), .ZN(n1293) );
  INV_X1 U1412 ( .A(n1293), .ZN(n1282) );
  NOR2_X1 U1413 ( .A1(n1283), .A2(n1282), .ZN(n1285) );
  NAND2_X1 U1414 ( .A1(G200), .A2(n1287), .ZN(n1284) );
  NAND2_X1 U1415 ( .A1(n1285), .A2(n1284), .ZN(n1295) );
  NAND2_X1 U1416 ( .A1(n1295), .A2(n1286), .ZN(n1290) );
  NAND2_X1 U1417 ( .A1(G169), .A2(n1287), .ZN(n1289) );
  OR2_X1 U1418 ( .A1(n1372), .A2(n1287), .ZN(n1288) );
  AND2_X1 U1419 ( .A1(n1289), .A2(n1288), .ZN(n1299) );
  NOR2_X1 U1420 ( .A1(n1299), .A2(n1293), .ZN(n1434) );
  INV_X1 U1421 ( .A(n1434), .ZN(n1296) );
  NAND2_X1 U1422 ( .A1(n1290), .A2(n1296), .ZN(n1291) );
  NAND2_X1 U1423 ( .A1(n1291), .A2(n1292), .ZN(n1335) );
  NOR2_X1 U1424 ( .A1(n1293), .A2(n1292), .ZN(n1294) );
  XNOR2_X1 U1425 ( .A(KEYINPUT5), .B(n1294), .ZN(n1298) );
  INV_X1 U1426 ( .A(n1298), .ZN(n1297) );
  NAND2_X1 U1427 ( .A1(n1296), .A2(n1295), .ZN(n1426) );
  NOR2_X1 U1428 ( .A1(n1297), .A2(n1426), .ZN(n1301) );
  NOR2_X1 U1429 ( .A1(n1299), .A2(n1298), .ZN(n1300) );
  NOR2_X1 U1430 ( .A1(n1301), .A2(n1300), .ZN(n1801) );
  OR2_X1 U1431 ( .A1(n1801), .A2(n1340), .ZN(n1302) );
  NAND2_X1 U1432 ( .A1(n1335), .A2(n1302), .ZN(n1334) );
  NAND2_X1 U1433 ( .A1(G77), .A2(n1401), .ZN(n1304) );
  NAND2_X1 U1434 ( .A1(G50), .A2(n1405), .ZN(n1303) );
  NAND2_X1 U1435 ( .A1(n1304), .A2(n1303), .ZN(n1307) );
  NOR2_X1 U1436 ( .A1(G68), .A2(n1305), .ZN(n1306) );
  NOR2_X1 U1437 ( .A1(n1307), .A2(n1306), .ZN(n1309) );
  NAND2_X1 U1438 ( .A1(G68), .A2(n1348), .ZN(n1308) );
  NAND2_X1 U1439 ( .A1(n1309), .A2(n1308), .ZN(n1321) );
  NAND2_X1 U1440 ( .A1(n1321), .A2(n1687), .ZN(n1329) );
  NAND2_X1 U1441 ( .A1(n1389), .A2(G97), .ZN(n1310) );
  NAND2_X1 U1442 ( .A1(n1391), .A2(n1310), .ZN(n1314) );
  NAND2_X1 U1443 ( .A1(G232), .A2(n1393), .ZN(n1312) );
  NAND2_X1 U1444 ( .A1(G226), .A2(n960), .ZN(n1311) );
  NAND2_X1 U1445 ( .A1(n1312), .A2(n1311), .ZN(n1313) );
  NOR2_X1 U1446 ( .A1(n1314), .A2(n1313), .ZN(n1316) );
  NAND2_X1 U1447 ( .A1(G238), .A2(n1392), .ZN(n1315) );
  NAND2_X1 U1448 ( .A1(n1316), .A2(n1315), .ZN(n1322) );
  NAND2_X1 U1449 ( .A1(n1400), .A2(n1322), .ZN(n1317) );
  NAND2_X1 U1450 ( .A1(n1321), .A2(n1317), .ZN(n1319) );
  NOR2_X1 U1451 ( .A1(G179), .A2(n1322), .ZN(n1318) );
  NOR2_X1 U1452 ( .A1(n1319), .A2(n1318), .ZN(n1336) );
  NAND2_X1 U1453 ( .A1(n1322), .A2(G200), .ZN(n1320) );
  XNOR2_X1 U1454 ( .A(n1320), .B(KEYINPUT27), .ZN(n1327) );
  INV_X1 U1455 ( .A(n1321), .ZN(n1325) );
  NOR2_X1 U1456 ( .A1(n1420), .A2(n1322), .ZN(n1323) );
  XOR2_X1 U1457 ( .A(KEYINPUT28), .B(n1323), .Z(n1324) );
  NAND2_X1 U1458 ( .A1(n1325), .A2(n1324), .ZN(n1326) );
  NOR2_X1 U1459 ( .A1(n1327), .A2(n1326), .ZN(n1328) );
  NOR2_X1 U1460 ( .A1(n1336), .A2(n1328), .ZN(n1433) );
  NAND2_X1 U1461 ( .A1(n1329), .A2(n1433), .ZN(n1331) );
  NAND2_X1 U1462 ( .A1(n1336), .A2(n1687), .ZN(n1330) );
  NAND2_X1 U1463 ( .A1(n1331), .A2(n1330), .ZN(n1332) );
  XNOR2_X1 U1464 ( .A(KEYINPUT29), .B(n1332), .ZN(n1598) );
  INV_X1 U1465 ( .A(n1560), .ZN(n1563) );
  NOR2_X1 U1466 ( .A1(n1335), .A2(n1598), .ZN(n1338) );
  INV_X1 U1467 ( .A(n1336), .ZN(n1436) );
  NOR2_X1 U1468 ( .A1(n1687), .A2(n1436), .ZN(n1337) );
  NOR2_X1 U1469 ( .A1(n1338), .A2(n1337), .ZN(n1456) );
  OR2_X1 U1470 ( .A1(n1598), .A2(n1801), .ZN(n1339) );
  XNOR2_X1 U1471 ( .A(KEYINPUT39), .B(n1341), .ZN(n1342) );
  NAND2_X1 U1472 ( .A1(n1456), .A2(n1342), .ZN(n1385) );
  NAND2_X1 U1473 ( .A1(n1344), .A2(n1343), .ZN(n1354) );
  NAND2_X1 U1474 ( .A1(n1405), .A2(G159), .ZN(n1347) );
  OR2_X1 U1475 ( .A1(n1345), .A2(G58), .ZN(n1346) );
  NAND2_X1 U1476 ( .A1(n1347), .A2(n1346), .ZN(n1352) );
  NAND2_X1 U1477 ( .A1(n1348), .A2(G58), .ZN(n1350) );
  NAND2_X1 U1478 ( .A1(n1401), .A2(G68), .ZN(n1349) );
  NAND2_X1 U1479 ( .A1(n1350), .A2(n1349), .ZN(n1351) );
  NOR2_X1 U1480 ( .A1(n1352), .A2(n1351), .ZN(n1353) );
  NAND2_X1 U1481 ( .A1(n1354), .A2(n1353), .ZN(n1355) );
  XOR2_X1 U1482 ( .A(n1355), .B(KEYINPUT30), .Z(n1378) );
  INV_X1 U1483 ( .A(n1378), .ZN(n1381) );
  NAND2_X1 U1484 ( .A1(n1392), .A2(G232), .ZN(n1358) );
  NAND2_X1 U1485 ( .A1(G87), .A2(n1389), .ZN(n1356) );
  XOR2_X1 U1486 ( .A(KEYINPUT31), .B(n1356), .Z(n1357) );
  NAND2_X1 U1487 ( .A1(n1358), .A2(n1357), .ZN(n1365) );
  NAND2_X1 U1488 ( .A1(n1393), .A2(G226), .ZN(n1359) );
  XNOR2_X1 U1489 ( .A(n1359), .B(KEYINPUT32), .ZN(n1361) );
  NAND2_X1 U1490 ( .A1(G223), .A2(n960), .ZN(n1360) );
  NAND2_X1 U1491 ( .A1(n1361), .A2(n1360), .ZN(n1362) );
  XNOR2_X1 U1492 ( .A(n1362), .B(KEYINPUT33), .ZN(n1363) );
  NAND2_X1 U1493 ( .A1(n1363), .A2(n1391), .ZN(n1364) );
  NOR2_X1 U1494 ( .A1(n1371), .A2(n1366), .ZN(n1367) );
  XNOR2_X1 U1495 ( .A(n1367), .B(KEYINPUT35), .ZN(n1369) );
  NAND2_X1 U1496 ( .A1(n1371), .A2(G190), .ZN(n1368) );
  NAND2_X1 U1497 ( .A1(n1369), .A2(n1368), .ZN(n1370) );
  NOR2_X1 U1498 ( .A1(n1381), .A2(n1370), .ZN(n1432) );
  INV_X1 U1499 ( .A(n1371), .ZN(n1374) );
  XOR2_X1 U1500 ( .A(n1373), .B(KEYINPUT34), .Z(n1376) );
  NAND2_X1 U1501 ( .A1(n1374), .A2(G169), .ZN(n1375) );
  NAND2_X1 U1502 ( .A1(n1376), .A2(n1375), .ZN(n1380) );
  NOR2_X1 U1503 ( .A1(n1380), .A2(n1458), .ZN(n1377) );
  NOR2_X1 U1504 ( .A1(n1378), .A2(n1377), .ZN(n1379) );
  NOR2_X1 U1505 ( .A1(n1432), .A2(n1379), .ZN(n1383) );
  NAND2_X1 U1506 ( .A1(n1381), .A2(n1380), .ZN(n1457) );
  INV_X1 U1507 ( .A(n1457), .ZN(n1427) );
  AND2_X1 U1508 ( .A1(n1427), .A2(n1458), .ZN(n1382) );
  NOR2_X1 U1509 ( .A1(n1383), .A2(n1382), .ZN(n1534) );
  XNOR2_X2 U1510 ( .A(n1385), .B(n1384), .ZN(n1557) );
  XNOR2_X1 U1511 ( .A(n1387), .B(n1386), .ZN(n1448) );
  NAND2_X1 U1512 ( .A1(G222), .A2(n960), .ZN(n1388) );
  XNOR2_X1 U1513 ( .A(n1388), .B(KEYINPUT36), .ZN(n1399) );
  NAND2_X1 U1514 ( .A1(n1389), .A2(G77), .ZN(n1390) );
  NAND2_X1 U1515 ( .A1(n1391), .A2(n1390), .ZN(n1397) );
  NAND2_X1 U1516 ( .A1(G226), .A2(n1392), .ZN(n1395) );
  NAND2_X1 U1517 ( .A1(G223), .A2(n1393), .ZN(n1394) );
  NAND2_X1 U1518 ( .A1(n1395), .A2(n1394), .ZN(n1396) );
  NOR2_X1 U1519 ( .A1(n1397), .A2(n1396), .ZN(n1398) );
  NAND2_X1 U1520 ( .A1(n1399), .A2(n1398), .ZN(n1419) );
  NAND2_X1 U1521 ( .A1(n1400), .A2(n1419), .ZN(n1414) );
  NAND2_X1 U1522 ( .A1(n1401), .A2(G58), .ZN(n1404) );
  NAND2_X1 U1523 ( .A1(n1402), .A2(n1894), .ZN(n1403) );
  NAND2_X1 U1524 ( .A1(n1404), .A2(n1403), .ZN(n1407) );
  AND2_X1 U1525 ( .A1(n1405), .A2(G150), .ZN(n1406) );
  NOR2_X1 U1526 ( .A1(n1407), .A2(n1406), .ZN(n1413) );
  NOR2_X1 U1527 ( .A1(n1408), .A2(n1894), .ZN(n1411) );
  NOR2_X1 U1528 ( .A1(n1409), .A2(n1895), .ZN(n1410) );
  NOR2_X1 U1529 ( .A1(n1411), .A2(n1410), .ZN(n1412) );
  NAND2_X1 U1530 ( .A1(n1413), .A2(n1412), .ZN(n1450) );
  NAND2_X1 U1531 ( .A1(n1414), .A2(n1450), .ZN(n1416) );
  NOR2_X1 U1532 ( .A1(G179), .A2(n1419), .ZN(n1415) );
  NOR2_X1 U1533 ( .A1(n1416), .A2(n1415), .ZN(n1453) );
  INV_X1 U1534 ( .A(n1450), .ZN(n1418) );
  NAND2_X1 U1535 ( .A1(G200), .A2(n1419), .ZN(n1417) );
  NAND2_X1 U1536 ( .A1(n1418), .A2(n1417), .ZN(n1422) );
  NOR2_X1 U1537 ( .A1(n1420), .A2(n1419), .ZN(n1421) );
  NOR2_X1 U1538 ( .A1(n1422), .A2(n1421), .ZN(n1423) );
  NOR2_X1 U1539 ( .A1(n1453), .A2(n1423), .ZN(n1424) );
  XOR2_X1 U1540 ( .A(KEYINPUT37), .B(n1424), .Z(n1451) );
  NAND2_X1 U1541 ( .A1(n1433), .A2(n1451), .ZN(n1425) );
  NOR2_X1 U1542 ( .A1(n1432), .A2(n1425), .ZN(n1429) );
  NAND2_X1 U1543 ( .A1(n1429), .A2(n1428), .ZN(n1869) );
  INV_X1 U1544 ( .A(n1869), .ZN(n1897) );
  NAND2_X1 U1545 ( .A1(G330), .A2(n1897), .ZN(n1431) );
  INV_X1 U1546 ( .A(n1430), .ZN(n1870) );
  INV_X1 U1547 ( .A(n1432), .ZN(n1438) );
  NAND2_X1 U1548 ( .A1(n1434), .A2(n1433), .ZN(n1435) );
  NAND2_X1 U1549 ( .A1(n1436), .A2(n1435), .ZN(n1437) );
  NAND2_X1 U1550 ( .A1(n1438), .A2(n1437), .ZN(n1439) );
  NAND2_X1 U1551 ( .A1(n1439), .A2(n1457), .ZN(n1440) );
  AND2_X1 U1552 ( .A1(n1440), .A2(n1451), .ZN(n1441) );
  NOR2_X1 U1553 ( .A1(n1453), .A2(n1441), .ZN(n1899) );
  INV_X1 U1554 ( .A(n1899), .ZN(n1444) );
  NOR2_X1 U1555 ( .A1(n1442), .A2(n1869), .ZN(n1443) );
  NOR2_X1 U1556 ( .A1(n1444), .A2(n1443), .ZN(n1867) );
  NAND2_X1 U1557 ( .A1(n1445), .A2(n1867), .ZN(n1446) );
  XNOR2_X1 U1558 ( .A(n1446), .B(KEYINPUT38), .ZN(n1561) );
  NOR2_X1 U1559 ( .A1(n1672), .A2(n1561), .ZN(n1447) );
  NAND2_X1 U1560 ( .A1(n1450), .A2(n1458), .ZN(n1452) );
  NAND2_X1 U1561 ( .A1(n1452), .A2(n1451), .ZN(n1455) );
  NAND2_X1 U1562 ( .A1(n1453), .A2(n1458), .ZN(n1454) );
  NAND2_X1 U1563 ( .A1(n1455), .A2(n1454), .ZN(n1507) );
  NOR2_X1 U1564 ( .A1(n1456), .A2(n1534), .ZN(n1460) );
  NOR2_X1 U1565 ( .A1(n1458), .A2(n1457), .ZN(n1459) );
  NOR2_X1 U1566 ( .A1(n1460), .A2(n1459), .ZN(n1868) );
  NOR2_X1 U1567 ( .A1(n1801), .A2(n1598), .ZN(n1462) );
  INV_X1 U1568 ( .A(n1534), .ZN(n1461) );
  NAND2_X1 U1569 ( .A1(n1462), .A2(n1461), .ZN(n1463) );
  NOR2_X1 U1570 ( .A1(n1870), .A2(n1463), .ZN(n1871) );
  NAND2_X1 U1571 ( .A1(G330), .A2(n1871), .ZN(n1464) );
  NAND2_X1 U1572 ( .A1(n1868), .A2(n1464), .ZN(n1465) );
  XOR2_X1 U1573 ( .A(n1507), .B(n1465), .Z(n1466) );
  NAND2_X1 U1574 ( .A1(n1467), .A2(n1466), .ZN(n1512) );
  NOR2_X1 U1575 ( .A1(G41), .A2(n1753), .ZN(n1502) );
  NAND2_X1 U1576 ( .A1(G132), .A2(n1775), .ZN(n1469) );
  NAND2_X1 U1577 ( .A1(G159), .A2(n1626), .ZN(n1468) );
  NAND2_X1 U1578 ( .A1(n1469), .A2(n1468), .ZN(n1470) );
  XNOR2_X1 U1579 ( .A(KEYINPUT44), .B(n1470), .ZN(n1483) );
  NAND2_X1 U1580 ( .A1(G125), .A2(n1782), .ZN(n1472) );
  NAND2_X1 U1581 ( .A1(G124), .A2(n1778), .ZN(n1471) );
  NAND2_X1 U1582 ( .A1(n1472), .A2(n1471), .ZN(n1474) );
  AND2_X1 U1583 ( .A1(n1786), .A2(G143), .ZN(n1473) );
  NOR2_X1 U1584 ( .A1(n1474), .A2(n1473), .ZN(n1481) );
  NAND2_X1 U1585 ( .A1(n1772), .A2(G128), .ZN(n1476) );
  NAND2_X1 U1586 ( .A1(G150), .A2(n1787), .ZN(n1475) );
  NAND2_X1 U1587 ( .A1(n1476), .A2(n1475), .ZN(n1479) );
  NAND2_X1 U1588 ( .A1(n1783), .A2(G137), .ZN(n1477) );
  XNOR2_X1 U1589 ( .A(KEYINPUT43), .B(n1477), .ZN(n1478) );
  NOR2_X1 U1590 ( .A1(n1479), .A2(n1478), .ZN(n1480) );
  NAND2_X1 U1591 ( .A1(n1481), .A2(n1480), .ZN(n1482) );
  NOR2_X1 U1592 ( .A1(n1483), .A2(n1482), .ZN(n1484) );
  NOR2_X1 U1593 ( .A1(G33), .A2(n1484), .ZN(n1500) );
  NOR2_X1 U1594 ( .A1(n1881), .A2(n1761), .ZN(n1607) );
  NAND2_X1 U1595 ( .A1(n1778), .A2(G283), .ZN(n1486) );
  NAND2_X1 U1596 ( .A1(n1782), .A2(G116), .ZN(n1485) );
  NAND2_X1 U1597 ( .A1(n1486), .A2(n1485), .ZN(n1487) );
  NOR2_X1 U1598 ( .A1(n1607), .A2(n1487), .ZN(n1494) );
  NAND2_X1 U1599 ( .A1(n1775), .A2(G97), .ZN(n1489) );
  NAND2_X1 U1600 ( .A1(n1783), .A2(G87), .ZN(n1488) );
  NAND2_X1 U1601 ( .A1(n1489), .A2(n1488), .ZN(n1492) );
  NAND2_X1 U1602 ( .A1(G107), .A2(n1772), .ZN(n1490) );
  XOR2_X1 U1603 ( .A(KEYINPUT42), .B(n1490), .Z(n1491) );
  NOR2_X1 U1604 ( .A1(n1492), .A2(n1491), .ZN(n1493) );
  NAND2_X1 U1605 ( .A1(n1494), .A2(n1493), .ZN(n1496) );
  NAND2_X1 U1606 ( .A1(G68), .A2(n1787), .ZN(n1705) );
  NAND2_X1 U1607 ( .A1(n1626), .A2(G58), .ZN(n1589) );
  NAND2_X1 U1608 ( .A1(n1705), .A2(n1589), .ZN(n1495) );
  NOR2_X1 U1609 ( .A1(n1496), .A2(n1495), .ZN(n1497) );
  NOR2_X1 U1610 ( .A1(n1498), .A2(n1497), .ZN(n1499) );
  NOR2_X1 U1611 ( .A1(n1500), .A2(n1499), .ZN(n1501) );
  NAND2_X1 U1612 ( .A1(n1502), .A2(n1501), .ZN(n1506) );
  INV_X1 U1613 ( .A(n1502), .ZN(n1504) );
  NOR2_X1 U1614 ( .A1(G50), .A2(n1747), .ZN(n1503) );
  NAND2_X1 U1615 ( .A1(n1504), .A2(n1503), .ZN(n1505) );
  NAND2_X1 U1616 ( .A1(n1506), .A2(n1505), .ZN(n1509) );
  NOR2_X1 U1617 ( .A1(n1654), .A2(n1507), .ZN(n1508) );
  NOR2_X1 U1618 ( .A1(n1509), .A2(n1508), .ZN(n1510) );
  NAND2_X1 U1619 ( .A1(n1510), .A2(n1620), .ZN(n1511) );
  INV_X1 U1620 ( .A(n1863), .ZN(n1515) );
  NOR2_X1 U1621 ( .A1(n1561), .A2(n1560), .ZN(n1513) );
  XNOR2_X1 U1622 ( .A(n1513), .B(n1557), .ZN(n1514) );
  NOR2_X1 U1623 ( .A1(n1515), .A2(n1514), .ZN(n1556) );
  NAND2_X1 U1624 ( .A1(n1654), .A2(n1753), .ZN(n1748) );
  NOR2_X1 U1625 ( .A1(G58), .A2(n1748), .ZN(n1516) );
  NOR2_X1 U1626 ( .A1(n1802), .A2(n1516), .ZN(n1533) );
  NAND2_X1 U1627 ( .A1(G125), .A2(n1778), .ZN(n1518) );
  NAND2_X1 U1628 ( .A1(G137), .A2(n1775), .ZN(n1517) );
  NAND2_X1 U1629 ( .A1(n1518), .A2(n1517), .ZN(n1523) );
  AND2_X1 U1630 ( .A1(n1786), .A2(G150), .ZN(n1519) );
  NOR2_X1 U1631 ( .A1(n1709), .A2(n1519), .ZN(n1521) );
  NAND2_X1 U1632 ( .A1(n1772), .A2(G132), .ZN(n1520) );
  NAND2_X1 U1633 ( .A1(n1521), .A2(n1520), .ZN(n1522) );
  NOR2_X1 U1634 ( .A1(n1523), .A2(n1522), .ZN(n1531) );
  NAND2_X1 U1635 ( .A1(G128), .A2(n1782), .ZN(n1525) );
  NAND2_X1 U1636 ( .A1(G50), .A2(n1626), .ZN(n1524) );
  NAND2_X1 U1637 ( .A1(n1525), .A2(n1524), .ZN(n1529) );
  NAND2_X1 U1638 ( .A1(n1783), .A2(G143), .ZN(n1527) );
  NAND2_X1 U1639 ( .A1(G159), .A2(n1787), .ZN(n1526) );
  NAND2_X1 U1640 ( .A1(n1527), .A2(n1526), .ZN(n1528) );
  NOR2_X1 U1641 ( .A1(n1529), .A2(n1528), .ZN(n1530) );
  NAND2_X1 U1642 ( .A1(n1531), .A2(n1530), .ZN(n1532) );
  NAND2_X1 U1643 ( .A1(n1533), .A2(n1532), .ZN(n1554) );
  NAND2_X1 U1644 ( .A1(n1747), .A2(n1534), .ZN(n1552) );
  NAND2_X1 U1645 ( .A1(G107), .A2(n1775), .ZN(n1535) );
  NAND2_X1 U1646 ( .A1(n1536), .A2(n1535), .ZN(n1545) );
  NAND2_X1 U1647 ( .A1(n1772), .A2(G116), .ZN(n1537) );
  XNOR2_X1 U1648 ( .A(KEYINPUT47), .B(n1537), .ZN(n1538) );
  NOR2_X1 U1649 ( .A1(n1624), .A2(n1538), .ZN(n1543) );
  AND2_X1 U1650 ( .A1(G283), .A2(n1782), .ZN(n1541) );
  NAND2_X1 U1651 ( .A1(G68), .A2(n1626), .ZN(n1774) );
  NAND2_X1 U1652 ( .A1(n1774), .A2(n1539), .ZN(n1540) );
  NOR2_X1 U1653 ( .A1(n1541), .A2(n1540), .ZN(n1542) );
  NAND2_X1 U1654 ( .A1(n1543), .A2(n1542), .ZN(n1544) );
  NOR2_X1 U1655 ( .A1(n1545), .A2(n1544), .ZN(n1550) );
  NAND2_X1 U1656 ( .A1(n1778), .A2(G294), .ZN(n1547) );
  NAND2_X1 U1657 ( .A1(n1783), .A2(G97), .ZN(n1546) );
  NAND2_X1 U1658 ( .A1(n1547), .A2(n1546), .ZN(n1548) );
  XOR2_X1 U1659 ( .A(KEYINPUT48), .B(n1548), .Z(n1549) );
  NAND2_X1 U1660 ( .A1(n1550), .A2(n1549), .ZN(n1551) );
  NAND2_X1 U1661 ( .A1(n1552), .A2(n1551), .ZN(n1553) );
  NOR2_X1 U1662 ( .A1(n1554), .A2(n1553), .ZN(n1555) );
  NOR2_X1 U1663 ( .A1(n1556), .A2(n1555), .ZN(n1559) );
  NAND2_X1 U1664 ( .A1(n1672), .A2(n1557), .ZN(n1558) );
  NAND2_X1 U1665 ( .A1(n1559), .A2(n1558), .ZN(G378) );
  NAND2_X1 U1666 ( .A1(n961), .A2(n1863), .ZN(n1604) );
  AND2_X1 U1667 ( .A1(n1563), .A2(n1672), .ZN(n1602) );
  NAND2_X1 U1668 ( .A1(G77), .A2(n1626), .ZN(n1711) );
  NAND2_X1 U1669 ( .A1(G97), .A2(n1786), .ZN(n1564) );
  NAND2_X1 U1670 ( .A1(n1711), .A2(n1564), .ZN(n1576) );
  NAND2_X1 U1671 ( .A1(n1782), .A2(G294), .ZN(n1566) );
  NAND2_X1 U1672 ( .A1(n1772), .A2(G283), .ZN(n1565) );
  NAND2_X1 U1673 ( .A1(n1566), .A2(n1565), .ZN(n1567) );
  NOR2_X1 U1674 ( .A1(n1624), .A2(n1567), .ZN(n1574) );
  NAND2_X1 U1675 ( .A1(G87), .A2(n1787), .ZN(n1613) );
  NAND2_X1 U1676 ( .A1(G116), .A2(n1775), .ZN(n1568) );
  NAND2_X1 U1677 ( .A1(n1613), .A2(n1568), .ZN(n1572) );
  NAND2_X1 U1678 ( .A1(n1778), .A2(G303), .ZN(n1570) );
  NAND2_X1 U1679 ( .A1(n1783), .A2(G107), .ZN(n1569) );
  NAND2_X1 U1680 ( .A1(n1570), .A2(n1569), .ZN(n1571) );
  NOR2_X1 U1681 ( .A1(n1572), .A2(n1571), .ZN(n1573) );
  NAND2_X1 U1682 ( .A1(n1574), .A2(n1573), .ZN(n1575) );
  NOR2_X1 U1683 ( .A1(n1576), .A2(n1575), .ZN(n1593) );
  NAND2_X1 U1684 ( .A1(G137), .A2(n1772), .ZN(n1578) );
  NAND2_X1 U1685 ( .A1(G132), .A2(n1782), .ZN(n1577) );
  NAND2_X1 U1686 ( .A1(n1578), .A2(n1577), .ZN(n1579) );
  NOR2_X1 U1687 ( .A1(n1709), .A2(n1579), .ZN(n1587) );
  NAND2_X1 U1688 ( .A1(G128), .A2(n1778), .ZN(n1581) );
  NAND2_X1 U1689 ( .A1(G150), .A2(n1783), .ZN(n1580) );
  NAND2_X1 U1690 ( .A1(n1581), .A2(n1580), .ZN(n1585) );
  NAND2_X1 U1691 ( .A1(n1775), .A2(G143), .ZN(n1583) );
  NAND2_X1 U1692 ( .A1(G50), .A2(n1787), .ZN(n1582) );
  NAND2_X1 U1693 ( .A1(n1583), .A2(n1582), .ZN(n1584) );
  NOR2_X1 U1694 ( .A1(n1585), .A2(n1584), .ZN(n1586) );
  NAND2_X1 U1695 ( .A1(n1587), .A2(n1586), .ZN(n1591) );
  NAND2_X1 U1696 ( .A1(n1786), .A2(G159), .ZN(n1588) );
  NAND2_X1 U1697 ( .A1(n1589), .A2(n1588), .ZN(n1590) );
  NOR2_X1 U1698 ( .A1(n1591), .A2(n1590), .ZN(n1592) );
  NOR2_X1 U1699 ( .A1(n1593), .A2(n1592), .ZN(n1594) );
  NAND2_X1 U1700 ( .A1(n1620), .A2(n1594), .ZN(n1596) );
  NOR2_X1 U1701 ( .A1(G68), .A2(n1748), .ZN(n1595) );
  NOR2_X1 U1702 ( .A1(n1596), .A2(n1595), .ZN(n1597) );
  XNOR2_X1 U1703 ( .A(n1597), .B(KEYINPUT45), .ZN(n1600) );
  AND2_X1 U1704 ( .A1(n1747), .A2(n1598), .ZN(n1599) );
  NOR2_X1 U1705 ( .A1(n1600), .A2(n1599), .ZN(n1601) );
  NOR2_X1 U1706 ( .A1(n1602), .A2(n1601), .ZN(n1603) );
  NAND2_X1 U1707 ( .A1(n1604), .A2(n1603), .ZN(G381) );
  NAND2_X1 U1708 ( .A1(G150), .A2(n1778), .ZN(n1606) );
  NAND2_X1 U1709 ( .A1(G58), .A2(n1775), .ZN(n1605) );
  NAND2_X1 U1710 ( .A1(n1606), .A2(n1605), .ZN(n1611) );
  NOR2_X1 U1711 ( .A1(n1607), .A2(n1709), .ZN(n1609) );
  NAND2_X1 U1712 ( .A1(n1782), .A2(G159), .ZN(n1608) );
  NAND2_X1 U1713 ( .A1(n1609), .A2(n1608), .ZN(n1610) );
  NOR2_X1 U1714 ( .A1(n1611), .A2(n1610), .ZN(n1618) );
  NAND2_X1 U1715 ( .A1(G97), .A2(n1626), .ZN(n1734) );
  NAND2_X1 U1716 ( .A1(n1772), .A2(G50), .ZN(n1612) );
  NAND2_X1 U1717 ( .A1(n1734), .A2(n1612), .ZN(n1616) );
  NAND2_X1 U1718 ( .A1(G68), .A2(n1783), .ZN(n1614) );
  NAND2_X1 U1719 ( .A1(n1614), .A2(n1613), .ZN(n1615) );
  NOR2_X1 U1720 ( .A1(n1616), .A2(n1615), .ZN(n1617) );
  NAND2_X1 U1721 ( .A1(n1618), .A2(n1617), .ZN(n1619) );
  NAND2_X1 U1722 ( .A1(n1620), .A2(n1619), .ZN(n1641) );
  NAND2_X1 U1723 ( .A1(G322), .A2(n1782), .ZN(n1622) );
  NAND2_X1 U1724 ( .A1(n1786), .A2(G294), .ZN(n1621) );
  NAND2_X1 U1725 ( .A1(n1622), .A2(n1621), .ZN(n1623) );
  XNOR2_X1 U1726 ( .A(KEYINPUT26), .B(n1623), .ZN(n1639) );
  INV_X1 U1727 ( .A(n1624), .ZN(n1727) );
  NAND2_X1 U1728 ( .A1(n1778), .A2(G326), .ZN(n1625) );
  NAND2_X1 U1729 ( .A1(n1727), .A2(n1625), .ZN(n1629) );
  NAND2_X1 U1730 ( .A1(G116), .A2(n1626), .ZN(n1627) );
  XNOR2_X1 U1731 ( .A(KEYINPUT25), .B(n1627), .ZN(n1628) );
  NOR2_X1 U1732 ( .A1(n1629), .A2(n1628), .ZN(n1637) );
  NAND2_X1 U1733 ( .A1(n1775), .A2(G311), .ZN(n1631) );
  NAND2_X1 U1734 ( .A1(G283), .A2(n1787), .ZN(n1630) );
  NAND2_X1 U1735 ( .A1(n1631), .A2(n1630), .ZN(n1635) );
  NAND2_X1 U1736 ( .A1(n1772), .A2(G317), .ZN(n1633) );
  NAND2_X1 U1737 ( .A1(n1783), .A2(G303), .ZN(n1632) );
  NAND2_X1 U1738 ( .A1(n1633), .A2(n1632), .ZN(n1634) );
  NOR2_X1 U1739 ( .A1(n1635), .A2(n1634), .ZN(n1636) );
  NAND2_X1 U1740 ( .A1(n1637), .A2(n1636), .ZN(n1638) );
  NOR2_X1 U1741 ( .A1(n1639), .A2(n1638), .ZN(n1640) );
  NOR2_X1 U1742 ( .A1(n1641), .A2(n1640), .ZN(n1661) );
  NAND2_X1 U1743 ( .A1(n1762), .A2(n1828), .ZN(n1658) );
  NOR2_X1 U1744 ( .A1(G116), .A2(n1642), .ZN(n1858) );
  NAND2_X1 U1745 ( .A1(G68), .A2(G77), .ZN(n1643) );
  NAND2_X1 U1746 ( .A1(n1858), .A2(n1643), .ZN(n1645) );
  NAND2_X1 U1747 ( .A1(G58), .A2(n1894), .ZN(n1644) );
  NOR2_X1 U1748 ( .A1(n1645), .A2(n1644), .ZN(n1646) );
  NOR2_X1 U1749 ( .A1(G45), .A2(n1646), .ZN(n1647) );
  XOR2_X1 U1750 ( .A(KEYINPUT23), .B(n1647), .Z(n1652) );
  XNOR2_X1 U1751 ( .A(G244), .B(G232), .ZN(n1648) );
  XNOR2_X1 U1752 ( .A(n1648), .B(G226), .ZN(n1649) );
  XNOR2_X1 U1753 ( .A(G238), .B(n1649), .ZN(n1900) );
  NOR2_X1 U1754 ( .A1(n1900), .A2(n1650), .ZN(n1651) );
  NOR2_X1 U1755 ( .A1(n1652), .A2(n1651), .ZN(n1653) );
  NOR2_X1 U1756 ( .A1(n1700), .A2(n1653), .ZN(n1656) );
  NOR2_X1 U1757 ( .A1(n1858), .A2(n1654), .ZN(n1655) );
  NOR2_X1 U1758 ( .A1(n1656), .A2(n1655), .ZN(n1657) );
  NAND2_X1 U1759 ( .A1(n1658), .A2(n1657), .ZN(n1659) );
  NAND2_X1 U1760 ( .A1(n1659), .A2(n1697), .ZN(n1660) );
  NAND2_X1 U1761 ( .A1(n1661), .A2(n1660), .ZN(n1664) );
  NOR2_X1 U1762 ( .A1(n1662), .A2(n1741), .ZN(n1663) );
  NOR2_X1 U1763 ( .A1(n1664), .A2(n1663), .ZN(n1667) );
  NAND2_X1 U1764 ( .A1(n1863), .A2(n1857), .ZN(n1665) );
  NOR2_X1 U1765 ( .A1(n1669), .A2(n1665), .ZN(n1666) );
  NOR2_X1 U1766 ( .A1(n1667), .A2(n1666), .ZN(n1671) );
  NAND2_X1 U1767 ( .A1(n1669), .A2(n1668), .ZN(n1670) );
  NAND2_X1 U1768 ( .A1(n1671), .A2(n1670), .ZN(G393) );
  NOR2_X1 U1769 ( .A1(n1673), .A2(n1672), .ZN(n1674) );
  NAND2_X1 U1770 ( .A1(n1675), .A2(n1674), .ZN(n1676) );
  NAND2_X1 U1771 ( .A1(n1676), .A2(n1802), .ZN(n1695) );
  NOR2_X1 U1772 ( .A1(n1677), .A2(n1855), .ZN(n1693) );
  NAND2_X1 U1773 ( .A1(n1679), .A2(n1678), .ZN(n1680) );
  XOR2_X1 U1774 ( .A(n963), .B(n1680), .Z(n1681) );
  NAND2_X1 U1775 ( .A1(n1681), .A2(n1292), .ZN(n1684) );
  NAND2_X1 U1776 ( .A1(n1687), .A2(n1682), .ZN(n1683) );
  NAND2_X1 U1777 ( .A1(n1684), .A2(n1683), .ZN(n1685) );
  XNOR2_X1 U1778 ( .A(n1685), .B(KEYINPUT53), .ZN(n1691) );
  NAND2_X1 U1779 ( .A1(n1687), .A2(n1686), .ZN(n1688) );
  NOR2_X1 U1780 ( .A1(n1689), .A2(n1688), .ZN(n1690) );
  NOR2_X1 U1781 ( .A1(n1691), .A2(n1690), .ZN(n1692) );
  XNOR2_X1 U1782 ( .A(n1693), .B(n1692), .ZN(n1694) );
  NOR2_X1 U1783 ( .A1(n1695), .A2(n1694), .ZN(n1745) );
  NAND2_X1 U1784 ( .A1(G87), .A2(n1828), .ZN(n1696) );
  NAND2_X1 U1785 ( .A1(n1697), .A2(n1696), .ZN(n1702) );
  XOR2_X1 U1786 ( .A(G264), .B(G270), .Z(n1699) );
  XNOR2_X1 U1787 ( .A(G250), .B(G257), .ZN(n1698) );
  XNOR2_X1 U1788 ( .A(n1699), .B(n1698), .ZN(n1901) );
  NOR2_X1 U1789 ( .A1(n1901), .A2(n1700), .ZN(n1701) );
  NOR2_X1 U1790 ( .A1(n1702), .A2(n1701), .ZN(n1703) );
  NOR2_X1 U1791 ( .A1(n1802), .A2(n1703), .ZN(n1740) );
  NAND2_X1 U1792 ( .A1(n1786), .A2(G58), .ZN(n1704) );
  NAND2_X1 U1793 ( .A1(n1705), .A2(n1704), .ZN(n1719) );
  NAND2_X1 U1794 ( .A1(G150), .A2(n1772), .ZN(n1707) );
  NAND2_X1 U1795 ( .A1(G143), .A2(n1782), .ZN(n1706) );
  NAND2_X1 U1796 ( .A1(n1707), .A2(n1706), .ZN(n1708) );
  NOR2_X1 U1797 ( .A1(n1709), .A2(n1708), .ZN(n1717) );
  NAND2_X1 U1798 ( .A1(n1775), .A2(G159), .ZN(n1710) );
  NAND2_X1 U1799 ( .A1(n1711), .A2(n1710), .ZN(n1715) );
  NAND2_X1 U1800 ( .A1(G137), .A2(n1778), .ZN(n1713) );
  NAND2_X1 U1801 ( .A1(G50), .A2(n1783), .ZN(n1712) );
  NAND2_X1 U1802 ( .A1(n1713), .A2(n1712), .ZN(n1714) );
  NOR2_X1 U1803 ( .A1(n1715), .A2(n1714), .ZN(n1716) );
  NAND2_X1 U1804 ( .A1(n1717), .A2(n1716), .ZN(n1718) );
  NOR2_X1 U1805 ( .A1(n1719), .A2(n1718), .ZN(n1738) );
  NAND2_X1 U1806 ( .A1(G303), .A2(n1772), .ZN(n1721) );
  NAND2_X1 U1807 ( .A1(G107), .A2(n1787), .ZN(n1720) );
  NAND2_X1 U1808 ( .A1(n1721), .A2(n1720), .ZN(n1723) );
  NOR2_X1 U1809 ( .A1(n1889), .A2(n1761), .ZN(n1722) );
  NOR2_X1 U1810 ( .A1(n1723), .A2(n1722), .ZN(n1732) );
  NAND2_X1 U1811 ( .A1(G294), .A2(n1775), .ZN(n1725) );
  NAND2_X1 U1812 ( .A1(n1778), .A2(G317), .ZN(n1724) );
  NAND2_X1 U1813 ( .A1(n1725), .A2(n1724), .ZN(n1730) );
  NAND2_X1 U1814 ( .A1(G311), .A2(n1782), .ZN(n1726) );
  XNOR2_X1 U1815 ( .A(n1726), .B(KEYINPUT54), .ZN(n1728) );
  NAND2_X1 U1816 ( .A1(n1728), .A2(n1727), .ZN(n1729) );
  NOR2_X1 U1817 ( .A1(n1730), .A2(n1729), .ZN(n1731) );
  NAND2_X1 U1818 ( .A1(n1732), .A2(n1731), .ZN(n1736) );
  NAND2_X1 U1819 ( .A1(G283), .A2(n1783), .ZN(n1733) );
  NAND2_X1 U1820 ( .A1(n1734), .A2(n1733), .ZN(n1735) );
  NOR2_X1 U1821 ( .A1(n1736), .A2(n1735), .ZN(n1737) );
  NOR2_X1 U1822 ( .A1(n1738), .A2(n1737), .ZN(n1739) );
  NAND2_X1 U1823 ( .A1(n1740), .A2(n1739), .ZN(n1743) );
  NOR2_X1 U1824 ( .A1(n1741), .A2(n963), .ZN(n1742) );
  NOR2_X1 U1825 ( .A1(n1743), .A2(n1742), .ZN(n1744) );
  NAND2_X1 U1826 ( .A1(n1801), .A2(n1747), .ZN(n1800) );
  NOR2_X1 U1827 ( .A1(G77), .A2(n1748), .ZN(n1749) );
  NOR2_X1 U1828 ( .A1(n1802), .A2(n1749), .ZN(n1771) );
  NAND2_X1 U1829 ( .A1(G311), .A2(n1778), .ZN(n1751) );
  NAND2_X1 U1830 ( .A1(n1775), .A2(G283), .ZN(n1750) );
  NAND2_X1 U1831 ( .A1(n1751), .A2(n1750), .ZN(n1752) );
  NOR2_X1 U1832 ( .A1(n1753), .A2(n1752), .ZN(n1755) );
  NAND2_X1 U1833 ( .A1(n1755), .A2(n1754), .ZN(n1758) );
  NAND2_X1 U1834 ( .A1(G116), .A2(n1783), .ZN(n1756) );
  XNOR2_X1 U1835 ( .A(KEYINPUT21), .B(n1756), .ZN(n1757) );
  NOR2_X1 U1836 ( .A1(n1758), .A2(n1757), .ZN(n1769) );
  NAND2_X1 U1837 ( .A1(n1772), .A2(G294), .ZN(n1760) );
  NAND2_X1 U1838 ( .A1(n1782), .A2(G303), .ZN(n1759) );
  NAND2_X1 U1839 ( .A1(n1760), .A2(n1759), .ZN(n1764) );
  NOR2_X1 U1840 ( .A1(n1762), .A2(n1761), .ZN(n1763) );
  NOR2_X1 U1841 ( .A1(n1764), .A2(n1763), .ZN(n1765) );
  NAND2_X1 U1842 ( .A1(G33), .A2(n1765), .ZN(n1766) );
  NOR2_X1 U1843 ( .A1(n1767), .A2(n1766), .ZN(n1768) );
  NAND2_X1 U1844 ( .A1(n1769), .A2(n1768), .ZN(n1770) );
  NAND2_X1 U1845 ( .A1(n1771), .A2(n1770), .ZN(n1798) );
  NAND2_X1 U1846 ( .A1(n1772), .A2(G143), .ZN(n1773) );
  NAND2_X1 U1847 ( .A1(n1774), .A2(n1773), .ZN(n1796) );
  NAND2_X1 U1848 ( .A1(n1775), .A2(G150), .ZN(n1776) );
  NAND2_X1 U1849 ( .A1(n1777), .A2(n1776), .ZN(n1781) );
  NAND2_X1 U1850 ( .A1(G132), .A2(n1778), .ZN(n1779) );
  XNOR2_X1 U1851 ( .A(KEYINPUT19), .B(n1779), .ZN(n1780) );
  NOR2_X1 U1852 ( .A1(n1781), .A2(n1780), .ZN(n1794) );
  NAND2_X1 U1853 ( .A1(G137), .A2(n1782), .ZN(n1785) );
  NAND2_X1 U1854 ( .A1(G159), .A2(n1783), .ZN(n1784) );
  NAND2_X1 U1855 ( .A1(n1785), .A2(n1784), .ZN(n1791) );
  NAND2_X1 U1856 ( .A1(n1786), .A2(G50), .ZN(n1789) );
  NAND2_X1 U1857 ( .A1(G58), .A2(n1787), .ZN(n1788) );
  NAND2_X1 U1858 ( .A1(n1789), .A2(n1788), .ZN(n1790) );
  NOR2_X1 U1859 ( .A1(n1791), .A2(n1790), .ZN(n1792) );
  XNOR2_X1 U1860 ( .A(n1792), .B(KEYINPUT20), .ZN(n1793) );
  NAND2_X1 U1861 ( .A1(n1794), .A2(n1793), .ZN(n1795) );
  NOR2_X1 U1862 ( .A1(n1796), .A2(n1795), .ZN(n1797) );
  NOR2_X1 U1863 ( .A1(n1798), .A2(n1797), .ZN(n1799) );
  NAND2_X1 U1864 ( .A1(n1800), .A2(n1799), .ZN(n1805) );
  XOR2_X1 U1865 ( .A(n1801), .B(n1857), .Z(n1803) );
  NAND2_X1 U1866 ( .A1(n1803), .A2(n1802), .ZN(n1804) );
  NAND2_X1 U1867 ( .A1(n1805), .A2(n1804), .ZN(G384) );
  NOR2_X1 U1868 ( .A1(G381), .A2(G390), .ZN(n1807) );
  NOR2_X1 U1869 ( .A1(G393), .A2(G396), .ZN(n1806) );
  NAND2_X1 U1870 ( .A1(n1807), .A2(n1806), .ZN(n1808) );
  NOR2_X1 U1871 ( .A1(n1811), .A2(n1808), .ZN(n1810) );
  NOR2_X1 U1872 ( .A1(G387), .A2(G384), .ZN(n1809) );
  NAND2_X1 U1873 ( .A1(n1810), .A2(n1809), .ZN(G407) );
  INV_X1 U1874 ( .A(G213), .ZN(n1815) );
  NOR2_X1 U1875 ( .A1(G343), .A2(n1811), .ZN(n1812) );
  NOR2_X1 U1876 ( .A1(n1815), .A2(n1812), .ZN(n1813) );
  NAND2_X1 U1877 ( .A1(n1813), .A2(G407), .ZN(G409) );
  NOR2_X1 U1878 ( .A1(G343), .A2(n1815), .ZN(n1816) );
  NOR2_X1 U1879 ( .A1(n1904), .A2(n1816), .ZN(n1819) );
  NAND2_X1 U1880 ( .A1(n1816), .A2(G2897), .ZN(n1817) );
  XNOR2_X1 U1881 ( .A(n1817), .B(KEYINPUT63), .ZN(n1818) );
  NOR2_X2 U1882 ( .A1(n1819), .A2(n1818), .ZN(n1825) );
  XNOR2_X1 U1883 ( .A(n1825), .B(n1905), .ZN(G405) );
  NOR2_X1 U1884 ( .A1(n1827), .A2(n1826), .ZN(n1891) );
  NAND2_X1 U1885 ( .A1(n1891), .A2(n1862), .ZN(n1832) );
  NOR2_X1 U1886 ( .A1(G257), .A2(G264), .ZN(n1829) );
  NOR2_X1 U1887 ( .A1(n1829), .A2(n1828), .ZN(n1830) );
  NAND2_X1 U1888 ( .A1(n1830), .A2(G250), .ZN(n1831) );
  NAND2_X1 U1889 ( .A1(n1832), .A2(n1831), .ZN(n1852) );
  NAND2_X1 U1890 ( .A1(G87), .A2(G250), .ZN(n1834) );
  NAND2_X1 U1891 ( .A1(G270), .A2(G116), .ZN(n1833) );
  NAND2_X1 U1892 ( .A1(n1834), .A2(n1833), .ZN(n1837) );
  NAND2_X1 U1893 ( .A1(G107), .A2(G264), .ZN(n1835) );
  XOR2_X1 U1894 ( .A(KEYINPUT50), .B(n1835), .Z(n1836) );
  NOR2_X1 U1895 ( .A1(n1837), .A2(n1836), .ZN(n1839) );
  NAND2_X1 U1896 ( .A1(G97), .A2(G257), .ZN(n1838) );
  NAND2_X1 U1897 ( .A1(n1839), .A2(n1838), .ZN(n1848) );
  NAND2_X1 U1898 ( .A1(G226), .A2(G50), .ZN(n1841) );
  NAND2_X1 U1899 ( .A1(G232), .A2(G58), .ZN(n1840) );
  NAND2_X1 U1900 ( .A1(n1841), .A2(n1840), .ZN(n1845) );
  NAND2_X1 U1901 ( .A1(G77), .A2(G244), .ZN(n1843) );
  NAND2_X1 U1902 ( .A1(G68), .A2(G238), .ZN(n1842) );
  NAND2_X1 U1903 ( .A1(n1843), .A2(n1842), .ZN(n1844) );
  NOR2_X1 U1904 ( .A1(n1845), .A2(n1844), .ZN(n1846) );
  XNOR2_X1 U1905 ( .A(KEYINPUT49), .B(n1846), .ZN(n1847) );
  NOR2_X1 U1906 ( .A1(n1848), .A2(n1847), .ZN(n1849) );
  NOR2_X1 U1907 ( .A1(n1850), .A2(n1849), .ZN(n1851) );
  NOR2_X1 U1908 ( .A1(n1852), .A2(n1851), .ZN(G361) );
  AND2_X1 U1909 ( .A1(n1853), .A2(n1897), .ZN(G372) );
  INV_X1 U1910 ( .A(n1854), .ZN(n1856) );
  NAND2_X1 U1911 ( .A1(n1856), .A2(n1855), .ZN(G399) );
  NOR2_X1 U1912 ( .A1(G1), .A2(n1857), .ZN(n1861) );
  NAND2_X1 U1913 ( .A1(G1), .A2(n1858), .ZN(n1859) );
  NOR2_X1 U1914 ( .A1(n1863), .A2(n1859), .ZN(n1860) );
  NOR2_X1 U1915 ( .A1(n1861), .A2(n1860), .ZN(n1865) );
  NAND2_X1 U1916 ( .A1(n1863), .A2(n1862), .ZN(n1864) );
  NAND2_X1 U1917 ( .A1(n1865), .A2(n1864), .ZN(G364) );
  NAND2_X1 U1918 ( .A1(n1866), .A2(G1), .ZN(n1879) );
  INV_X1 U1919 ( .A(n1891), .ZN(n1877) );
  XOR2_X1 U1920 ( .A(n1868), .B(n1867), .Z(n1875) );
  NOR2_X1 U1921 ( .A1(n1870), .A2(n1869), .ZN(n1872) );
  XOR2_X1 U1922 ( .A(n1872), .B(n1871), .Z(n1873) );
  NAND2_X1 U1923 ( .A1(n1873), .A2(G330), .ZN(n1874) );
  XNOR2_X1 U1924 ( .A(n1875), .B(n1874), .ZN(n1876) );
  NAND2_X1 U1925 ( .A1(n1877), .A2(n1876), .ZN(n1878) );
  NAND2_X1 U1926 ( .A1(n1879), .A2(n1878), .ZN(n1887) );
  INV_X1 U1927 ( .A(n1879), .ZN(n1885) );
  NAND2_X1 U1928 ( .A1(G58), .A2(G50), .ZN(n1880) );
  XNOR2_X1 U1929 ( .A(n1880), .B(G68), .ZN(n1883) );
  NAND2_X1 U1930 ( .A1(n1881), .A2(G50), .ZN(n1882) );
  NAND2_X1 U1931 ( .A1(n1883), .A2(n1882), .ZN(n1884) );
  NAND2_X1 U1932 ( .A1(n1885), .A2(n1884), .ZN(n1886) );
  NAND2_X1 U1933 ( .A1(n1887), .A2(n1886), .ZN(n1893) );
  NOR2_X1 U1934 ( .A1(n1889), .A2(n1888), .ZN(n1890) );
  NAND2_X1 U1935 ( .A1(n1891), .A2(n1890), .ZN(n1892) );
  NAND2_X1 U1936 ( .A1(n1893), .A2(n1892), .ZN(G367) );
  NAND2_X1 U1937 ( .A1(n1895), .A2(n1894), .ZN(n1896) );
  NOR2_X1 U1938 ( .A1(G77), .A2(n1896), .ZN(G353) );
  NAND2_X1 U1939 ( .A1(n1897), .A2(n1286), .ZN(n1898) );
  NAND2_X1 U1940 ( .A1(n1899), .A2(n1898), .ZN(G369) );
  XOR2_X1 U1941 ( .A(n1901), .B(n1900), .Z(G358) );
  XOR2_X1 U1942 ( .A(n1903), .B(n1902), .Z(G351) );
  XNOR2_X1 U1943 ( .A(n1905), .B(n1904), .ZN(G402) );
endmodule

