//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT85), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n202), .A2(KEYINPUT85), .ZN(new_n205));
  OAI21_X1  g004(.A(G36gat), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(new_n202), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT84), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(KEYINPUT14), .A3(new_n210), .ZN(new_n211));
  OR2_X1    g010(.A1(new_n210), .A2(KEYINPUT14), .ZN(new_n212));
  NOR2_X1   g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(G43gat), .A2(G50gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n206), .A2(new_n211), .A3(new_n212), .A4(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n215), .B1(new_n214), .B2(new_n216), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n216), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n221), .A2(new_n213), .A3(KEYINPUT15), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT85), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G29gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n208), .B1(new_n203), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n219), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n226), .A2(new_n227), .A3(new_n211), .A4(new_n212), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n220), .A2(new_n228), .A3(KEYINPUT17), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT86), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n220), .A2(new_n228), .A3(KEYINPUT86), .A4(KEYINPUT17), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(G1gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT16), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n237), .B1(G1gat), .B2(new_n234), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G8gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n220), .A2(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n233), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n239), .ZN(new_n245));
  INV_X1    g044(.A(new_n240), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n243), .A2(new_n244), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT87), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(G113gat), .B(G141gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT11), .ZN(new_n253));
  INV_X1    g052(.A(G169gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G197gat), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n256), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT12), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT12), .B1(new_n257), .B2(new_n258), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n239), .B(new_n240), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n244), .B(KEYINPUT13), .Z(new_n264));
  AOI22_X1  g063(.A1(new_n249), .A2(new_n250), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n247), .B1(new_n233), .B2(new_n242), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT18), .A3(new_n244), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n265), .B(new_n267), .C1(new_n251), .C2(new_n261), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT88), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n269), .A2(new_n270), .A3(KEYINPUT88), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT0), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G57gat), .ZN(new_n279));
  INV_X1    g078(.A(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  INV_X1    g081(.A(G120gat), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT1), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n284), .B1(new_n282), .B2(new_n283), .ZN(new_n285));
  XOR2_X1   g084(.A(G127gat), .B(G134gat), .Z(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n286), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT67), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G155gat), .B(G162gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(G141gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G148gat), .ZN(new_n297));
  INV_X1    g096(.A(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(G141gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n301));
  INV_X1    g100(.A(G155gat), .ZN(new_n302));
  INV_X1    g101(.A(G162gat), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT2), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n295), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n294), .A2(KEYINPUT77), .ZN(new_n308));
  OR3_X1    g107(.A1(new_n296), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(KEYINPUT76), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n294), .A2(KEYINPUT77), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n308), .A2(new_n311), .A3(new_n304), .A4(new_n312), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n293), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n307), .A2(new_n313), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT4), .B1(new_n317), .B2(new_n289), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT5), .ZN(new_n320));
  NAND2_X1  g119(.A1(G225gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n287), .A2(new_n288), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n325), .B1(new_n317), .B2(KEYINPUT3), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n322), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n319), .A2(new_n320), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n324), .A2(new_n326), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n293), .A2(new_n314), .A3(KEYINPUT4), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n315), .B1(new_n317), .B2(new_n289), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n321), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT78), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n327), .A2(new_n334), .A3(new_n331), .A4(new_n330), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n317), .B(new_n325), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT5), .B1(new_n337), .B2(new_n321), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n281), .B(new_n328), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n281), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n338), .B1(new_n333), .B2(new_n335), .ZN(new_n341));
  INV_X1    g140(.A(new_n328), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n340), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT6), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT82), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT82), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n339), .A2(new_n343), .A3(new_n347), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n328), .B1(new_n336), .B2(new_n338), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n350), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n254), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT23), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n254), .A2(new_n353), .A3(KEYINPUT23), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n356), .B(new_n357), .C1(new_n254), .C2(new_n353), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(G183gat), .A2(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT64), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n361), .B1(new_n363), .B2(KEYINPUT24), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(KEYINPUT24), .B2(new_n363), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n360), .A2(KEYINPUT65), .A3(new_n365), .ZN(new_n369));
  AND3_X1   g168(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  AOI211_X1 g170(.A(new_n361), .B(new_n370), .C1(new_n371), .C2(new_n362), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n359), .B1(new_n372), .B2(new_n358), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n354), .A2(KEYINPUT26), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n354), .A2(KEYINPUT26), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n375), .B(new_n376), .C1(new_n254), .C2(new_n353), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT27), .B(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379));
  INV_X1    g178(.A(G190gat), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n378), .A2(KEYINPUT66), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n380), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n377), .A2(new_n362), .A3(new_n381), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n293), .ZN(new_n387));
  INV_X1    g186(.A(new_n293), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n374), .A3(new_n385), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n387), .A2(G227gat), .A3(G233gat), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT32), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT33), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(G15gat), .B(G43gat), .Z(new_n394));
  XNOR2_X1  g193(.A(G71gat), .B(G99gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G227gat), .A2(G233gat), .ZN(new_n398));
  INV_X1    g197(.A(new_n389), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n388), .B1(new_n374), .B2(new_n385), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT34), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g202(.A(KEYINPUT34), .B(new_n398), .C1(new_n399), .C2(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n396), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n390), .B(KEYINPUT32), .C1(new_n392), .C2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n397), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT69), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n397), .A2(new_n405), .A3(KEYINPUT69), .A4(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT70), .B(G197gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(G204gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT71), .ZN(new_n415));
  AOI22_X1  g214(.A1(new_n415), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(new_n415), .B2(KEYINPUT22), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  XOR2_X1   g217(.A(G211gat), .B(G218gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT29), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n314), .B1(new_n422), .B2(new_n323), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n420), .B1(new_n421), .B2(new_n324), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT81), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n426), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT81), .B(new_n428), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT80), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G50gat), .ZN(new_n432));
  NAND2_X1  g231(.A1(G228gat), .A2(G233gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G22gat), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n432), .B(new_n434), .Z(new_n435));
  AND3_X1   g234(.A1(new_n427), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n435), .B1(new_n427), .B2(new_n429), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n397), .A2(new_n407), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n440), .A2(new_n403), .A3(new_n404), .ZN(new_n441));
  AND3_X1   g240(.A1(new_n412), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n420), .ZN(new_n443));
  INV_X1    g242(.A(G226gat), .ZN(new_n444));
  INV_X1    g243(.A(G233gat), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n386), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(KEYINPUT29), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n374), .B2(new_n385), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n374), .B(new_n385), .C1(new_n444), .C2(new_n445), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n420), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n451), .A2(KEYINPUT72), .A3(new_n420), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G64gat), .B(G92gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(G36gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT73), .B(G8gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  INV_X1    g262(.A(new_n457), .ZN(new_n464));
  XOR2_X1   g263(.A(new_n461), .B(KEYINPUT74), .Z(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n462), .A2(new_n463), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT35), .ZN(new_n468));
  INV_X1    g267(.A(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n469), .B1(new_n455), .B2(new_n456), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT30), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n352), .A2(new_n442), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT83), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n352), .A2(new_n442), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  OAI22_X1  g276(.A1(new_n470), .A2(KEYINPUT30), .B1(new_n457), .B2(new_n465), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(KEYINPUT30), .B2(new_n470), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n345), .A2(new_n351), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n405), .A2(KEYINPUT68), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n405), .A2(KEYINPUT68), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n482), .A2(new_n440), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n412), .A2(new_n439), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT35), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n475), .A2(new_n477), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n471), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n319), .A2(new_n329), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n322), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n490), .A2(KEYINPUT39), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n337), .A2(new_n321), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(KEYINPUT39), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n281), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n491), .A2(KEYINPUT40), .A3(new_n281), .A4(new_n493), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n496), .A2(new_n343), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n438), .B1(new_n488), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n461), .B1(new_n457), .B2(KEYINPUT38), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n450), .A2(new_n453), .ZN(new_n501));
  AOI211_X1 g300(.A(KEYINPUT38), .B(new_n465), .C1(new_n501), .C2(KEYINPUT37), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n457), .B(KEYINPUT37), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT38), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n500), .B(new_n503), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n499), .B1(new_n352), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n481), .A2(new_n438), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT36), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n412), .A2(new_n509), .A3(new_n441), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n509), .B1(new_n412), .B2(new_n484), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n508), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n276), .B1(new_n487), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G57gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G64gat), .ZN(new_n522));
  INV_X1    g321(.A(G64gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G57gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G71gat), .B(G78gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n519), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n520), .A2(new_n528), .A3(KEYINPUT90), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n239), .B1(KEYINPUT21), .B2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(new_n534), .B(G183gat), .Z(new_n535));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT89), .ZN(new_n537));
  XOR2_X1   g336(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n535), .B(new_n539), .Z(new_n540));
  AOI21_X1  g339(.A(KEYINPUT21), .B1(new_n520), .B2(new_n528), .ZN(new_n541));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(G211gat), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n540), .A2(new_n544), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(KEYINPUT41), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT91), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G134gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n303), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT92), .Z(new_n553));
  XNOR2_X1  g352(.A(G99gat), .B(G106gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(KEYINPUT8), .ZN(new_n560));
  NAND4_X1  g359(.A1(KEYINPUT93), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(KEYINPUT94), .A2(G85gat), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n564), .A2(new_n565), .A3(G92gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n555), .B1(new_n562), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g366(.A1(new_n560), .A2(new_n561), .ZN(new_n568));
  INV_X1    g367(.A(new_n565), .ZN(new_n569));
  INV_X1    g368(.A(G92gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n563), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n568), .A2(new_n571), .A3(new_n554), .A4(new_n558), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n574), .B1(new_n240), .B2(new_n241), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n233), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n240), .A2(new_n574), .B1(KEYINPUT41), .B2(new_n548), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G190gat), .B(G218gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT95), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n578), .A2(new_n581), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n578), .A2(KEYINPUT96), .A3(new_n581), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n553), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n582), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n583), .A3(new_n552), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n591));
  AND3_X1   g390(.A1(new_n520), .A2(new_n528), .A3(KEYINPUT90), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT90), .B1(new_n520), .B2(new_n528), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT10), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n591), .B1(new_n594), .B2(new_n573), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n520), .A2(new_n528), .A3(KEYINPUT97), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n520), .A2(new_n528), .A3(KEYINPUT97), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT97), .B1(new_n520), .B2(new_n528), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n596), .B(new_n598), .C1(new_n601), .C2(new_n573), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n533), .A2(new_n574), .A3(KEYINPUT98), .A4(KEYINPUT10), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n595), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G230gat), .A2(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G176gat), .ZN(new_n608));
  INV_X1    g407(.A(G204gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n598), .B1(new_n601), .B2(new_n573), .ZN(new_n611));
  INV_X1    g410(.A(new_n605), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n606), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT99), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n604), .A2(new_n615), .A3(new_n605), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n604), .B2(new_n605), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619));
  INV_X1    g418(.A(new_n610), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n614), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n547), .A2(new_n590), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n514), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n625), .A2(new_n480), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT101), .B(G1gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(G1324gat));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n514), .A2(new_n488), .A3(new_n624), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT102), .Z(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT16), .B(G8gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n630), .A2(new_n629), .A3(new_n632), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n634), .B1(new_n631), .B2(G8gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(G1325gat));
  INV_X1    g435(.A(G15gat), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n625), .A2(new_n637), .A3(new_n512), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n412), .A2(new_n441), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n637), .B1(new_n625), .B2(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(KEYINPUT103), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n638), .B1(new_n642), .B2(new_n643), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n625), .A2(new_n439), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  INV_X1    g446(.A(new_n623), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n547), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n590), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n514), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n480), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n204), .A2(new_n205), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT45), .ZN(new_n657));
  INV_X1    g456(.A(new_n271), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n649), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n351), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n346), .B2(new_n348), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n412), .A2(new_n439), .A3(new_n441), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n662), .A2(new_n663), .A3(new_n472), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n486), .B1(new_n664), .B2(new_n476), .ZN(new_n665));
  INV_X1    g464(.A(new_n477), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n513), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n590), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n650), .B1(new_n487), .B2(new_n513), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n660), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n673), .A2(new_n654), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n657), .B1(new_n655), .B2(new_n674), .ZN(G1328gat));
  NAND3_X1  g474(.A1(new_n653), .A2(new_n208), .A3(new_n488), .ZN(new_n676));
  AND2_X1   g475(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n677));
  NOR2_X1   g476(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n673), .A2(new_n488), .ZN(new_n680));
  OAI221_X1 g479(.A(new_n679), .B1(new_n677), .B2(new_n676), .C1(new_n680), .C2(new_n208), .ZN(G1329gat));
  INV_X1    g480(.A(G43gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n512), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n673), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n652), .A2(G43gat), .A3(new_n640), .ZN(new_n686));
  OR3_X1    g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1330gat));
  AOI211_X1 g488(.A(KEYINPUT44), .B(new_n650), .C1(new_n487), .C2(new_n513), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n671), .B1(new_n667), .B2(new_n590), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n438), .B(new_n659), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n667), .A2(new_n693), .A3(new_n275), .A4(new_n651), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n439), .A2(G50gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT106), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n693), .B1(new_n514), .B2(new_n651), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI22_X1  g499(.A1(new_n692), .A2(G50gat), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT107), .B1(new_n692), .B2(G50gat), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n697), .A2(new_n699), .ZN(new_n705));
  AOI221_X4 g504(.A(new_n705), .B1(KEYINPUT107), .B2(KEYINPUT48), .C1(G50gat), .C2(new_n692), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(G1331gat));
  INV_X1    g506(.A(new_n547), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n648), .A2(new_n271), .ZN(new_n709));
  AND4_X1   g508(.A1(new_n667), .A2(new_n708), .A3(new_n650), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n654), .ZN(new_n711));
  XOR2_X1   g510(.A(KEYINPUT108), .B(G57gat), .Z(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1332gat));
  AOI21_X1  g512(.A(new_n479), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT109), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT110), .ZN(new_n717));
  OR2_X1    g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1333gat));
  NAND2_X1  g518(.A1(new_n710), .A2(new_n683), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n640), .A2(G71gat), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n720), .A2(G71gat), .B1(new_n710), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g522(.A1(new_n710), .A2(new_n438), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT111), .B(G78gat), .Z(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(G1335gat));
  NAND2_X1  g525(.A1(new_n569), .A2(new_n563), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n480), .A2(new_n648), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n708), .A2(new_n271), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT51), .B1(new_n670), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n670), .A2(KEYINPUT51), .A3(new_n730), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n729), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n733), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n735), .A2(KEYINPUT112), .A3(new_n731), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n728), .B1(new_n734), .B2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n547), .B(new_n709), .C1(new_n690), .C2(new_n691), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n727), .B1(new_n738), .B2(new_n480), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1336gat));
  OAI21_X1  g539(.A(G92gat), .B1(new_n738), .B2(new_n479), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n479), .A2(G92gat), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n623), .B(new_n742), .C1(new_n735), .C2(new_n731), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n741), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n741), .B2(new_n743), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(G1337gat));
  XOR2_X1   g546(.A(KEYINPUT114), .B(G99gat), .Z(new_n748));
  NOR3_X1   g547(.A1(new_n640), .A2(new_n648), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n734), .B2(new_n736), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n748), .B1(new_n738), .B2(new_n512), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(G1338gat));
  OAI21_X1  g551(.A(G106gat), .B1(new_n738), .B2(new_n439), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n439), .A2(G106gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n623), .B(new_n754), .C1(new_n735), .C2(new_n731), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT53), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n753), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1339gat));
  NAND2_X1  g559(.A1(new_n606), .A2(KEYINPUT99), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT54), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n604), .A2(new_n615), .A3(new_n605), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n595), .A2(new_n602), .A3(new_n612), .A4(new_n603), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n765), .A2(new_n606), .A3(KEYINPUT54), .A4(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n762), .B1(new_n604), .B2(new_n605), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n765), .B1(new_n768), .B2(new_n766), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n620), .B(new_n764), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT55), .ZN(new_n771));
  OAI21_X1  g570(.A(KEYINPUT116), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n614), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n770), .B2(new_n771), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n616), .A2(new_n617), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n610), .B1(new_n775), .B2(new_n762), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n766), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT115), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n768), .A2(new_n765), .A3(new_n766), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n776), .A2(new_n780), .A3(new_n781), .A4(KEYINPUT55), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n772), .A2(new_n774), .A3(new_n271), .A4(new_n782), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n266), .A2(new_n244), .B1(new_n263), .B2(new_n264), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n257), .A2(new_n258), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n265), .A2(new_n261), .A3(new_n267), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n623), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n590), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n786), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n587), .B2(new_n589), .ZN(new_n791));
  AND4_X1   g590(.A1(new_n782), .A2(new_n791), .A3(new_n772), .A4(new_n774), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n547), .B1(new_n789), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n624), .A2(new_n658), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n793), .A2(KEYINPUT117), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT117), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n663), .A2(new_n480), .A3(new_n488), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n276), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n795), .A2(new_n796), .A3(new_n480), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n485), .A2(new_n488), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(KEYINPUT118), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n271), .A2(new_n282), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n800), .B1(new_n808), .B2(new_n809), .ZN(G1340gat));
  OAI21_X1  g609(.A(G120gat), .B1(new_n799), .B2(new_n648), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(KEYINPUT119), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n623), .A2(new_n283), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n812), .B(KEYINPUT120), .C1(new_n808), .C2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n811), .B(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n813), .B1(new_n805), .B2(new_n807), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(G1341gat));
  NAND4_X1  g619(.A1(new_n797), .A2(G127gat), .A3(new_n708), .A4(new_n798), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT121), .ZN(new_n822));
  AOI21_X1  g621(.A(G127gat), .B1(new_n804), .B2(new_n708), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(G1342gat));
  OR3_X1    g623(.A1(new_n803), .A2(G134gat), .A3(new_n650), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n799), .B2(new_n650), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(KEYINPUT56), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(G1343gat));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n683), .A2(new_n439), .A3(new_n488), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n801), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n833), .A2(new_n296), .A3(new_n275), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n439), .A2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n772), .A2(new_n774), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n275), .A3(new_n782), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n590), .B1(new_n839), .B2(new_n788), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n547), .B1(new_n840), .B2(new_n792), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n837), .B1(new_n841), .B2(new_n794), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n793), .A2(new_n794), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n793), .A2(KEYINPUT117), .A3(new_n794), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(new_n438), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n842), .B1(new_n847), .B2(new_n835), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n512), .A2(new_n654), .A3(new_n479), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n276), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G141gat), .B1(new_n850), .B2(KEYINPUT123), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n848), .A2(new_n849), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n852), .A2(KEYINPUT123), .A3(new_n275), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n830), .B(new_n834), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n841), .A2(new_n794), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n836), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n795), .A2(new_n796), .A3(new_n439), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(KEYINPUT57), .ZN(new_n858));
  INV_X1    g657(.A(new_n849), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n271), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(G141gat), .ZN(new_n861));
  AOI211_X1 g660(.A(KEYINPUT122), .B(new_n830), .C1(new_n861), .C2(new_n834), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n848), .A2(new_n658), .A3(new_n849), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n834), .B1(new_n864), .B2(new_n296), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(KEYINPUT58), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n854), .B1(new_n862), .B2(new_n866), .ZN(G1344gat));
  NAND3_X1  g666(.A1(new_n833), .A2(new_n298), .A3(new_n623), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n869));
  INV_X1    g668(.A(new_n624), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n841), .B1(new_n275), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n871), .B2(new_n438), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n795), .A2(new_n796), .A3(new_n837), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n623), .A3(new_n859), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n869), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  AOI211_X1 g676(.A(KEYINPUT59), .B(new_n298), .C1(new_n852), .C2(new_n623), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n868), .B1(new_n877), .B2(new_n878), .ZN(G1345gat));
  NAND3_X1  g678(.A1(new_n833), .A2(new_n302), .A3(new_n708), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n848), .A2(new_n547), .A3(new_n849), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n302), .ZN(G1346gat));
  NAND3_X1  g681(.A1(new_n833), .A2(new_n303), .A3(new_n590), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n848), .A2(new_n650), .A3(new_n849), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n884), .B2(new_n303), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n479), .A2(new_n654), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n797), .A2(new_n442), .A3(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n254), .A3(new_n276), .ZN(new_n888));
  INV_X1    g687(.A(new_n485), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n797), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n271), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n888), .B1(new_n892), .B2(new_n254), .ZN(G1348gat));
  OAI21_X1  g692(.A(G176gat), .B1(new_n887), .B2(new_n648), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n623), .A2(new_n353), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n890), .B2(new_n895), .ZN(G1349gat));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n708), .A2(new_n378), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n890), .B2(new_n898), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n797), .A2(new_n886), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n442), .A3(new_n708), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n903), .A2(G183gat), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n904));
  OR2_X1    g703(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n901), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n905), .B1(new_n901), .B2(new_n904), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n380), .A3(new_n590), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n902), .A2(new_n442), .A3(new_n590), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(G190gat), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n910), .B(G190gat), .C1(new_n887), .C2(new_n650), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n909), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(KEYINPUT126), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n909), .B(new_n917), .C1(new_n912), .C2(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1351gat));
  NAND2_X1  g718(.A1(new_n512), .A2(new_n886), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n857), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(G197gat), .B1(new_n923), .B2(new_n271), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n875), .A2(KEYINPUT127), .ZN(new_n925));
  OR3_X1    g724(.A1(new_n872), .A2(KEYINPUT127), .A3(new_n873), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n920), .A2(new_n256), .A3(new_n276), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(G1352gat));
  NOR3_X1   g728(.A1(new_n922), .A2(G204gat), .A3(new_n648), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT62), .ZN(new_n931));
  AOI211_X1 g730(.A(new_n648), .B(new_n920), .C1(new_n925), .C2(new_n926), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n932), .B2(new_n609), .ZN(G1353gat));
  OR3_X1    g732(.A1(new_n922), .A2(G211gat), .A3(new_n547), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n875), .A2(new_n708), .A3(new_n921), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n936));
  AOI21_X1  g735(.A(KEYINPUT63), .B1(new_n935), .B2(G211gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  AOI21_X1  g737(.A(G218gat), .B1(new_n923), .B2(new_n590), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n921), .A2(G218gat), .A3(new_n590), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n927), .B2(new_n940), .ZN(G1355gat));
endmodule


