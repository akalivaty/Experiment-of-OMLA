

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n607), .A2(n563), .ZN(n797) );
  NOR2_X1 U551 ( .A1(n718), .A2(n655), .ZN(n545) );
  NAND2_X1 U552 ( .A1(G8), .A2(n724), .ZN(n750) );
  INV_X1 U553 ( .A(n698), .ZN(n724) );
  NOR2_X2 U554 ( .A1(G164), .A2(n524), .ZN(n698) );
  XNOR2_X1 U555 ( .A(n526), .B(n525), .ZN(G164) );
  OR2_X1 U556 ( .A1(n655), .A2(n541), .ZN(n540) );
  OR2_X1 U557 ( .A1(n720), .A2(n542), .ZN(n541) );
  INV_X1 U558 ( .A(G8), .ZN(n542) );
  AND2_X1 U559 ( .A1(n746), .A2(n522), .ZN(n543) );
  OR2_X1 U560 ( .A1(n651), .A2(G1384), .ZN(n524) );
  NAND2_X1 U561 ( .A1(n533), .A2(n531), .ZN(n530) );
  NAND2_X1 U562 ( .A1(n743), .A2(n532), .ZN(n531) );
  NAND2_X1 U563 ( .A1(n534), .A2(KEYINPUT107), .ZN(n533) );
  NAND2_X1 U564 ( .A1(n750), .A2(KEYINPUT107), .ZN(n532) );
  NAND2_X1 U565 ( .A1(n547), .A2(n551), .ZN(n546) );
  INV_X1 U566 ( .A(G2105), .ZN(n547) );
  NAND2_X1 U567 ( .A1(n518), .A2(n521), .ZN(n539) );
  NOR2_X1 U568 ( .A1(n754), .A2(n520), .ZN(n538) );
  XNOR2_X1 U569 ( .A(n540), .B(KEYINPUT30), .ZN(n656) );
  XNOR2_X1 U570 ( .A(KEYINPUT31), .B(KEYINPUT103), .ZN(n662) );
  INV_X1 U571 ( .A(n743), .ZN(n534) );
  XNOR2_X1 U572 ( .A(n732), .B(KEYINPUT32), .ZN(n746) );
  NAND2_X1 U573 ( .A1(n528), .A2(n519), .ZN(n527) );
  AND2_X1 U574 ( .A1(n535), .A2(n530), .ZN(n529) );
  XNOR2_X1 U575 ( .A(KEYINPUT15), .B(n689), .ZN(n1024) );
  NAND2_X1 U576 ( .A1(n537), .A2(n770), .ZN(n771) );
  INV_X1 U577 ( .A(KEYINPUT86), .ZN(n525) );
  OR2_X1 U578 ( .A1(n577), .A2(n576), .ZN(n526) );
  NOR2_X2 U579 ( .A1(n555), .A2(n554), .ZN(G160) );
  AND2_X1 U580 ( .A1(n753), .A2(n752), .ZN(n518) );
  AND2_X1 U581 ( .A1(n743), .A2(KEYINPUT107), .ZN(n519) );
  NOR2_X2 U582 ( .A1(G2105), .A2(n551), .ZN(n573) );
  AND2_X1 U583 ( .A1(n859), .A2(n767), .ZN(n520) );
  OR2_X1 U584 ( .A1(n750), .A2(n653), .ZN(n521) );
  AND2_X1 U585 ( .A1(n853), .A2(n733), .ZN(n522) );
  AND2_X1 U586 ( .A1(n740), .A2(n744), .ZN(n523) );
  NAND2_X1 U587 ( .A1(n529), .A2(n527), .ZN(n536) );
  INV_X1 U588 ( .A(n739), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n739), .A2(n523), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n848), .ZN(n753) );
  NAND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n745), .A2(n543), .ZN(n738) );
  NAND2_X1 U593 ( .A1(n544), .A2(n722), .ZN(n745) );
  XNOR2_X1 U594 ( .A(n545), .B(n719), .ZN(n544) );
  XNOR2_X2 U595 ( .A(n546), .B(KEYINPUT17), .ZN(n1000) );
  NOR2_X1 U596 ( .A1(n695), .A2(n781), .ZN(n690) );
  INV_X1 U597 ( .A(KEYINPUT105), .ZN(n719) );
  INV_X1 U598 ( .A(KEYINPUT107), .ZN(n744) );
  INV_X1 U599 ( .A(KEYINPUT13), .ZN(n672) );
  XNOR2_X1 U600 ( .A(n672), .B(KEYINPUT68), .ZN(n673) );
  XNOR2_X1 U601 ( .A(n674), .B(n673), .ZN(n675) );
  NOR2_X1 U602 ( .A1(G651), .A2(n607), .ZN(n801) );
  INV_X1 U603 ( .A(G2104), .ZN(n551) );
  AND2_X1 U604 ( .A1(G2105), .A2(G2104), .ZN(n995) );
  NAND2_X1 U605 ( .A1(n995), .A2(G113), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G101), .A2(n573), .ZN(n548) );
  XOR2_X1 U607 ( .A(KEYINPUT23), .B(n548), .Z(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n555) );
  NAND2_X1 U609 ( .A1(G137), .A2(n1000), .ZN(n553) );
  AND2_X1 U610 ( .A1(n551), .A2(G2105), .ZN(n996) );
  NAND2_X1 U611 ( .A1(G125), .A2(n996), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U613 ( .A1(G543), .A2(G651), .ZN(n556) );
  XNOR2_X1 U614 ( .A(n556), .B(KEYINPUT64), .ZN(n798) );
  NAND2_X1 U615 ( .A1(G89), .A2(n798), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n557), .B(KEYINPUT4), .ZN(n560) );
  XNOR2_X1 U617 ( .A(G543), .B(KEYINPUT0), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT65), .ZN(n607) );
  XOR2_X1 U619 ( .A(G651), .B(KEYINPUT66), .Z(n563) );
  NAND2_X1 U620 ( .A1(G76), .A2(n797), .ZN(n559) );
  NAND2_X1 U621 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n561), .B(KEYINPUT5), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n801), .A2(G51), .ZN(n562) );
  XNOR2_X1 U624 ( .A(n562), .B(KEYINPUT72), .ZN(n566) );
  NOR2_X1 U625 ( .A1(G543), .A2(n563), .ZN(n564) );
  XOR2_X2 U626 ( .A(KEYINPUT1), .B(n564), .Z(n796) );
  NAND2_X1 U627 ( .A1(G63), .A2(n796), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n567), .Z(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(G138), .A2(n1000), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G126), .A2(n996), .ZN(n571) );
  NAND2_X1 U635 ( .A1(n572), .A2(n571), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G102), .A2(n573), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G114), .A2(n995), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U639 ( .A1(G73), .A2(n797), .ZN(n578) );
  XNOR2_X1 U640 ( .A(n578), .B(KEYINPUT2), .ZN(n585) );
  NAND2_X1 U641 ( .A1(G61), .A2(n796), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G48), .A2(n801), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U644 ( .A1(G86), .A2(n798), .ZN(n581) );
  XNOR2_X1 U645 ( .A(KEYINPUT79), .B(n581), .ZN(n582) );
  NOR2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n585), .A2(n584), .ZN(G305) );
  NAND2_X1 U648 ( .A1(n801), .A2(G52), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n796), .A2(G64), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U651 ( .A1(n797), .A2(G77), .ZN(n589) );
  NAND2_X1 U652 ( .A1(G90), .A2(n798), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT9), .B(n590), .Z(n591) );
  NOR2_X1 U655 ( .A1(n592), .A2(n591), .ZN(G171) );
  NAND2_X1 U656 ( .A1(G65), .A2(n796), .ZN(n594) );
  NAND2_X1 U657 ( .A1(G53), .A2(n801), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U659 ( .A1(n797), .A2(G78), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G91), .A2(n798), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n597) );
  OR2_X1 U662 ( .A1(n598), .A2(n597), .ZN(G299) );
  NAND2_X1 U663 ( .A1(n797), .A2(G75), .ZN(n600) );
  NAND2_X1 U664 ( .A1(G88), .A2(n798), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U666 ( .A(KEYINPUT80), .B(n601), .Z(n605) );
  NAND2_X1 U667 ( .A1(G62), .A2(n796), .ZN(n603) );
  NAND2_X1 U668 ( .A1(G50), .A2(n801), .ZN(n602) );
  AND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U670 ( .A1(n605), .A2(n604), .ZN(G303) );
  NAND2_X1 U671 ( .A1(G49), .A2(n801), .ZN(n606) );
  XNOR2_X1 U672 ( .A(n606), .B(KEYINPUT78), .ZN(n612) );
  NAND2_X1 U673 ( .A1(G87), .A2(n607), .ZN(n609) );
  NAND2_X1 U674 ( .A1(G74), .A2(G651), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U676 ( .A1(n796), .A2(n610), .ZN(n611) );
  NAND2_X1 U677 ( .A1(n612), .A2(n611), .ZN(G288) );
  NAND2_X1 U678 ( .A1(G60), .A2(n796), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G47), .A2(n801), .ZN(n613) );
  NAND2_X1 U680 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U681 ( .A(KEYINPUT67), .B(n615), .ZN(n619) );
  NAND2_X1 U682 ( .A1(n798), .A2(G85), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n797), .A2(G72), .ZN(n616) );
  AND2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n619), .A2(n618), .ZN(G290) );
  NOR2_X1 U686 ( .A1(G1384), .A2(G164), .ZN(n620) );
  NAND2_X1 U687 ( .A1(G160), .A2(G40), .ZN(n651) );
  NOR2_X1 U688 ( .A1(n620), .A2(n651), .ZN(n767) );
  NAND2_X1 U689 ( .A1(n1000), .A2(G140), .ZN(n621) );
  XOR2_X1 U690 ( .A(KEYINPUT87), .B(n621), .Z(n623) );
  NAND2_X1 U691 ( .A1(n573), .A2(G104), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U693 ( .A(KEYINPUT34), .B(n624), .ZN(n629) );
  NAND2_X1 U694 ( .A1(G116), .A2(n995), .ZN(n626) );
  NAND2_X1 U695 ( .A1(G128), .A2(n996), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U697 ( .A(KEYINPUT35), .B(n627), .Z(n628) );
  NOR2_X1 U698 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U699 ( .A(KEYINPUT36), .B(n630), .ZN(n1012) );
  XNOR2_X1 U700 ( .A(G2067), .B(KEYINPUT37), .ZN(n765) );
  NOR2_X1 U701 ( .A1(n1012), .A2(n765), .ZN(n946) );
  NAND2_X1 U702 ( .A1(n767), .A2(n946), .ZN(n764) );
  INV_X1 U703 ( .A(G1996), .ZN(n985) );
  NAND2_X1 U704 ( .A1(G141), .A2(n1000), .ZN(n639) );
  XOR2_X1 U705 ( .A(KEYINPUT38), .B(KEYINPUT90), .Z(n632) );
  NAND2_X1 U706 ( .A1(G105), .A2(n573), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n632), .B(n631), .ZN(n636) );
  NAND2_X1 U708 ( .A1(G117), .A2(n995), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G129), .A2(n996), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U712 ( .A(KEYINPUT91), .B(n637), .Z(n638) );
  NAND2_X1 U713 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U714 ( .A(n640), .B(KEYINPUT92), .Z(n1011) );
  NOR2_X1 U715 ( .A1(n985), .A2(n1011), .ZN(n649) );
  NAND2_X1 U716 ( .A1(G95), .A2(n573), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G131), .A2(n1000), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U719 ( .A(KEYINPUT88), .B(n643), .Z(n647) );
  NAND2_X1 U720 ( .A1(G107), .A2(n995), .ZN(n645) );
  NAND2_X1 U721 ( .A1(G119), .A2(n996), .ZN(n644) );
  AND2_X1 U722 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n1018) );
  XOR2_X1 U724 ( .A(G1991), .B(KEYINPUT89), .Z(n900) );
  AND2_X1 U725 ( .A1(n1018), .A2(n900), .ZN(n648) );
  NOR2_X1 U726 ( .A1(n649), .A2(n648), .ZN(n922) );
  INV_X1 U727 ( .A(n922), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n650), .A2(n767), .ZN(n755) );
  NAND2_X1 U729 ( .A1(n764), .A2(n755), .ZN(n754) );
  NOR2_X1 U730 ( .A1(G1981), .A2(G305), .ZN(n652) );
  XOR2_X1 U731 ( .A(n652), .B(KEYINPUT24), .Z(n653) );
  NOR2_X1 U732 ( .A1(G1966), .A2(n750), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n654), .B(KEYINPUT94), .ZN(n655) );
  NOR2_X1 U734 ( .A1(G2084), .A2(n724), .ZN(n720) );
  NOR2_X1 U735 ( .A1(G168), .A2(n656), .ZN(n661) );
  XOR2_X1 U736 ( .A(G2078), .B(KEYINPUT25), .Z(n903) );
  NOR2_X1 U737 ( .A1(n903), .A2(n724), .ZN(n657) );
  XNOR2_X1 U738 ( .A(n657), .B(KEYINPUT95), .ZN(n659) );
  INV_X1 U739 ( .A(G1961), .ZN(n990) );
  NAND2_X1 U740 ( .A1(n990), .A2(n724), .ZN(n658) );
  NAND2_X1 U741 ( .A1(n659), .A2(n658), .ZN(n713) );
  NOR2_X1 U742 ( .A1(G171), .A2(n713), .ZN(n660) );
  NOR2_X1 U743 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U744 ( .A(n663), .B(n662), .ZN(n717) );
  XOR2_X1 U745 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n665) );
  XNOR2_X1 U746 ( .A(n985), .B(KEYINPUT97), .ZN(n909) );
  NAND2_X1 U747 ( .A1(n909), .A2(n698), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n665), .B(n664), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n796), .A2(G56), .ZN(n666) );
  XNOR2_X1 U750 ( .A(n666), .B(KEYINPUT14), .ZN(n668) );
  NAND2_X1 U751 ( .A1(G43), .A2(n801), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n676) );
  NAND2_X1 U753 ( .A1(G81), .A2(n798), .ZN(n669) );
  XNOR2_X1 U754 ( .A(n669), .B(KEYINPUT12), .ZN(n671) );
  NAND2_X1 U755 ( .A1(G68), .A2(n797), .ZN(n670) );
  NAND2_X1 U756 ( .A1(n671), .A2(n670), .ZN(n674) );
  NOR2_X1 U757 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U758 ( .A(KEYINPUT69), .B(n677), .ZN(n774) );
  NOR2_X1 U759 ( .A1(n678), .A2(n774), .ZN(n680) );
  NAND2_X1 U760 ( .A1(G1341), .A2(n724), .ZN(n679) );
  NAND2_X1 U761 ( .A1(n680), .A2(n679), .ZN(n695) );
  NAND2_X1 U762 ( .A1(G66), .A2(n796), .ZN(n681) );
  XNOR2_X1 U763 ( .A(n681), .B(KEYINPUT70), .ZN(n688) );
  NAND2_X1 U764 ( .A1(n801), .A2(G54), .ZN(n683) );
  NAND2_X1 U765 ( .A1(G92), .A2(n798), .ZN(n682) );
  NAND2_X1 U766 ( .A1(n683), .A2(n682), .ZN(n686) );
  NAND2_X1 U767 ( .A1(G79), .A2(n797), .ZN(n684) );
  XNOR2_X1 U768 ( .A(KEYINPUT71), .B(n684), .ZN(n685) );
  NOR2_X1 U769 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n688), .A2(n687), .ZN(n689) );
  INV_X1 U771 ( .A(n1024), .ZN(n781) );
  XNOR2_X1 U772 ( .A(n690), .B(KEYINPUT99), .ZN(n694) );
  NOR2_X1 U773 ( .A1(G2067), .A2(n724), .ZN(n692) );
  NOR2_X1 U774 ( .A1(n698), .A2(G1348), .ZN(n691) );
  NOR2_X1 U775 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U776 ( .A1(n694), .A2(n693), .ZN(n697) );
  NAND2_X1 U777 ( .A1(n695), .A2(n781), .ZN(n696) );
  NAND2_X1 U778 ( .A1(n697), .A2(n696), .ZN(n705) );
  NAND2_X1 U779 ( .A1(n724), .A2(G1956), .ZN(n701) );
  NAND2_X1 U780 ( .A1(n698), .A2(G2072), .ZN(n699) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(n699), .Z(n700) );
  NAND2_X1 U782 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U783 ( .A(n702), .B(KEYINPUT96), .ZN(n706) );
  NOR2_X1 U784 ( .A1(n706), .A2(G299), .ZN(n703) );
  XOR2_X1 U785 ( .A(KEYINPUT100), .B(n703), .Z(n704) );
  NAND2_X1 U786 ( .A1(n705), .A2(n704), .ZN(n709) );
  NAND2_X1 U787 ( .A1(n706), .A2(G299), .ZN(n707) );
  XNOR2_X1 U788 ( .A(n707), .B(KEYINPUT28), .ZN(n708) );
  NAND2_X1 U789 ( .A1(n709), .A2(n708), .ZN(n712) );
  XNOR2_X1 U790 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n710) );
  XNOR2_X1 U791 ( .A(n710), .B(KEYINPUT29), .ZN(n711) );
  XNOR2_X1 U792 ( .A(n712), .B(n711), .ZN(n715) );
  NAND2_X1 U793 ( .A1(n713), .A2(G171), .ZN(n714) );
  NAND2_X1 U794 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U795 ( .A1(n717), .A2(n716), .ZN(n723) );
  XOR2_X1 U796 ( .A(n723), .B(KEYINPUT104), .Z(n718) );
  NAND2_X1 U797 ( .A1(G8), .A2(n720), .ZN(n721) );
  XOR2_X1 U798 ( .A(KEYINPUT93), .B(n721), .Z(n722) );
  NAND2_X1 U799 ( .A1(n723), .A2(G286), .ZN(n730) );
  NOR2_X1 U800 ( .A1(G1971), .A2(n750), .ZN(n726) );
  NOR2_X1 U801 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U802 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U803 ( .A1(n727), .A2(G303), .ZN(n728) );
  XNOR2_X1 U804 ( .A(n728), .B(KEYINPUT106), .ZN(n729) );
  NAND2_X1 U805 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U806 ( .A1(n731), .A2(G8), .ZN(n732) );
  NAND2_X1 U807 ( .A1(G1976), .A2(G288), .ZN(n853) );
  INV_X1 U808 ( .A(KEYINPUT33), .ZN(n733) );
  INV_X1 U809 ( .A(n853), .ZN(n735) );
  NOR2_X1 U810 ( .A1(G1976), .A2(G288), .ZN(n741) );
  NOR2_X1 U811 ( .A1(G1971), .A2(G303), .ZN(n734) );
  NOR2_X1 U812 ( .A1(n741), .A2(n734), .ZN(n861) );
  OR2_X1 U813 ( .A1(n735), .A2(n861), .ZN(n736) );
  OR2_X1 U814 ( .A1(KEYINPUT33), .A2(n736), .ZN(n737) );
  NAND2_X1 U815 ( .A1(n738), .A2(n737), .ZN(n739) );
  INV_X1 U816 ( .A(n750), .ZN(n740) );
  NAND2_X1 U817 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U818 ( .A1(n742), .A2(KEYINPUT33), .ZN(n743) );
  XOR2_X1 U819 ( .A(G1981), .B(G305), .Z(n848) );
  NAND2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n749) );
  NOR2_X1 U821 ( .A1(G2090), .A2(G303), .ZN(n747) );
  NAND2_X1 U822 ( .A1(G8), .A2(n747), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n749), .A2(n748), .ZN(n751) );
  NAND2_X1 U824 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U825 ( .A(G1986), .B(G290), .ZN(n859) );
  XOR2_X1 U826 ( .A(KEYINPUT39), .B(KEYINPUT109), .Z(n762) );
  AND2_X1 U827 ( .A1(n985), .A2(n1011), .ZN(n939) );
  INV_X1 U828 ( .A(n755), .ZN(n758) );
  NOR2_X1 U829 ( .A1(G1986), .A2(G290), .ZN(n756) );
  NOR2_X1 U830 ( .A1(n900), .A2(n1018), .ZN(n924) );
  NOR2_X1 U831 ( .A1(n756), .A2(n924), .ZN(n757) );
  NOR2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U833 ( .A1(n939), .A2(n759), .ZN(n760) );
  XNOR2_X1 U834 ( .A(n760), .B(KEYINPUT108), .ZN(n761) );
  XNOR2_X1 U835 ( .A(n762), .B(n761), .ZN(n763) );
  NAND2_X1 U836 ( .A1(n764), .A2(n763), .ZN(n766) );
  NAND2_X1 U837 ( .A1(n1012), .A2(n765), .ZN(n936) );
  NAND2_X1 U838 ( .A1(n766), .A2(n936), .ZN(n768) );
  NAND2_X1 U839 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U840 ( .A(KEYINPUT110), .B(n769), .ZN(n770) );
  XNOR2_X1 U841 ( .A(n771), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(G171), .ZN(G301) );
  INV_X1 U844 ( .A(G57), .ZN(G237) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n772) );
  XOR2_X1 U846 ( .A(n772), .B(KEYINPUT10), .Z(n836) );
  NAND2_X1 U847 ( .A1(n836), .A2(G567), .ZN(n773) );
  XOR2_X1 U848 ( .A(KEYINPUT11), .B(n773), .Z(G234) );
  INV_X1 U849 ( .A(n774), .ZN(n1027) );
  NAND2_X1 U850 ( .A1(n1027), .A2(G860), .ZN(G153) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n776) );
  INV_X1 U852 ( .A(G868), .ZN(n808) );
  NAND2_X1 U853 ( .A1(n781), .A2(n808), .ZN(n775) );
  NAND2_X1 U854 ( .A1(n776), .A2(n775), .ZN(G284) );
  NOR2_X1 U855 ( .A1(G286), .A2(n808), .ZN(n778) );
  NOR2_X1 U856 ( .A1(G868), .A2(G299), .ZN(n777) );
  NOR2_X1 U857 ( .A1(n778), .A2(n777), .ZN(G297) );
  INV_X1 U858 ( .A(G860), .ZN(n959) );
  NAND2_X1 U859 ( .A1(n959), .A2(G559), .ZN(n779) );
  NAND2_X1 U860 ( .A1(n779), .A2(n1024), .ZN(n780) );
  XNOR2_X1 U861 ( .A(n780), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U862 ( .A1(G559), .A2(n781), .ZN(n782) );
  NOR2_X1 U863 ( .A1(n808), .A2(n782), .ZN(n784) );
  NOR2_X1 U864 ( .A1(n1027), .A2(G868), .ZN(n783) );
  NOR2_X1 U865 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U866 ( .A(KEYINPUT73), .B(n785), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G99), .A2(n573), .ZN(n787) );
  NAND2_X1 U868 ( .A1(G111), .A2(n995), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n787), .A2(n786), .ZN(n794) );
  NAND2_X1 U870 ( .A1(G123), .A2(n996), .ZN(n788) );
  XNOR2_X1 U871 ( .A(n788), .B(KEYINPUT18), .ZN(n789) );
  XNOR2_X1 U872 ( .A(n789), .B(KEYINPUT74), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G135), .A2(n1000), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n792) );
  XOR2_X1 U875 ( .A(KEYINPUT75), .B(n792), .Z(n793) );
  NOR2_X1 U876 ( .A1(n794), .A2(n793), .ZN(n1007) );
  XNOR2_X1 U877 ( .A(n1007), .B(G2096), .ZN(n795) );
  INV_X1 U878 ( .A(G2100), .ZN(n978) );
  NAND2_X1 U879 ( .A1(n795), .A2(n978), .ZN(G156) );
  NAND2_X1 U880 ( .A1(n796), .A2(G67), .ZN(n806) );
  NAND2_X1 U881 ( .A1(n797), .A2(G80), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G93), .A2(n798), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n804) );
  NAND2_X1 U884 ( .A1(n801), .A2(G55), .ZN(n802) );
  XOR2_X1 U885 ( .A(KEYINPUT76), .B(n802), .Z(n803) );
  NOR2_X1 U886 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U887 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U888 ( .A(KEYINPUT77), .B(n807), .ZN(n960) );
  INV_X1 U889 ( .A(n960), .ZN(n810) );
  NAND2_X1 U890 ( .A1(n808), .A2(n810), .ZN(n809) );
  XNOR2_X1 U891 ( .A(n809), .B(KEYINPUT82), .ZN(n820) );
  XOR2_X1 U892 ( .A(n810), .B(G290), .Z(n816) );
  XNOR2_X1 U893 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n812) );
  XOR2_X1 U894 ( .A(G299), .B(G303), .Z(n811) );
  XNOR2_X1 U895 ( .A(n812), .B(n811), .ZN(n813) );
  XOR2_X1 U896 ( .A(n813), .B(G305), .Z(n814) );
  XNOR2_X1 U897 ( .A(G288), .B(n814), .ZN(n815) );
  XNOR2_X1 U898 ( .A(n816), .B(n815), .ZN(n1023) );
  NAND2_X1 U899 ( .A1(G559), .A2(n1024), .ZN(n817) );
  XNOR2_X1 U900 ( .A(n1027), .B(n817), .ZN(n958) );
  XNOR2_X1 U901 ( .A(n1023), .B(n958), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G868), .A2(n818), .ZN(n819) );
  NAND2_X1 U903 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U904 ( .A(KEYINPUT83), .B(n821), .Z(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n822) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n822), .Z(n823) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n823), .ZN(n824) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n824), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(KEYINPUT84), .B(G44), .ZN(n826) );
  XNOR2_X1 U911 ( .A(n826), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(KEYINPUT85), .Z(n828) );
  NAND2_X1 U913 ( .A1(G132), .A2(G82), .ZN(n827) );
  XNOR2_X1 U914 ( .A(n828), .B(n827), .ZN(n829) );
  NOR2_X1 U915 ( .A1(G218), .A2(n829), .ZN(n830) );
  NAND2_X1 U916 ( .A1(G96), .A2(n830), .ZN(n956) );
  NAND2_X1 U917 ( .A1(n956), .A2(G2106), .ZN(n834) );
  NAND2_X1 U918 ( .A1(G69), .A2(G120), .ZN(n831) );
  NOR2_X1 U919 ( .A1(G237), .A2(n831), .ZN(n832) );
  NAND2_X1 U920 ( .A1(G108), .A2(n832), .ZN(n957) );
  NAND2_X1 U921 ( .A1(n957), .A2(G567), .ZN(n833) );
  NAND2_X1 U922 ( .A1(n834), .A2(n833), .ZN(n972) );
  NAND2_X1 U923 ( .A1(G483), .A2(G661), .ZN(n835) );
  NOR2_X1 U924 ( .A1(n972), .A2(n835), .ZN(n838) );
  NAND2_X1 U925 ( .A1(n838), .A2(G36), .ZN(G176) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n836), .ZN(G217) );
  INV_X1 U927 ( .A(n836), .ZN(G223) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U929 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G1), .A2(G3), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U932 ( .A(n840), .B(KEYINPUT112), .ZN(G188) );
  NAND2_X1 U934 ( .A1(G124), .A2(n996), .ZN(n841) );
  XNOR2_X1 U935 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U936 ( .A1(n995), .A2(G112), .ZN(n842) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U938 ( .A1(G100), .A2(n573), .ZN(n845) );
  NAND2_X1 U939 ( .A1(G136), .A2(n1000), .ZN(n844) );
  NAND2_X1 U940 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U941 ( .A1(n847), .A2(n846), .ZN(G162) );
  XNOR2_X1 U942 ( .A(G1966), .B(G168), .ZN(n849) );
  NAND2_X1 U943 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U944 ( .A(n850), .B(KEYINPUT57), .ZN(n851) );
  XNOR2_X1 U945 ( .A(KEYINPUT124), .B(n851), .ZN(n865) );
  XOR2_X1 U946 ( .A(G301), .B(G1961), .Z(n857) );
  NAND2_X1 U947 ( .A1(G1971), .A2(G303), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n853), .A2(n852), .ZN(n855) );
  XNOR2_X1 U949 ( .A(G1956), .B(G299), .ZN(n854) );
  NOR2_X1 U950 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U951 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U952 ( .A1(n859), .A2(n858), .ZN(n860) );
  NAND2_X1 U953 ( .A1(n861), .A2(n860), .ZN(n863) );
  XOR2_X1 U954 ( .A(G1341), .B(n1027), .Z(n862) );
  NOR2_X1 U955 ( .A1(n863), .A2(n862), .ZN(n864) );
  NAND2_X1 U956 ( .A1(n865), .A2(n864), .ZN(n867) );
  XOR2_X1 U957 ( .A(G1348), .B(n1024), .Z(n866) );
  NOR2_X1 U958 ( .A1(n867), .A2(n866), .ZN(n869) );
  INV_X1 U959 ( .A(G16), .ZN(n892) );
  XNOR2_X1 U960 ( .A(n892), .B(KEYINPUT56), .ZN(n868) );
  NOR2_X1 U961 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U962 ( .A(KEYINPUT125), .B(n870), .ZN(n954) );
  XOR2_X1 U963 ( .A(G1986), .B(G24), .Z(n874) );
  XNOR2_X1 U964 ( .A(G1971), .B(G22), .ZN(n872) );
  XNOR2_X1 U965 ( .A(G23), .B(G1976), .ZN(n871) );
  NOR2_X1 U966 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U967 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U968 ( .A(KEYINPUT58), .B(n875), .ZN(n890) );
  XNOR2_X1 U969 ( .A(G1348), .B(KEYINPUT59), .ZN(n876) );
  XNOR2_X1 U970 ( .A(n876), .B(G4), .ZN(n880) );
  XNOR2_X1 U971 ( .A(G1341), .B(G19), .ZN(n878) );
  XNOR2_X1 U972 ( .A(G1981), .B(G6), .ZN(n877) );
  NOR2_X1 U973 ( .A1(n878), .A2(n877), .ZN(n879) );
  NAND2_X1 U974 ( .A1(n880), .A2(n879), .ZN(n882) );
  XNOR2_X1 U975 ( .A(G20), .B(G1956), .ZN(n881) );
  NOR2_X1 U976 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U977 ( .A(KEYINPUT60), .B(n883), .Z(n885) );
  XNOR2_X1 U978 ( .A(G1966), .B(G21), .ZN(n884) );
  NOR2_X1 U979 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U980 ( .A(KEYINPUT126), .B(n886), .ZN(n888) );
  XOR2_X1 U981 ( .A(G1961), .B(G5), .Z(n887) );
  NAND2_X1 U982 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U983 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U984 ( .A(KEYINPUT61), .B(n891), .ZN(n893) );
  NAND2_X1 U985 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U986 ( .A1(n894), .A2(G11), .ZN(n952) );
  XOR2_X1 U987 ( .A(KEYINPUT123), .B(G34), .Z(n896) );
  XNOR2_X1 U988 ( .A(G2084), .B(KEYINPUT54), .ZN(n895) );
  XNOR2_X1 U989 ( .A(n896), .B(n895), .ZN(n917) );
  XOR2_X1 U990 ( .A(G2090), .B(G35), .Z(n897) );
  XNOR2_X1 U991 ( .A(KEYINPUT119), .B(n897), .ZN(n914) );
  XNOR2_X1 U992 ( .A(G2067), .B(G26), .ZN(n899) );
  XNOR2_X1 U993 ( .A(G33), .B(G2072), .ZN(n898) );
  NOR2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n908) );
  XOR2_X1 U995 ( .A(n900), .B(G25), .Z(n901) );
  NAND2_X1 U996 ( .A1(n901), .A2(G28), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n902), .B(KEYINPUT120), .ZN(n906) );
  XOR2_X1 U998 ( .A(G27), .B(n903), .Z(n904) );
  XNOR2_X1 U999 ( .A(KEYINPUT121), .B(n904), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(n906), .A2(n905), .ZN(n907) );
  NAND2_X1 U1001 ( .A1(n908), .A2(n907), .ZN(n911) );
  XNOR2_X1 U1002 ( .A(G32), .B(n909), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1004 ( .A(n912), .B(KEYINPUT53), .ZN(n913) );
  NOR2_X1 U1005 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1006 ( .A(KEYINPUT122), .B(n915), .Z(n916) );
  NOR2_X1 U1007 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1008 ( .A1(G29), .A2(n918), .ZN(n919) );
  XNOR2_X1 U1009 ( .A(n919), .B(KEYINPUT55), .ZN(n950) );
  XOR2_X1 U1010 ( .A(G2084), .B(G160), .Z(n920) );
  NOR2_X1 U1011 ( .A1(n1007), .A2(n920), .ZN(n921) );
  NAND2_X1 U1012 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n944) );
  NAND2_X1 U1014 ( .A1(G103), .A2(n573), .ZN(n926) );
  NAND2_X1 U1015 ( .A1(G139), .A2(n1000), .ZN(n925) );
  NAND2_X1 U1016 ( .A1(n926), .A2(n925), .ZN(n932) );
  NAND2_X1 U1017 ( .A1(G115), .A2(n995), .ZN(n928) );
  NAND2_X1 U1018 ( .A1(G127), .A2(n996), .ZN(n927) );
  NAND2_X1 U1019 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1020 ( .A(KEYINPUT47), .B(n929), .Z(n930) );
  XNOR2_X1 U1021 ( .A(KEYINPUT116), .B(n930), .ZN(n931) );
  NOR2_X1 U1022 ( .A1(n932), .A2(n931), .ZN(n1017) );
  XOR2_X1 U1023 ( .A(G2072), .B(n1017), .Z(n934) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(n935), .B(KEYINPUT50), .ZN(n937) );
  NAND2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n942) );
  XOR2_X1 U1028 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1029 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(n940), .B(KEYINPUT51), .ZN(n941) );
  NOR2_X1 U1031 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1032 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1033 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1034 ( .A(KEYINPUT52), .B(n947), .Z(n948) );
  NAND2_X1 U1035 ( .A1(G29), .A2(n948), .ZN(n949) );
  NAND2_X1 U1036 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1037 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1038 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1039 ( .A(KEYINPUT62), .B(n955), .Z(G311) );
  XNOR2_X1 U1040 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1041 ( .A(G132), .ZN(G219) );
  INV_X1 U1042 ( .A(G120), .ZN(G236) );
  INV_X1 U1043 ( .A(G96), .ZN(G221) );
  INV_X1 U1044 ( .A(G82), .ZN(G220) );
  INV_X1 U1045 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1046 ( .A1(n957), .A2(n956), .ZN(G325) );
  INV_X1 U1047 ( .A(G325), .ZN(G261) );
  NAND2_X1 U1048 ( .A1(n959), .A2(n958), .ZN(n961) );
  XOR2_X1 U1049 ( .A(n961), .B(n960), .Z(G145) );
  XNOR2_X1 U1050 ( .A(G1348), .B(G2454), .ZN(n962) );
  XNOR2_X1 U1051 ( .A(n962), .B(G2430), .ZN(n963) );
  XNOR2_X1 U1052 ( .A(n963), .B(G1341), .ZN(n969) );
  XOR2_X1 U1053 ( .A(G2443), .B(G2427), .Z(n965) );
  XNOR2_X1 U1054 ( .A(G2438), .B(G2446), .ZN(n964) );
  XNOR2_X1 U1055 ( .A(n965), .B(n964), .ZN(n967) );
  XOR2_X1 U1056 ( .A(G2451), .B(G2435), .Z(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(n969), .B(n968), .ZN(n970) );
  NAND2_X1 U1059 ( .A1(n970), .A2(G14), .ZN(n971) );
  XNOR2_X1 U1060 ( .A(KEYINPUT111), .B(n971), .ZN(G401) );
  INV_X1 U1061 ( .A(n972), .ZN(G319) );
  XOR2_X1 U1062 ( .A(G2678), .B(G2067), .Z(n974) );
  XNOR2_X1 U1063 ( .A(G2084), .B(G2078), .ZN(n973) );
  XNOR2_X1 U1064 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1065 ( .A(n975), .B(KEYINPUT42), .Z(n977) );
  XNOR2_X1 U1066 ( .A(G2072), .B(KEYINPUT113), .ZN(n976) );
  XNOR2_X1 U1067 ( .A(n977), .B(n976), .ZN(n982) );
  XNOR2_X1 U1068 ( .A(n978), .B(G2096), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G2090), .B(KEYINPUT43), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n980), .B(n979), .ZN(n981) );
  XOR2_X1 U1071 ( .A(n982), .B(n981), .Z(G227) );
  XNOR2_X1 U1072 ( .A(G1976), .B(KEYINPUT41), .ZN(n994) );
  XOR2_X1 U1073 ( .A(G1986), .B(G1981), .Z(n984) );
  XNOR2_X1 U1074 ( .A(G1966), .B(G1956), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n984), .B(n983), .ZN(n989) );
  XOR2_X1 U1076 ( .A(G2474), .B(KEYINPUT114), .Z(n987) );
  XOR2_X1 U1077 ( .A(n985), .B(G1991), .Z(n986) );
  XNOR2_X1 U1078 ( .A(n987), .B(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(n989), .B(n988), .Z(n992) );
  XOR2_X1 U1080 ( .A(n990), .B(G1971), .Z(n991) );
  XNOR2_X1 U1081 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(n994), .B(n993), .ZN(G229) );
  NAND2_X1 U1083 ( .A1(G118), .A2(n995), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(G130), .A2(n996), .ZN(n997) );
  NAND2_X1 U1085 ( .A1(n998), .A2(n997), .ZN(n1005) );
  NAND2_X1 U1086 ( .A1(n573), .A2(G106), .ZN(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT115), .B(n999), .Z(n1002) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(G142), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(KEYINPUT45), .B(n1003), .Z(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1007), .B(n1006), .ZN(n1016) );
  XNOR2_X1 U1093 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G164), .B(KEYINPUT46), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(n1009), .B(n1008), .ZN(n1010) );
  XNOR2_X1 U1096 ( .A(G162), .B(n1010), .ZN(n1014) );
  XOR2_X1 U1097 ( .A(n1012), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1098 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(n1016), .B(n1015), .ZN(n1021) );
  XNOR2_X1 U1100 ( .A(G160), .B(n1017), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(n1019), .B(n1018), .ZN(n1020) );
  XOR2_X1 U1102 ( .A(n1021), .B(n1020), .Z(n1022) );
  NOR2_X1 U1103 ( .A1(G37), .A2(n1022), .ZN(G395) );
  XOR2_X1 U1104 ( .A(n1023), .B(G286), .Z(n1026) );
  XOR2_X1 U1105 ( .A(G301), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1106 ( .A(n1026), .B(n1025), .ZN(n1028) );
  XNOR2_X1 U1107 ( .A(n1028), .B(n1027), .ZN(n1029) );
  NOR2_X1 U1108 ( .A1(G37), .A2(n1029), .ZN(G397) );
  NOR2_X1 U1109 ( .A1(G227), .A2(G229), .ZN(n1030) );
  XOR2_X1 U1110 ( .A(KEYINPUT49), .B(n1030), .Z(n1031) );
  NAND2_X1 U1111 ( .A1(G319), .A2(n1031), .ZN(n1032) );
  NOR2_X1 U1112 ( .A1(G401), .A2(n1032), .ZN(n1033) );
  XNOR2_X1 U1113 ( .A(KEYINPUT118), .B(n1033), .ZN(n1035) );
  NOR2_X1 U1114 ( .A1(G395), .A2(G397), .ZN(n1034) );
  NAND2_X1 U1115 ( .A1(n1035), .A2(n1034), .ZN(G225) );
  INV_X1 U1116 ( .A(G225), .ZN(G308) );
  INV_X1 U1117 ( .A(G303), .ZN(G166) );
  INV_X1 U1118 ( .A(G108), .ZN(G238) );
endmodule

