

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589;

  INV_X1 U324 ( .A(n553), .ZN(n568) );
  NOR2_X2 U325 ( .A1(n457), .A2(n557), .ZN(n458) );
  XOR2_X1 U326 ( .A(G92GAT), .B(G85GAT), .Z(n385) );
  XNOR2_X1 U327 ( .A(n363), .B(n362), .ZN(n368) );
  NOR2_X1 U328 ( .A1(n536), .A2(n452), .ZN(n576) );
  XOR2_X1 U329 ( .A(G155GAT), .B(G211GAT), .Z(n292) );
  AND2_X1 U330 ( .A1(G231GAT), .A2(G233GAT), .ZN(n293) );
  NOR2_X1 U331 ( .A1(n405), .A2(n404), .ZN(n406) );
  XNOR2_X1 U332 ( .A(KEYINPUT47), .B(KEYINPUT107), .ZN(n399) );
  XNOR2_X1 U333 ( .A(n400), .B(n399), .ZN(n409) );
  XNOR2_X1 U334 ( .A(KEYINPUT71), .B(KEYINPUT31), .ZN(n362) );
  XNOR2_X1 U335 ( .A(n356), .B(n293), .ZN(n327) );
  XNOR2_X1 U336 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U337 ( .A(n373), .B(n385), .ZN(n374) );
  XNOR2_X1 U338 ( .A(n375), .B(n374), .ZN(n377) );
  XNOR2_X1 U339 ( .A(n344), .B(n343), .ZN(n575) );
  XOR2_X1 U340 ( .A(n469), .B(KEYINPUT28), .Z(n538) );
  XNOR2_X1 U341 ( .A(n459), .B(G211GAT), .ZN(n460) );
  XNOR2_X1 U342 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U343 ( .A(n461), .B(n460), .ZN(G1354GAT) );
  XNOR2_X1 U344 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(G43GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n294), .B(G113GAT), .ZN(n358) );
  XOR2_X1 U347 ( .A(n358), .B(KEYINPUT85), .Z(n296) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n299) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G134GAT), .Z(n392) );
  XNOR2_X1 U351 ( .A(n392), .B(G176GAT), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n297), .B(KEYINPUT20), .ZN(n298) );
  XOR2_X1 U353 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U354 ( .A(G127GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U355 ( .A(KEYINPUT82), .B(KEYINPUT83), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n428) );
  XNOR2_X1 U357 ( .A(G99GAT), .B(G71GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n302), .B(G120GAT), .ZN(n372) );
  XNOR2_X1 U359 ( .A(n428), .B(n372), .ZN(n303) );
  XNOR2_X1 U360 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U361 ( .A(KEYINPUT84), .B(G183GAT), .Z(n306) );
  XNOR2_X1 U362 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U364 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U365 ( .A(n308), .B(n307), .ZN(n419) );
  XOR2_X1 U366 ( .A(n309), .B(n419), .Z(n504) );
  INV_X1 U367 ( .A(n504), .ZN(n536) );
  XOR2_X1 U368 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n311) );
  XNOR2_X1 U369 ( .A(G50GAT), .B(KEYINPUT87), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n325) );
  XOR2_X1 U371 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n313) );
  NAND2_X1 U372 ( .A1(G228GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U374 ( .A(n314), .B(KEYINPUT24), .Z(n319) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n316) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(G204GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n363) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n317), .B(G211GAT), .ZN(n412) );
  XNOR2_X1 U380 ( .A(n363), .B(n412), .ZN(n318) );
  XNOR2_X1 U381 ( .A(n319), .B(n318), .ZN(n321) );
  XNOR2_X1 U382 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n320), .B(KEYINPUT2), .ZN(n441) );
  XOR2_X1 U384 ( .A(n321), .B(n441), .Z(n323) );
  XOR2_X1 U385 ( .A(G141GAT), .B(G22GAT), .Z(n359) );
  XOR2_X1 U386 ( .A(G218GAT), .B(G162GAT), .Z(n384) );
  XNOR2_X1 U387 ( .A(n359), .B(n384), .ZN(n322) );
  XNOR2_X1 U388 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U389 ( .A(n325), .B(n324), .Z(n469) );
  INV_X1 U390 ( .A(KEYINPUT64), .ZN(n450) );
  XNOR2_X1 U391 ( .A(G22GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U392 ( .A(n292), .B(n326), .ZN(n328) );
  XOR2_X1 U393 ( .A(G8GAT), .B(G1GAT), .Z(n356) );
  XOR2_X1 U394 ( .A(n329), .B(KEYINPUT78), .Z(n332) );
  XNOR2_X1 U395 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n330), .B(KEYINPUT13), .ZN(n371) );
  XNOR2_X1 U397 ( .A(n371), .B(KEYINPUT79), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U399 ( .A(G71GAT), .B(G127GAT), .Z(n334) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(G183GAT), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U402 ( .A(n336), .B(n335), .Z(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT75), .B(KEYINPUT15), .Z(n338) );
  XNOR2_X1 U404 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n337) );
  XNOR2_X1 U405 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U406 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n340) );
  XNOR2_X1 U407 ( .A(KEYINPUT74), .B(G64GAT), .ZN(n339) );
  XNOR2_X1 U408 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U410 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n346) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U412 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U413 ( .A(n347), .B(KEYINPUT66), .Z(n355) );
  XOR2_X1 U414 ( .A(KEYINPUT7), .B(G50GAT), .Z(n349) );
  XNOR2_X1 U415 ( .A(G36GAT), .B(G29GAT), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U417 ( .A(KEYINPUT8), .B(n350), .Z(n393) );
  XOR2_X1 U418 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n352) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G197GAT), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n393), .B(n353), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n357) );
  XOR2_X1 U423 ( .A(n357), .B(n356), .Z(n361) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n578) );
  INV_X1 U426 ( .A(n368), .ZN(n366) );
  XOR2_X1 U427 ( .A(G176GAT), .B(G64GAT), .Z(n411) );
  XNOR2_X1 U428 ( .A(n411), .B(KEYINPUT32), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(KEYINPUT33), .ZN(n367) );
  INV_X1 U430 ( .A(n367), .ZN(n365) );
  NAND2_X1 U431 ( .A1(n366), .A2(n365), .ZN(n370) );
  NAND2_X1 U432 ( .A1(n368), .A2(n367), .ZN(n369) );
  NAND2_X1 U433 ( .A1(n370), .A2(n369), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n372), .B(n371), .ZN(n373) );
  NAND2_X1 U435 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n404) );
  XOR2_X1 U437 ( .A(KEYINPUT41), .B(n404), .Z(n561) );
  AND2_X1 U438 ( .A1(n578), .A2(n561), .ZN(n380) );
  XOR2_X1 U439 ( .A(KEYINPUT46), .B(KEYINPUT106), .Z(n378) );
  XNOR2_X1 U440 ( .A(KEYINPUT105), .B(n378), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  NOR2_X1 U442 ( .A1(n575), .A2(n381), .ZN(n398) );
  XOR2_X1 U443 ( .A(KEYINPUT72), .B(KEYINPUT9), .Z(n383) );
  XNOR2_X1 U444 ( .A(KEYINPUT11), .B(KEYINPUT73), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n397) );
  XOR2_X1 U446 ( .A(n385), .B(n384), .Z(n387) );
  NAND2_X1 U447 ( .A1(G232GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U449 ( .A(KEYINPUT10), .B(G106GAT), .Z(n389) );
  XNOR2_X1 U450 ( .A(G43GAT), .B(G99GAT), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U452 ( .A(n391), .B(n390), .Z(n395) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X2 U455 ( .A(n397), .B(n396), .Z(n553) );
  NAND2_X1 U456 ( .A1(n398), .A2(n553), .ZN(n400) );
  XNOR2_X1 U457 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n403) );
  XNOR2_X1 U458 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n401) );
  XNOR2_X1 U459 ( .A(n401), .B(n568), .ZN(n587) );
  NAND2_X1 U460 ( .A1(n575), .A2(n587), .ZN(n402) );
  XOR2_X1 U461 ( .A(n403), .B(n402), .Z(n405) );
  XOR2_X1 U462 ( .A(n578), .B(KEYINPUT69), .Z(n573) );
  INV_X1 U463 ( .A(n573), .ZN(n539) );
  NAND2_X1 U464 ( .A1(n406), .A2(n539), .ZN(n407) );
  XNOR2_X1 U465 ( .A(KEYINPUT108), .B(n407), .ZN(n408) );
  NAND2_X1 U466 ( .A1(n409), .A2(n408), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n410), .B(KEYINPUT48), .ZN(n533) );
  XOR2_X1 U468 ( .A(n412), .B(n411), .Z(n414) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT74), .B(KEYINPUT92), .Z(n416) );
  XNOR2_X1 U472 ( .A(G8GAT), .B(G204GAT), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U474 ( .A(n418), .B(n417), .Z(n425) );
  INV_X1 U475 ( .A(n419), .ZN(n423) );
  XOR2_X1 U476 ( .A(G92GAT), .B(G218GAT), .Z(n421) );
  XNOR2_X1 U477 ( .A(G36GAT), .B(G190GAT), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n502) );
  NAND2_X1 U481 ( .A1(n533), .A2(n502), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n448) );
  XOR2_X1 U484 ( .A(G85GAT), .B(n428), .Z(n430) );
  NAND2_X1 U485 ( .A1(G225GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(G29GAT), .B(n431), .ZN(n447) );
  XOR2_X1 U488 ( .A(G57GAT), .B(G120GAT), .Z(n433) );
  XNOR2_X1 U489 ( .A(G113GAT), .B(G1GAT), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U491 ( .A(G162GAT), .B(G148GAT), .Z(n435) );
  XNOR2_X1 U492 ( .A(G141GAT), .B(G134GAT), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n445) );
  XOR2_X1 U495 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n439) );
  XNOR2_X1 U497 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n498) );
  NOR2_X1 U503 ( .A1(n448), .A2(n498), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n457) );
  NOR2_X1 U505 ( .A1(n469), .A2(n457), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  NAND2_X1 U507 ( .A1(n576), .A2(n561), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n453) );
  XNOR2_X1 U509 ( .A(n453), .B(G176GAT), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  NAND2_X1 U511 ( .A1(n469), .A2(n536), .ZN(n456) );
  XNOR2_X1 U512 ( .A(n456), .B(KEYINPUT26), .ZN(n557) );
  XOR2_X1 U513 ( .A(KEYINPUT123), .B(n458), .Z(n586) );
  NAND2_X1 U514 ( .A1(n586), .A2(n575), .ZN(n461) );
  XOR2_X1 U515 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n459) );
  NAND2_X1 U516 ( .A1(n576), .A2(n568), .ZN(n465) );
  XOR2_X1 U517 ( .A(KEYINPUT58), .B(KEYINPUT122), .Z(n463) );
  INV_X1 U518 ( .A(G190GAT), .ZN(n462) );
  INV_X1 U519 ( .A(n498), .ZN(n522) );
  NOR2_X1 U520 ( .A1(n404), .A2(n539), .ZN(n496) );
  XOR2_X1 U521 ( .A(n502), .B(KEYINPUT27), .Z(n472) );
  NOR2_X1 U522 ( .A1(n472), .A2(n522), .ZN(n534) );
  NAND2_X1 U523 ( .A1(n534), .A2(n538), .ZN(n467) );
  XOR2_X1 U524 ( .A(n536), .B(KEYINPUT86), .Z(n466) );
  NOR2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n477) );
  INV_X1 U526 ( .A(n502), .ZN(n525) );
  NOR2_X1 U527 ( .A1(n536), .A2(n525), .ZN(n468) );
  NOR2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U529 ( .A(n470), .B(KEYINPUT93), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT25), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n557), .A2(n472), .ZN(n473) );
  NOR2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n498), .A2(n475), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n493) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n479) );
  NAND2_X1 U536 ( .A1(n575), .A2(n553), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n480), .B(KEYINPUT80), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n493), .A2(n481), .ZN(n511) );
  NAND2_X1 U540 ( .A1(n496), .A2(n511), .ZN(n490) );
  NOR2_X1 U541 ( .A1(n522), .A2(n490), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(n482), .Z(n483) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n525), .A2(n490), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n486), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n536), .A2(n490), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT96), .B(KEYINPUT35), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(n489), .ZN(G1326GAT) );
  NOR2_X1 U552 ( .A1(n538), .A2(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(G22GAT), .B(KEYINPUT97), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT99), .B(KEYINPUT39), .Z(n500) );
  NOR2_X1 U556 ( .A1(n575), .A2(n493), .ZN(n494) );
  NAND2_X1 U557 ( .A1(n494), .A2(n587), .ZN(n495) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n495), .ZN(n521) );
  NAND2_X1 U559 ( .A1(n521), .A2(n496), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT38), .B(n497), .Z(n507) );
  NAND2_X1 U561 ( .A1(n498), .A2(n507), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U563 ( .A(G29GAT), .B(n501), .Z(G1328GAT) );
  NAND2_X1 U564 ( .A1(n507), .A2(n502), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n504), .A2(n507), .ZN(n505) );
  XNOR2_X1 U567 ( .A(KEYINPUT40), .B(n505), .ZN(n506) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  XNOR2_X1 U569 ( .A(G50GAT), .B(KEYINPUT100), .ZN(n510) );
  INV_X1 U570 ( .A(n538), .ZN(n508) );
  NAND2_X1 U571 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1331GAT) );
  INV_X1 U573 ( .A(n561), .ZN(n541) );
  NOR2_X1 U574 ( .A1(n578), .A2(n541), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n520), .A2(n511), .ZN(n517) );
  NOR2_X1 U576 ( .A1(n522), .A2(n517), .ZN(n512) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n525), .A2(n517), .ZN(n514) );
  XOR2_X1 U580 ( .A(G64GAT), .B(n514), .Z(G1333GAT) );
  NOR2_X1 U581 ( .A1(n536), .A2(n517), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G71GAT), .B(KEYINPUT101), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(G1334GAT) );
  NOR2_X1 U584 ( .A1(n538), .A2(n517), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n530) );
  NOR2_X1 U588 ( .A1(n522), .A2(n530), .ZN(n523) );
  XOR2_X1 U589 ( .A(G85GAT), .B(n523), .Z(n524) );
  XNOR2_X1 U590 ( .A(KEYINPUT102), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U591 ( .A1(n525), .A2(n530), .ZN(n526) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n536), .A2(n530), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NOR2_X1 U597 ( .A1(n538), .A2(n530), .ZN(n531) );
  XOR2_X1 U598 ( .A(KEYINPUT44), .B(n531), .Z(n532) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U601 ( .A(KEYINPUT109), .B(n535), .Z(n558) );
  NOR2_X1 U602 ( .A1(n536), .A2(n558), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n538), .A2(n537), .ZN(n552) );
  NOR2_X1 U604 ( .A1(n539), .A2(n552), .ZN(n540) );
  XOR2_X1 U605 ( .A(G113GAT), .B(n540), .Z(G1340GAT) );
  NOR2_X1 U606 ( .A1(n552), .A2(n541), .ZN(n545) );
  XOR2_X1 U607 ( .A(KEYINPUT110), .B(KEYINPUT49), .Z(n543) );
  XNOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT111), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(KEYINPUT113), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(n550) );
  INV_X1 U614 ( .A(n575), .ZN(n548) );
  NOR2_X1 U615 ( .A1(n548), .A2(n552), .ZN(n549) );
  XOR2_X1 U616 ( .A(n550), .B(n549), .Z(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT112), .B(n551), .ZN(G1342GAT) );
  NOR2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U619 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U621 ( .A(G134GAT), .B(n556), .Z(G1343GAT) );
  NOR2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n559), .B(KEYINPUT116), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n578), .A2(n569), .ZN(n560) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n560), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n563) );
  NAND2_X1 U627 ( .A1(n561), .A2(n569), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U629 ( .A(G148GAT), .B(KEYINPUT53), .Z(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U631 ( .A1(n569), .A2(n575), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(KEYINPUT118), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G155GAT), .B(n567), .ZN(G1346GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n571) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G162GAT), .B(n572), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n576), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n580) );
  NAND2_X1 U643 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n583) );
  NAND2_X1 U647 ( .A1(n586), .A2(n404), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n585) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT124), .Z(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(KEYINPUT62), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

