

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775;

  NAND2_X1 U374 ( .A1(n741), .A2(n641), .ZN(n735) );
  NAND2_X1 U375 ( .A1(n578), .A2(n577), .ZN(n719) );
  BUF_X1 U376 ( .A(G107), .Z(n352) );
  XNOR2_X1 U377 ( .A(n751), .B(KEYINPUT69), .ZN(n507) );
  XNOR2_X2 U378 ( .A(n513), .B(n512), .ZN(n540) );
  INV_X2 U379 ( .A(G953), .ZN(n767) );
  AND2_X2 U380 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X2 U381 ( .A1(n402), .A2(n400), .ZN(n401) );
  XNOR2_X2 U382 ( .A(n401), .B(KEYINPUT103), .ZN(n613) );
  XNOR2_X1 U383 ( .A(n439), .B(n410), .ZN(n508) );
  AND2_X1 U384 ( .A1(n735), .A2(G472), .ZN(n374) );
  AND2_X1 U385 ( .A1(n775), .A2(n622), .ZN(n631) );
  OR2_X1 U386 ( .A1(n678), .A2(n580), .ZN(n528) );
  OR2_X1 U387 ( .A1(n562), .A2(n661), .ZN(n667) );
  OR2_X1 U388 ( .A1(G902), .A2(n739), .ZN(n498) );
  XNOR2_X1 U389 ( .A(G143), .B(G128), .ZN(n493) );
  INV_X1 U390 ( .A(n701), .ZN(n392) );
  BUF_X1 U391 ( .A(n604), .Z(n609) );
  NOR2_X2 U392 ( .A1(n540), .A2(n661), .ZN(n363) );
  XNOR2_X2 U393 ( .A(n441), .B(n440), .ZN(n751) );
  XNOR2_X2 U394 ( .A(KEYINPUT87), .B(G107), .ZN(n441) );
  OR2_X2 U395 ( .A1(n702), .A2(n688), .ZN(n513) );
  XNOR2_X2 U396 ( .A(n555), .B(KEYINPUT22), .ZN(n620) );
  XNOR2_X2 U397 ( .A(n552), .B(KEYINPUT0), .ZN(n604) );
  XNOR2_X1 U398 ( .A(G122), .B(G104), .ZN(n506) );
  XNOR2_X1 U399 ( .A(n508), .B(n431), .ZN(n693) );
  NAND2_X1 U400 ( .A1(n701), .A2(n358), .ZN(n396) );
  AND2_X2 U401 ( .A1(n737), .A2(n735), .ZN(n701) );
  INV_X1 U402 ( .A(KEYINPUT46), .ZN(n570) );
  INV_X1 U403 ( .A(KEYINPUT80), .ZN(n628) );
  NOR2_X1 U404 ( .A1(G953), .A2(G237), .ZN(n477) );
  INV_X1 U405 ( .A(G237), .ZN(n433) );
  XNOR2_X1 U406 ( .A(n748), .B(n504), .ZN(n366) );
  OR2_X1 U407 ( .A1(n698), .A2(G902), .ZN(n461) );
  OR2_X1 U408 ( .A1(n693), .A2(G902), .ZN(n432) );
  AND2_X1 U409 ( .A1(n396), .A2(n353), .ZN(n387) );
  XNOR2_X1 U410 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U411 ( .A(KEYINPUT77), .ZN(n378) );
  XNOR2_X1 U412 ( .A(G146), .B(G125), .ZN(n501) );
  XNOR2_X1 U413 ( .A(n571), .B(n570), .ZN(n589) );
  OR2_X1 U414 ( .A1(n633), .A2(n632), .ZN(n423) );
  AND2_X1 U415 ( .A1(G234), .A2(n767), .ZN(n448) );
  XNOR2_X1 U416 ( .A(G131), .B(G140), .ZN(n471) );
  XNOR2_X1 U417 ( .A(G143), .B(G113), .ZN(n478) );
  XNOR2_X1 U418 ( .A(n501), .B(KEYINPUT10), .ZN(n760) );
  AND2_X1 U419 ( .A1(n687), .A2(n385), .ZN(n384) );
  NAND2_X1 U420 ( .A1(n509), .A2(KEYINPUT76), .ZN(n385) );
  XNOR2_X1 U421 ( .A(G137), .B(G140), .ZN(n446) );
  XNOR2_X1 U422 ( .A(G134), .B(G131), .ZN(n761) );
  XNOR2_X1 U423 ( .A(n493), .B(KEYINPUT4), .ZN(n763) );
  INV_X1 U424 ( .A(n679), .ZN(n407) );
  INV_X1 U425 ( .A(KEYINPUT34), .ZN(n416) );
  XNOR2_X1 U426 ( .A(n511), .B(KEYINPUT74), .ZN(n512) );
  XNOR2_X1 U427 ( .A(G119), .B(G113), .ZN(n424) );
  INV_X1 U428 ( .A(G110), .ZN(n440) );
  XNOR2_X1 U429 ( .A(G128), .B(G119), .ZN(n453) );
  XNOR2_X1 U430 ( .A(n352), .B(G122), .ZN(n491) );
  INV_X1 U431 ( .A(G104), .ZN(n434) );
  XNOR2_X1 U432 ( .A(n763), .B(G101), .ZN(n439) );
  NOR2_X1 U433 ( .A1(n395), .A2(n740), .ZN(n394) );
  NOR2_X1 U434 ( .A1(n399), .A2(G210), .ZN(n395) );
  AND2_X1 U435 ( .A1(G234), .A2(G237), .ZN(n469) );
  INV_X1 U436 ( .A(KEYINPUT75), .ZN(n637) );
  XNOR2_X1 U437 ( .A(n411), .B(KEYINPUT71), .ZN(n563) );
  NAND2_X1 U438 ( .A1(n413), .A2(n412), .ZN(n411) );
  AND2_X1 U439 ( .A1(n650), .A2(n354), .ZN(n412) );
  XNOR2_X1 U440 ( .A(n363), .B(n362), .ZN(n582) );
  INV_X1 U441 ( .A(KEYINPUT19), .ZN(n362) );
  XNOR2_X1 U442 ( .A(n486), .B(n485), .ZN(n578) );
  XNOR2_X1 U443 ( .A(n484), .B(G475), .ZN(n485) );
  XNOR2_X1 U444 ( .A(n568), .B(n567), .ZN(n684) );
  INV_X1 U445 ( .A(KEYINPUT40), .ZN(n567) );
  NOR2_X1 U446 ( .A1(n593), .A2(n719), .ZN(n568) );
  OR2_X1 U447 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X2 U448 ( .A1(n620), .A2(n561), .ZN(n400) );
  AND2_X1 U449 ( .A1(n372), .A2(n398), .ZN(n697) );
  XNOR2_X1 U450 ( .A(n368), .B(n376), .ZN(n375) );
  INV_X1 U451 ( .A(n739), .ZN(n376) );
  NAND2_X1 U452 ( .A1(n701), .A2(G478), .ZN(n368) );
  XNOR2_X1 U453 ( .A(n369), .B(n361), .ZN(G60) );
  NAND2_X1 U454 ( .A1(n370), .A2(n398), .ZN(n369) );
  XNOR2_X1 U455 ( .A(n371), .B(n357), .ZN(n370) );
  NAND2_X1 U456 ( .A1(n387), .A2(n386), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n392), .A2(n704), .ZN(n386) );
  NAND2_X1 U458 ( .A1(n377), .A2(n355), .ZN(n682) );
  AND2_X1 U459 ( .A1(n394), .A2(KEYINPUT56), .ZN(n353) );
  AND2_X1 U460 ( .A1(n409), .A2(n521), .ZN(n354) );
  AND2_X1 U461 ( .A1(n422), .A2(n767), .ZN(n355) );
  XOR2_X1 U462 ( .A(n690), .B(KEYINPUT65), .Z(n356) );
  XOR2_X1 U463 ( .A(n738), .B(n420), .Z(n357) );
  AND2_X1 U464 ( .A1(n399), .A2(G210), .ZN(n358) );
  AND2_X1 U465 ( .A1(n704), .A2(n397), .ZN(n359) );
  AND2_X1 U466 ( .A1(n356), .A2(n383), .ZN(n360) );
  XNOR2_X1 U467 ( .A(KEYINPUT60), .B(KEYINPUT123), .ZN(n361) );
  AND2_X1 U468 ( .A1(n695), .A2(G953), .ZN(n740) );
  INV_X1 U469 ( .A(n740), .ZN(n398) );
  INV_X1 U470 ( .A(KEYINPUT56), .ZN(n397) );
  NAND2_X1 U471 ( .A1(n613), .A2(n611), .ZN(n612) );
  NAND2_X1 U472 ( .A1(n415), .A2(n384), .ZN(n382) );
  NAND2_X1 U473 ( .A1(n364), .A2(n416), .ZN(n406) );
  NAND2_X1 U474 ( .A1(n408), .A2(n407), .ZN(n364) );
  AND2_X1 U475 ( .A1(n375), .A2(n398), .ZN(G63) );
  NAND2_X1 U476 ( .A1(n634), .A2(n423), .ZN(n635) );
  XNOR2_X1 U477 ( .A(n365), .B(n508), .ZN(n702) );
  XNOR2_X1 U478 ( .A(n367), .B(n366), .ZN(n365) );
  XNOR2_X1 U479 ( .A(n507), .B(n505), .ZN(n367) );
  NAND2_X2 U480 ( .A1(n380), .A2(n382), .ZN(n737) );
  NAND2_X1 U481 ( .A1(n736), .A2(n737), .ZN(n371) );
  XNOR2_X1 U482 ( .A(n373), .B(n694), .ZN(n372) );
  NAND2_X1 U483 ( .A1(n737), .A2(n374), .ZN(n373) );
  NAND2_X1 U484 ( .A1(n642), .A2(n735), .ZN(n379) );
  AND2_X2 U485 ( .A1(n381), .A2(n360), .ZN(n380) );
  NAND2_X1 U486 ( .A1(n685), .A2(n686), .ZN(n381) );
  NAND2_X2 U487 ( .A1(n639), .A2(n766), .ZN(n685) );
  NAND2_X1 U488 ( .A1(n384), .A2(n686), .ZN(n383) );
  NAND2_X1 U489 ( .A1(n396), .A2(n394), .ZN(n393) );
  NAND2_X1 U490 ( .A1(n389), .A2(n388), .ZN(G51) );
  NAND2_X1 U491 ( .A1(n392), .A2(n359), .ZN(n390) );
  NAND2_X1 U492 ( .A1(n393), .A2(n397), .ZN(n391) );
  INV_X1 U493 ( .A(n704), .ZN(n399) );
  XNOR2_X1 U494 ( .A(n400), .B(G101), .ZN(G3) );
  NAND2_X1 U495 ( .A1(n403), .A2(n610), .ZN(n402) );
  NAND2_X1 U496 ( .A1(n722), .A2(n707), .ZN(n403) );
  NAND2_X1 U497 ( .A1(n406), .A2(n404), .ZN(n418) );
  NAND2_X1 U498 ( .A1(n405), .A2(n407), .ZN(n404) );
  NOR2_X1 U499 ( .A1(n609), .A2(n416), .ZN(n405) );
  INV_X1 U500 ( .A(n609), .ZN(n408) );
  AND2_X1 U501 ( .A1(n650), .A2(n409), .ZN(n607) );
  XNOR2_X2 U502 ( .A(n409), .B(n536), .ZN(n651) );
  NAND2_X1 U503 ( .A1(n525), .A2(n409), .ZN(n580) );
  XNOR2_X2 U504 ( .A(n445), .B(G469), .ZN(n409) );
  INV_X1 U505 ( .A(n749), .ZN(n410) );
  XNOR2_X1 U506 ( .A(n414), .B(KEYINPUT30), .ZN(n413) );
  NOR2_X1 U507 ( .A1(n648), .A2(n661), .ZN(n414) );
  INV_X1 U508 ( .A(n685), .ZN(n415) );
  XNOR2_X2 U509 ( .A(n417), .B(KEYINPUT35), .ZN(n774) );
  NAND2_X1 U510 ( .A1(n418), .A2(n601), .ZN(n417) );
  BUF_X1 U511 ( .A(n639), .Z(n741) );
  AND2_X1 U512 ( .A1(n553), .A2(n643), .ZN(n419) );
  XNOR2_X1 U513 ( .A(KEYINPUT59), .B(KEYINPUT85), .ZN(n420) );
  NOR2_X1 U514 ( .A1(n725), .A2(n588), .ZN(n421) );
  AND2_X1 U515 ( .A1(n681), .A2(n680), .ZN(n422) );
  AND2_X1 U516 ( .A1(n650), .A2(n651), .ZN(n597) );
  XNOR2_X1 U517 ( .A(n435), .B(n434), .ZN(n436) );
  INV_X1 U518 ( .A(KEYINPUT104), .ZN(n533) );
  XNOR2_X1 U519 ( .A(n424), .B(KEYINPUT3), .ZN(n426) );
  XNOR2_X1 U520 ( .A(G116), .B(KEYINPUT68), .ZN(n425) );
  XNOR2_X1 U521 ( .A(n426), .B(n425), .ZN(n749) );
  NAND2_X1 U522 ( .A1(n477), .A2(G210), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n427), .B(G137), .ZN(n429) );
  XNOR2_X1 U524 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n428) );
  XNOR2_X1 U525 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U526 ( .A(n761), .B(G146), .ZN(n437) );
  XNOR2_X1 U527 ( .A(n430), .B(n437), .ZN(n431) );
  INV_X1 U528 ( .A(G472), .ZN(n691) );
  XNOR2_X2 U529 ( .A(n432), .B(n691), .ZN(n648) );
  INV_X1 U530 ( .A(G902), .ZN(n444) );
  NAND2_X1 U531 ( .A1(n444), .A2(n433), .ZN(n510) );
  AND2_X1 U532 ( .A1(n510), .A2(G214), .ZN(n661) );
  NAND2_X1 U533 ( .A1(G227), .A2(n767), .ZN(n435) );
  XNOR2_X1 U534 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U535 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U536 ( .A(n446), .B(KEYINPUT90), .ZN(n759) );
  XNOR2_X1 U537 ( .A(n507), .B(n759), .ZN(n442) );
  XNOR2_X1 U538 ( .A(n443), .B(n442), .ZN(n731) );
  NAND2_X1 U539 ( .A1(n731), .A2(n444), .ZN(n445) );
  INV_X1 U540 ( .A(n446), .ZN(n447) );
  XNOR2_X1 U541 ( .A(n760), .B(n447), .ZN(n450) );
  XNOR2_X1 U542 ( .A(n448), .B(KEYINPUT8), .ZN(n487) );
  NAND2_X1 U543 ( .A1(n487), .A2(G221), .ZN(n449) );
  XNOR2_X1 U544 ( .A(n450), .B(n449), .ZN(n457) );
  XNOR2_X1 U545 ( .A(G110), .B(KEYINPUT23), .ZN(n452) );
  XNOR2_X1 U546 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n451) );
  XNOR2_X1 U547 ( .A(n452), .B(n451), .ZN(n455) );
  XNOR2_X1 U548 ( .A(n453), .B(KEYINPUT24), .ZN(n454) );
  XNOR2_X1 U549 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U550 ( .A(n457), .B(n456), .ZN(n698) );
  XNOR2_X1 U551 ( .A(G902), .B(KEYINPUT15), .ZN(n509) );
  NAND2_X1 U552 ( .A1(n509), .A2(G234), .ZN(n458) );
  XNOR2_X1 U553 ( .A(n458), .B(KEYINPUT20), .ZN(n462) );
  AND2_X1 U554 ( .A1(n462), .A2(G217), .ZN(n459) );
  XNOR2_X1 U555 ( .A(n459), .B(KEYINPUT25), .ZN(n460) );
  XNOR2_X2 U556 ( .A(n461), .B(n460), .ZN(n520) );
  INV_X1 U557 ( .A(n462), .ZN(n464) );
  INV_X1 U558 ( .A(G221), .ZN(n463) );
  OR2_X1 U559 ( .A1(n464), .A2(n463), .ZN(n466) );
  INV_X1 U560 ( .A(KEYINPUT21), .ZN(n465) );
  XNOR2_X1 U561 ( .A(n466), .B(n465), .ZN(n643) );
  AND2_X1 U562 ( .A1(n520), .A2(n643), .ZN(n650) );
  NAND2_X1 U563 ( .A1(G953), .A2(G902), .ZN(n541) );
  NOR2_X1 U564 ( .A1(G900), .A2(n541), .ZN(n468) );
  NAND2_X1 U565 ( .A1(n767), .A2(G952), .ZN(n543) );
  INV_X1 U566 ( .A(n543), .ZN(n467) );
  OR2_X1 U567 ( .A1(n468), .A2(n467), .ZN(n470) );
  XNOR2_X1 U568 ( .A(KEYINPUT14), .B(n469), .ZN(n676) );
  INV_X1 U569 ( .A(n676), .ZN(n546) );
  AND2_X1 U570 ( .A1(n470), .A2(n546), .ZN(n521) );
  XOR2_X1 U571 ( .A(KEYINPUT94), .B(KEYINPUT12), .Z(n472) );
  XNOR2_X1 U572 ( .A(n472), .B(n471), .ZN(n476) );
  XOR2_X1 U573 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n474) );
  XNOR2_X1 U574 ( .A(KEYINPUT11), .B(KEYINPUT95), .ZN(n473) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U576 ( .A(n476), .B(n475), .Z(n483) );
  NAND2_X1 U577 ( .A1(n477), .A2(G214), .ZN(n479) );
  XNOR2_X1 U578 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U579 ( .A(n480), .B(n506), .ZN(n481) );
  XNOR2_X1 U580 ( .A(n481), .B(n760), .ZN(n482) );
  XNOR2_X1 U581 ( .A(n483), .B(n482), .ZN(n738) );
  NOR2_X1 U582 ( .A1(G902), .A2(n738), .ZN(n486) );
  XNOR2_X1 U583 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n484) );
  XOR2_X1 U584 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n489) );
  NAND2_X1 U585 ( .A1(G217), .A2(n487), .ZN(n488) );
  XNOR2_X1 U586 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U587 ( .A(n490), .B(G134), .Z(n497) );
  XOR2_X1 U588 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n492) );
  XNOR2_X1 U589 ( .A(n492), .B(n491), .ZN(n495) );
  XNOR2_X1 U590 ( .A(n493), .B(G116), .ZN(n494) );
  XNOR2_X1 U591 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U592 ( .A(n497), .B(n496), .ZN(n739) );
  XNOR2_X1 U593 ( .A(G478), .B(n498), .ZN(n529) );
  NAND2_X1 U594 ( .A1(n578), .A2(n529), .ZN(n600) );
  NAND2_X1 U595 ( .A1(n767), .A2(G224), .ZN(n499) );
  XNOR2_X1 U596 ( .A(n499), .B(KEYINPUT18), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n501), .B(n500), .ZN(n505) );
  XNOR2_X1 U598 ( .A(KEYINPUT73), .B(KEYINPUT83), .ZN(n503) );
  XNOR2_X1 U599 ( .A(KEYINPUT17), .B(KEYINPUT72), .ZN(n502) );
  XNOR2_X1 U600 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U601 ( .A(n506), .B(KEYINPUT16), .ZN(n748) );
  INV_X1 U602 ( .A(n509), .ZN(n688) );
  NAND2_X1 U603 ( .A1(n510), .A2(G210), .ZN(n511) );
  BUF_X1 U604 ( .A(n540), .Z(n514) );
  NOR2_X1 U605 ( .A1(n600), .A2(n514), .ZN(n515) );
  NAND2_X1 U606 ( .A1(n563), .A2(n515), .ZN(n586) );
  XNOR2_X1 U607 ( .A(G143), .B(KEYINPUT112), .ZN(n516) );
  XNOR2_X1 U608 ( .A(n586), .B(n516), .ZN(G45) );
  INV_X1 U609 ( .A(KEYINPUT38), .ZN(n517) );
  XNOR2_X1 U610 ( .A(n514), .B(n517), .ZN(n562) );
  OR2_X1 U611 ( .A1(n578), .A2(n529), .ZN(n666) );
  NOR2_X1 U612 ( .A1(n667), .A2(n666), .ZN(n519) );
  XNOR2_X1 U613 ( .A(KEYINPUT106), .B(KEYINPUT41), .ZN(n518) );
  XNOR2_X1 U614 ( .A(n519), .B(n518), .ZN(n678) );
  NAND2_X1 U615 ( .A1(n643), .A2(n521), .ZN(n522) );
  OR2_X1 U616 ( .A1(n520), .A2(n522), .ZN(n530) );
  OR2_X1 U617 ( .A1(n648), .A2(n530), .ZN(n524) );
  INV_X1 U618 ( .A(KEYINPUT28), .ZN(n523) );
  XNOR2_X1 U619 ( .A(n524), .B(n523), .ZN(n525) );
  INV_X1 U620 ( .A(KEYINPUT107), .ZN(n526) );
  XNOR2_X1 U621 ( .A(n526), .B(KEYINPUT42), .ZN(n527) );
  XNOR2_X1 U622 ( .A(n528), .B(n527), .ZN(n569) );
  XNOR2_X1 U623 ( .A(n569), .B(G137), .ZN(G39) );
  INV_X1 U624 ( .A(n529), .ZN(n577) );
  NOR2_X1 U625 ( .A1(n719), .A2(n530), .ZN(n532) );
  XNOR2_X1 U626 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n531) );
  XNOR2_X1 U627 ( .A(n648), .B(n531), .ZN(n616) );
  AND2_X1 U628 ( .A1(n532), .A2(n616), .ZN(n534) );
  XNOR2_X1 U629 ( .A(n534), .B(n533), .ZN(n535) );
  OR2_X1 U630 ( .A1(n535), .A2(n661), .ZN(n572) );
  XNOR2_X1 U631 ( .A(KEYINPUT64), .B(KEYINPUT1), .ZN(n536) );
  NOR2_X1 U632 ( .A1(n572), .A2(n651), .ZN(n538) );
  XNOR2_X1 U633 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n537) );
  XNOR2_X1 U634 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U635 ( .A1(n539), .A2(n514), .ZN(n594) );
  XNOR2_X1 U636 ( .A(n594), .B(G140), .ZN(G42) );
  XNOR2_X1 U637 ( .A(KEYINPUT88), .B(G898), .ZN(n754) );
  NOR2_X1 U638 ( .A1(n541), .A2(n754), .ZN(n547) );
  INV_X1 U639 ( .A(KEYINPUT89), .ZN(n542) );
  NAND2_X1 U640 ( .A1(n547), .A2(n542), .ZN(n544) );
  NAND2_X1 U641 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U642 ( .A1(n545), .A2(n546), .ZN(n550) );
  NAND2_X1 U643 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U644 ( .A1(n548), .A2(KEYINPUT89), .ZN(n549) );
  NAND2_X1 U645 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U646 ( .A1(n582), .A2(n551), .ZN(n552) );
  INV_X1 U647 ( .A(n604), .ZN(n554) );
  INV_X1 U648 ( .A(n666), .ZN(n553) );
  NAND2_X1 U649 ( .A1(n554), .A2(n419), .ZN(n555) );
  INV_X1 U650 ( .A(n620), .ZN(n558) );
  INV_X1 U651 ( .A(n520), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n648), .A2(n559), .ZN(n556) );
  NOR2_X1 U653 ( .A1(n651), .A2(n556), .ZN(n557) );
  NAND2_X1 U654 ( .A1(n558), .A2(n557), .ZN(n622) );
  XNOR2_X1 U655 ( .A(n622), .B(G110), .ZN(G12) );
  OR2_X1 U656 ( .A1(n651), .A2(n559), .ZN(n560) );
  OR2_X1 U657 ( .A1(n560), .A2(n616), .ZN(n561) );
  INV_X1 U658 ( .A(KEYINPUT53), .ZN(n683) );
  INV_X1 U659 ( .A(n562), .ZN(n663) );
  NAND2_X1 U660 ( .A1(n563), .A2(n663), .ZN(n566) );
  INV_X1 U661 ( .A(KEYINPUT70), .ZN(n564) );
  XNOR2_X1 U662 ( .A(n564), .B(KEYINPUT39), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n566), .B(n565), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n684), .A2(n569), .ZN(n571) );
  NOR2_X1 U665 ( .A1(n572), .A2(n514), .ZN(n575) );
  XNOR2_X1 U666 ( .A(KEYINPUT108), .B(KEYINPUT36), .ZN(n573) );
  XNOR2_X1 U667 ( .A(n573), .B(KEYINPUT82), .ZN(n574) );
  XNOR2_X1 U668 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U669 ( .A(n651), .B(KEYINPUT84), .ZN(n618) );
  AND2_X1 U670 ( .A1(n576), .A2(n618), .ZN(n725) );
  OR2_X1 U671 ( .A1(n578), .A2(n577), .ZN(n723) );
  INV_X1 U672 ( .A(KEYINPUT101), .ZN(n579) );
  XNOR2_X1 U673 ( .A(n723), .B(n579), .ZN(n592) );
  AND2_X1 U674 ( .A1(n592), .A2(n719), .ZN(n668) );
  NOR2_X1 U675 ( .A1(n668), .A2(KEYINPUT67), .ZN(n583) );
  INV_X1 U676 ( .A(n580), .ZN(n581) );
  AND2_X1 U677 ( .A1(n582), .A2(n581), .ZN(n716) );
  NAND2_X1 U678 ( .A1(n583), .A2(n716), .ZN(n585) );
  INV_X1 U679 ( .A(KEYINPUT47), .ZN(n584) );
  XNOR2_X1 U680 ( .A(n585), .B(n584), .ZN(n587) );
  NAND2_X1 U681 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U682 ( .A1(n589), .A2(n421), .ZN(n591) );
  INV_X1 U683 ( .A(KEYINPUT48), .ZN(n590) );
  XNOR2_X1 U684 ( .A(n591), .B(n590), .ZN(n596) );
  OR2_X1 U685 ( .A1(n593), .A2(n592), .ZN(n727) );
  AND2_X1 U686 ( .A1(n594), .A2(n727), .ZN(n595) );
  NAND2_X1 U687 ( .A1(n596), .A2(n595), .ZN(n640) );
  XNOR2_X2 U688 ( .A(n640), .B(KEYINPUT79), .ZN(n766) );
  NAND2_X1 U689 ( .A1(n597), .A2(n616), .ZN(n599) );
  INV_X1 U690 ( .A(KEYINPUT33), .ZN(n598) );
  XNOR2_X2 U691 ( .A(n599), .B(n598), .ZN(n679) );
  INV_X1 U692 ( .A(n600), .ZN(n601) );
  NAND2_X1 U693 ( .A1(n774), .A2(KEYINPUT44), .ZN(n611) );
  INV_X1 U694 ( .A(n650), .ZN(n602) );
  NOR2_X1 U695 ( .A1(n648), .A2(n602), .ZN(n603) );
  NAND2_X1 U696 ( .A1(n651), .A2(n603), .ZN(n656) );
  OR2_X2 U697 ( .A1(n604), .A2(n656), .ZN(n606) );
  INV_X1 U698 ( .A(KEYINPUT31), .ZN(n605) );
  XNOR2_X2 U699 ( .A(n606), .B(n605), .ZN(n722) );
  NAND2_X1 U700 ( .A1(n607), .A2(n648), .ZN(n608) );
  OR2_X1 U701 ( .A1(n609), .A2(n608), .ZN(n707) );
  INV_X1 U702 ( .A(n668), .ZN(n610) );
  NAND2_X1 U703 ( .A1(n612), .A2(KEYINPUT81), .ZN(n615) );
  INV_X1 U704 ( .A(KEYINPUT81), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n613), .A2(n623), .ZN(n614) );
  NAND2_X1 U706 ( .A1(n615), .A2(n614), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n616), .A2(n520), .ZN(n617) );
  NAND2_X1 U708 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X2 U709 ( .A(n621), .B(KEYINPUT32), .ZN(n775) );
  NAND2_X1 U710 ( .A1(n774), .A2(n623), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n631), .A2(n624), .ZN(n625) );
  NAND2_X1 U712 ( .A1(n625), .A2(KEYINPUT44), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n629) );
  XNOR2_X1 U714 ( .A(n629), .B(n628), .ZN(n634) );
  OR2_X2 U715 ( .A1(n774), .A2(KEYINPUT44), .ZN(n630) );
  XNOR2_X1 U716 ( .A(n630), .B(KEYINPUT66), .ZN(n633) );
  INV_X1 U717 ( .A(n631), .ZN(n632) );
  XNOR2_X2 U718 ( .A(n635), .B(KEYINPUT45), .ZN(n639) );
  INV_X1 U719 ( .A(KEYINPUT2), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n685), .A2(n636), .ZN(n638) );
  XNOR2_X1 U721 ( .A(n638), .B(n637), .ZN(n642) );
  NOR2_X1 U722 ( .A1(n640), .A2(n636), .ZN(n641) );
  NOR2_X1 U723 ( .A1(n520), .A2(n643), .ZN(n646) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n644) );
  XNOR2_X1 U725 ( .A(n644), .B(KEYINPUT116), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n646), .B(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(KEYINPUT118), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U730 ( .A(n652), .B(KEYINPUT50), .ZN(n653) );
  NOR2_X1 U731 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U732 ( .A(KEYINPUT119), .B(n655), .ZN(n657) );
  NAND2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n658), .B(KEYINPUT51), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n659), .B(KEYINPUT120), .ZN(n660) );
  NOR2_X1 U736 ( .A1(n678), .A2(n660), .ZN(n673) );
  INV_X1 U737 ( .A(n661), .ZN(n662) );
  NOR2_X1 U738 ( .A1(n663), .A2(n662), .ZN(n664) );
  XOR2_X1 U739 ( .A(KEYINPUT121), .B(n664), .Z(n665) );
  NOR2_X1 U740 ( .A1(n666), .A2(n665), .ZN(n670) );
  NOR2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U742 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U743 ( .A1(n671), .A2(n679), .ZN(n672) );
  NOR2_X1 U744 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U745 ( .A(n674), .B(KEYINPUT52), .ZN(n675) );
  NOR2_X1 U746 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U747 ( .A1(G952), .A2(n677), .ZN(n681) );
  OR2_X1 U748 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n683), .B(n682), .ZN(G75) );
  XNOR2_X1 U750 ( .A(n684), .B(G131), .ZN(G33) );
  INV_X1 U751 ( .A(KEYINPUT76), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n688), .A2(n686), .ZN(n687) );
  XNOR2_X1 U753 ( .A(n688), .B(KEYINPUT78), .ZN(n689) );
  NAND2_X1 U754 ( .A1(n689), .A2(KEYINPUT2), .ZN(n690) );
  XNOR2_X1 U755 ( .A(KEYINPUT109), .B(KEYINPUT62), .ZN(n692) );
  XNOR2_X1 U756 ( .A(n693), .B(n692), .ZN(n694) );
  INV_X1 U757 ( .A(G952), .ZN(n695) );
  XOR2_X1 U758 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n696) );
  XNOR2_X1 U759 ( .A(n697), .B(n696), .ZN(G57) );
  NAND2_X1 U760 ( .A1(n701), .A2(G217), .ZN(n699) );
  XNOR2_X1 U761 ( .A(n699), .B(n698), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n700), .A2(n740), .ZN(G66) );
  XOR2_X1 U763 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n703) );
  XNOR2_X1 U764 ( .A(n702), .B(n703), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n707), .A2(n719), .ZN(n705) );
  XOR2_X1 U766 ( .A(KEYINPUT110), .B(n705), .Z(n706) );
  XNOR2_X1 U767 ( .A(G104), .B(n706), .ZN(G6) );
  NOR2_X1 U768 ( .A1(n707), .A2(n723), .ZN(n711) );
  XOR2_X1 U769 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n709) );
  XNOR2_X1 U770 ( .A(n352), .B(KEYINPUT111), .ZN(n708) );
  XNOR2_X1 U771 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U772 ( .A(n711), .B(n710), .ZN(G9) );
  XOR2_X1 U773 ( .A(G128), .B(KEYINPUT29), .Z(n714) );
  INV_X1 U774 ( .A(n723), .ZN(n712) );
  NAND2_X1 U775 ( .A1(n716), .A2(n712), .ZN(n713) );
  XNOR2_X1 U776 ( .A(n714), .B(n713), .ZN(G30) );
  XOR2_X1 U777 ( .A(G146), .B(KEYINPUT113), .Z(n718) );
  INV_X1 U778 ( .A(n719), .ZN(n715) );
  NAND2_X1 U779 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U780 ( .A(n718), .B(n717), .ZN(G48) );
  NOR2_X1 U781 ( .A1(n719), .A2(n722), .ZN(n720) );
  XOR2_X1 U782 ( .A(KEYINPUT114), .B(n720), .Z(n721) );
  XNOR2_X1 U783 ( .A(G113), .B(n721), .ZN(G15) );
  NOR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U785 ( .A(G116), .B(n724), .Z(G18) );
  XNOR2_X1 U786 ( .A(G125), .B(n725), .ZN(n726) );
  XNOR2_X1 U787 ( .A(n726), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U788 ( .A(G134), .B(n727), .Z(n728) );
  XNOR2_X1 U789 ( .A(n728), .B(KEYINPUT115), .ZN(G36) );
  NAND2_X1 U790 ( .A1(n701), .A2(G469), .ZN(n733) );
  XNOR2_X1 U791 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n729) );
  XNOR2_X1 U792 ( .A(n729), .B(KEYINPUT57), .ZN(n730) );
  XNOR2_X1 U793 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U794 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U795 ( .A1(n740), .A2(n734), .ZN(G54) );
  AND2_X1 U796 ( .A1(n735), .A2(G475), .ZN(n736) );
  NAND2_X1 U797 ( .A1(n741), .A2(n767), .ZN(n747) );
  NAND2_X1 U798 ( .A1(G224), .A2(G953), .ZN(n742) );
  XNOR2_X1 U799 ( .A(n742), .B(KEYINPUT61), .ZN(n743) );
  XNOR2_X1 U800 ( .A(n743), .B(KEYINPUT124), .ZN(n744) );
  NAND2_X1 U801 ( .A1(n744), .A2(n754), .ZN(n745) );
  XOR2_X1 U802 ( .A(KEYINPUT125), .B(n745), .Z(n746) );
  NAND2_X1 U803 ( .A1(n747), .A2(n746), .ZN(n758) );
  XNOR2_X1 U804 ( .A(n749), .B(n748), .ZN(n753) );
  XNOR2_X1 U805 ( .A(G101), .B(KEYINPUT126), .ZN(n750) );
  XNOR2_X1 U806 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U807 ( .A(n753), .B(n752), .ZN(n756) );
  NOR2_X1 U808 ( .A1(n767), .A2(n754), .ZN(n755) );
  NOR2_X1 U809 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n758), .B(n757), .ZN(G69) );
  XNOR2_X1 U811 ( .A(n760), .B(n759), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n761), .B(KEYINPUT127), .ZN(n762) );
  XNOR2_X1 U813 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U814 ( .A(n765), .B(n764), .ZN(n769) );
  XOR2_X1 U815 ( .A(n769), .B(n766), .Z(n768) );
  NAND2_X1 U816 ( .A1(n768), .A2(n767), .ZN(n773) );
  XNOR2_X1 U817 ( .A(G227), .B(n769), .ZN(n770) );
  NAND2_X1 U818 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U819 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U820 ( .A1(n773), .A2(n772), .ZN(G72) );
  XOR2_X1 U821 ( .A(n774), .B(G122), .Z(G24) );
  XNOR2_X1 U822 ( .A(n775), .B(G119), .ZN(G21) );
endmodule

