//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT28), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(G190gat), .ZN(new_n203));
  AND2_X1   g002(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT65), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n203), .B(new_n208), .C1(new_n205), .C2(new_n204), .ZN(new_n209));
  AND2_X1   g008(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(KEYINPUT64), .A2(G183gat), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT27), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n205), .ZN(new_n213));
  AOI21_X1  g012(.A(G190gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n207), .B(new_n209), .C1(new_n214), .C2(KEYINPUT28), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT66), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n219), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  INV_X1    g020(.A(G169gat), .ZN(new_n222));
  INV_X1    g021(.A(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT67), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n229), .A3(new_n226), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(G127gat), .B(G134gat), .ZN(new_n232));
  INV_X1    g031(.A(G113gat), .ZN(new_n233));
  INV_X1    g032(.A(G120gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT1), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n233), .A2(KEYINPUT69), .ZN(new_n238));
  OAI21_X1  g037(.A(G120gat), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(G127gat), .A2(G134gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT68), .B(G127gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(G134gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n235), .B1(new_n233), .B2(new_n234), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT23), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT23), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(G169gat), .B2(G176gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n247), .A2(new_n249), .A3(new_n218), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n226), .A2(KEYINPUT24), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT24), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(G183gat), .A3(G190gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT64), .B(G183gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(G190gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n253), .B2(new_n255), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n251), .B1(new_n261), .B2(new_n250), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n231), .A2(new_n246), .A3(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n231), .A2(KEYINPUT70), .A3(new_n246), .A4(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n231), .A2(new_n263), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n240), .A2(new_n245), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT34), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n271), .A2(KEYINPUT71), .A3(new_n272), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT71), .B1(new_n271), .B2(new_n272), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT32), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT33), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n275), .B2(new_n276), .ZN(new_n279));
  XOR2_X1   g078(.A(G15gat), .B(G43gat), .Z(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n283));
  XOR2_X1   g082(.A(new_n282), .B(new_n283), .Z(new_n284));
  NAND3_X1  g083(.A1(new_n277), .A2(new_n279), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n277), .A2(new_n279), .A3(KEYINPUT74), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n272), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n271), .A2(KEYINPUT71), .A3(new_n272), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(KEYINPUT33), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT32), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n274), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n274), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n298), .B1(new_n287), .B2(new_n288), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT36), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n298), .ZN(new_n301));
  INV_X1    g100(.A(new_n284), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n294), .B2(new_n278), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT74), .B1(new_n303), .B2(new_n277), .ZN(new_n304));
  AND4_X1   g103(.A1(KEYINPUT74), .A2(new_n277), .A3(new_n279), .A4(new_n284), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT36), .ZN(new_n307));
  INV_X1    g106(.A(new_n296), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n308), .B1(new_n287), .B2(new_n288), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n306), .B(new_n307), .C1(new_n309), .C2(new_n274), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n300), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n231), .A2(KEYINPUT76), .A3(new_n263), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT76), .B1(new_n231), .B2(new_n263), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AND2_X1   g115(.A1(G211gat), .A2(G218gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(G211gat), .A2(G218gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT75), .ZN(new_n320));
  OR2_X1    g119(.A1(G197gat), .A2(G204gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G197gat), .A2(G204gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n321), .A2(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n320), .B(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT29), .B1(new_n231), .B2(new_n263), .ZN(new_n327));
  INV_X1    g126(.A(new_n315), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n312), .B1(new_n316), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n268), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n231), .A2(KEYINPUT76), .A3(new_n263), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(new_n328), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n259), .A2(new_n262), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n207), .A2(new_n209), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n205), .B1(new_n257), .B2(KEYINPUT27), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n202), .B1(new_n337), .B2(G190gat), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n336), .A2(new_n338), .B1(KEYINPUT67), .B2(new_n227), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n339), .B2(new_n230), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n315), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n334), .A2(KEYINPUT77), .A3(new_n341), .A4(new_n326), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT37), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n328), .A2(KEYINPUT29), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n332), .A2(new_n333), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n326), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n328), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n330), .A2(new_n342), .A3(new_n343), .A4(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(KEYINPUT78), .ZN(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n330), .A2(new_n348), .A3(new_n342), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(KEYINPUT37), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n355), .B2(KEYINPUT93), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT93), .ZN(new_n357));
  AOI211_X1 g156(.A(new_n357), .B(new_n353), .C1(new_n354), .C2(KEYINPUT37), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT38), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G155gat), .ZN(new_n360));
  INV_X1    g159(.A(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(KEYINPUT80), .B(KEYINPUT2), .Z(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  INV_X1    g166(.A(G141gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G148gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n364), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n373));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n368), .B2(G148gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n366), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n369), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n363), .B1(new_n362), .B2(KEYINPUT2), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n377), .B2(new_n378), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n372), .B(new_n373), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n378), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT82), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n371), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n382), .B(new_n269), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n372), .B1(new_n380), .B2(new_n381), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(new_n269), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n246), .A3(KEYINPUT4), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n388), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n386), .A2(new_n246), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n391), .A2(new_n269), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n389), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n394), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n392), .A2(new_n393), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(KEYINPUT5), .A3(new_n389), .A4(new_n388), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT91), .ZN(new_n403));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(G57gat), .B(G85gat), .ZN(new_n406));
  XOR2_X1   g205(.A(new_n405), .B(new_n406), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n399), .A2(new_n401), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n403), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT6), .B1(new_n402), .B2(new_n407), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT6), .A4(new_n408), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT92), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n342), .A2(new_n348), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n417), .A2(KEYINPUT79), .A3(new_n330), .A4(new_n353), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n345), .A2(new_n326), .A3(new_n347), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n341), .A2(new_n346), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n419), .B(KEYINPUT37), .C1(new_n316), .C2(new_n420), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n353), .A2(KEYINPUT38), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n349), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n330), .A2(new_n342), .A3(new_n348), .A4(new_n353), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n418), .A2(new_n423), .A3(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n416), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n325), .A2(new_n319), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT29), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n325), .B2(new_n319), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n373), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n391), .A2(new_n432), .A3(KEYINPUT85), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT85), .B1(new_n391), .B2(new_n432), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n326), .B1(new_n382), .B2(new_n430), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n436), .A2(new_n438), .B1(G228gat), .B2(G233gat), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT3), .B1(new_n326), .B2(new_n430), .ZN(new_n440));
  OAI211_X1 g239(.A(G228gat), .B(G233gat), .C1(new_n440), .C2(new_n386), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n382), .A2(KEYINPUT86), .A3(new_n430), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n382), .A2(new_n430), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n326), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(G22gat), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(G228gat), .A2(G233gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n391), .A2(new_n432), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n433), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n452), .B2(new_n437), .ZN(new_n453));
  INV_X1    g252(.A(G22gat), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n445), .A2(new_n442), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(new_n441), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT87), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n447), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT88), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n447), .A2(new_n456), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT87), .ZN(new_n461));
  XOR2_X1   g260(.A(G78gat), .B(G106gat), .Z(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT84), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(KEYINPUT31), .ZN(new_n464));
  INV_X1    g263(.A(G50gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT88), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n447), .A2(new_n456), .A3(new_n457), .A4(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n459), .A2(new_n461), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n459), .A2(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n461), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n359), .A2(new_n428), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT30), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n418), .A2(new_n475), .A3(new_n426), .ZN(new_n476));
  OR2_X1    g275(.A1(new_n424), .A2(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(new_n353), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n354), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n483));
  INV_X1    g282(.A(new_n389), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n396), .A2(new_n397), .A3(new_n389), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n485), .A2(KEYINPUT39), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n407), .B1(new_n485), .B2(KEYINPUT39), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT40), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n491), .A2(new_n411), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n418), .A2(new_n475), .A3(new_n426), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(KEYINPUT89), .A3(new_n479), .A4(new_n477), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n481), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n472), .A2(new_n469), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n412), .B1(new_n407), .B2(new_n402), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n414), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n493), .A2(new_n499), .A3(new_n479), .A4(new_n477), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n473), .A2(new_n495), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n306), .B(new_n496), .C1(new_n309), .C2(new_n274), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT35), .B1(new_n502), .B2(new_n500), .ZN(new_n503));
  INV_X1    g302(.A(new_n297), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n481), .A2(new_n494), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n289), .A2(new_n301), .B1(new_n472), .B2(new_n469), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT35), .B1(new_n413), .B2(new_n415), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n311), .A2(new_n501), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  OR2_X1    g309(.A1(new_n510), .A2(G1gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT98), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n513), .B2(G1gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n515), .A3(G8gat), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n510), .A2(G1gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT98), .ZN(new_n518));
  OAI21_X1  g317(.A(G8gat), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n511), .A3(new_n514), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT95), .B(G29gat), .Z(new_n522));
  INV_X1    g321(.A(G36gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT97), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(KEYINPUT96), .A3(KEYINPUT15), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT15), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT96), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n525), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT94), .A3(new_n527), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  INV_X1    g338(.A(new_n527), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(new_n525), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n538), .B(new_n541), .C1(new_n523), .C2(new_n522), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n530), .A2(new_n532), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n536), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n521), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g346(.A1(new_n528), .A2(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT17), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n545), .A2(new_n521), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT18), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n515), .B(new_n519), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(new_n548), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(new_n547), .B2(new_n549), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT18), .A3(new_n551), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n545), .B2(new_n521), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(KEYINPUT99), .A3(new_n548), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n552), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n551), .B(KEYINPUT13), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n555), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G113gat), .B(G141gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(KEYINPUT11), .B(G169gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n555), .A2(new_n559), .A3(new_n571), .A4(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OR2_X1    g375(.A1(G57gat), .A2(G64gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(G57gat), .A2(G64gat), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT9), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n579), .A2(new_n580), .A3(new_n584), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(new_n577), .A3(new_n578), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT100), .B1(new_n582), .B2(new_n583), .ZN(new_n589));
  OR2_X1    g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n580), .A3(new_n581), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(KEYINPUT101), .B(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AND2_X1   g395(.A1(G231gat), .A2(G233gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G127gat), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n521), .B1(KEYINPUT21), .B2(new_n593), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G155gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G134gat), .B(G162gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT102), .B(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(G92gat), .ZN(new_n611));
  OAI21_X1  g410(.A(KEYINPUT7), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n613), .A2(G85gat), .A3(G92gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT8), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n610), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G99gat), .B(G106gat), .Z(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n608), .A2(new_n609), .B1(KEYINPUT8), .B2(new_n616), .ZN(new_n621));
  INV_X1    g420(.A(new_n619), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n621), .A2(new_n622), .A3(new_n615), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625));
  INV_X1    g424(.A(G232gat), .ZN(new_n626));
  INV_X1    g425(.A(G233gat), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI22_X1  g428(.A1(new_n548), .A2(new_n624), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n620), .A2(new_n623), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n545), .B2(new_n546), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n630), .B1(new_n632), .B2(new_n549), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n607), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n635), .ZN(new_n637));
  INV_X1    g436(.A(new_n607), .ZN(new_n638));
  INV_X1    g437(.A(new_n549), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n624), .B1(new_n548), .B2(KEYINPUT17), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n637), .B(new_n638), .C1(new_n641), .C2(new_n630), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n629), .A2(new_n625), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n634), .A2(KEYINPUT103), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n636), .A2(new_n642), .A3(new_n646), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n606), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n624), .A2(new_n594), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n620), .A2(new_n593), .A3(new_n623), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n654), .A2(KEYINPUT104), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT104), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n624), .A2(new_n657), .A3(new_n594), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT10), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT10), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n655), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n653), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n653), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n656), .A2(new_n663), .A3(new_n658), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n662), .A2(new_n664), .A3(new_n668), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n652), .A2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n509), .A2(new_n576), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n499), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT105), .B(G1gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  INV_X1    g478(.A(new_n505), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G8gat), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT16), .B(G8gat), .Z(new_n684));
  NAND3_X1  g483(.A1(new_n675), .A2(new_n680), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n683), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(KEYINPUT106), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(KEYINPUT106), .ZN(new_n688));
  OAI221_X1 g487(.A(new_n682), .B1(new_n683), .B2(new_n685), .C1(new_n687), .C2(new_n688), .ZN(G1325gat));
  INV_X1    g488(.A(G15gat), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n297), .A2(new_n299), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n311), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n675), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n694), .B2(new_n690), .ZN(G1326gat));
  NAND2_X1  g494(.A1(new_n675), .A2(new_n497), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  NAND2_X1  g497(.A1(new_n503), .A2(new_n508), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n473), .A2(new_n495), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n497), .A2(new_n500), .ZN(new_n701));
  NAND4_X1  g500(.A1(new_n700), .A2(new_n300), .A3(new_n310), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n606), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(new_n576), .A3(new_n672), .ZN(new_n705));
  AND3_X1   g504(.A1(new_n703), .A2(new_n651), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n706), .A2(new_n676), .A3(new_n522), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n509), .B2(new_n650), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n651), .ZN(new_n711));
  AND2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n712), .A2(new_n705), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n713), .A2(new_n676), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n708), .B1(new_n714), .B2(new_n522), .ZN(G1328gat));
  NAND3_X1  g514(.A1(new_n706), .A2(new_n523), .A3(new_n680), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n716), .B(KEYINPUT46), .Z(new_n717));
  AND2_X1   g516(.A1(new_n713), .A2(new_n680), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n523), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n710), .A2(new_n693), .A3(new_n711), .A4(new_n705), .ZN(new_n720));
  INV_X1    g519(.A(new_n691), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n721), .A2(G43gat), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n720), .A2(G43gat), .B1(new_n706), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n497), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n465), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n496), .A2(new_n465), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n710), .A2(new_n711), .A3(new_n705), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(KEYINPUT108), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT48), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n726), .A2(new_n734), .A3(new_n728), .A4(new_n729), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n731), .A2(new_n733), .A3(new_n735), .ZN(G1331gat));
  NOR4_X1   g535(.A1(new_n606), .A2(new_n575), .A3(new_n651), .A4(new_n673), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n703), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n499), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT109), .B(G57gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1332gat));
  OR2_X1    g540(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n505), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  OR2_X1    g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n311), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n742), .A2(new_n743), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n703), .A2(new_n691), .A3(new_n737), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n750), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n742), .A2(new_n753), .A3(new_n743), .A4(new_n751), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n756), .B2(new_n758), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n497), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n606), .A2(new_n576), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT113), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n765), .A2(new_n672), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n712), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n499), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n703), .A2(new_n651), .A3(new_n765), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n703), .A2(KEYINPUT51), .A3(new_n651), .A4(new_n765), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n676), .A2(new_n609), .A3(new_n672), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  NAND4_X1  g575(.A1(new_n710), .A2(new_n680), .A3(new_n711), .A4(new_n766), .ZN(new_n777));
  INV_X1    g576(.A(new_n608), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n680), .A2(new_n611), .A3(new_n672), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT52), .ZN(G1337gat));
  OAI21_X1  g581(.A(G99gat), .B1(new_n767), .B2(new_n311), .ZN(new_n783));
  OR3_X1    g582(.A1(new_n721), .A2(G99gat), .A3(new_n673), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n774), .B2(new_n784), .ZN(G1338gat));
  NAND4_X1  g584(.A1(new_n710), .A2(new_n497), .A3(new_n711), .A4(new_n766), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n496), .A2(G106gat), .A3(new_n673), .ZN(new_n787));
  AOI22_X1  g586(.A1(G106gat), .A2(new_n786), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT114), .B1(new_n786), .B2(G106gat), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n788), .A2(KEYINPUT53), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(G106gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n773), .A2(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(KEYINPUT53), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n790), .A2(new_n795), .ZN(G1339gat));
  OAI21_X1  g595(.A(new_n669), .B1(new_n662), .B2(KEYINPUT54), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n655), .A2(KEYINPUT104), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n593), .B1(new_n623), .B2(new_n620), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n658), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n660), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n661), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n800), .B1(new_n807), .B2(new_n653), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n805), .A2(new_n663), .A3(new_n806), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n799), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n809), .A2(new_n662), .A3(new_n799), .A4(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n798), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(new_n564), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n561), .A2(new_n562), .A3(new_n552), .A4(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n558), .B2(new_n551), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(new_n570), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n818), .A2(KEYINPUT116), .A3(new_n570), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n574), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n650), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n662), .A3(KEYINPUT54), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT115), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n797), .B1(new_n826), .B2(new_n811), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT55), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n815), .A2(new_n671), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n671), .B1(new_n827), .B2(KEYINPUT55), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n833), .A2(KEYINPUT117), .A3(new_n828), .A4(new_n824), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n815), .A2(new_n575), .A3(new_n671), .A4(new_n828), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n823), .A2(new_n673), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n651), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n606), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n652), .A2(new_n576), .A3(new_n673), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n499), .B1(new_n481), .B2(new_n494), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n502), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n575), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n237), .A2(new_n238), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n233), .B2(new_n847), .ZN(G1340gat));
  AOI22_X1  g649(.A1(new_n846), .A2(new_n672), .B1(KEYINPUT118), .B2(new_n234), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n234), .A2(KEYINPUT118), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(G1341gat));
  NAND2_X1  g652(.A1(new_n846), .A2(new_n704), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(new_n242), .ZN(G1342gat));
  AOI21_X1  g654(.A(new_n650), .B1(KEYINPUT56), .B2(G134gat), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n844), .A2(new_n845), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT119), .ZN(new_n858));
  NOR2_X1   g657(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n858), .B(new_n859), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n693), .A2(new_n496), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n368), .A2(new_n844), .A3(new_n575), .A4(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(KEYINPUT58), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n300), .A2(new_n310), .A3(new_n843), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n300), .A2(KEYINPUT120), .A3(new_n310), .A4(new_n843), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n842), .B2(new_n497), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  AOI211_X1 g670(.A(new_n871), .B(new_n496), .C1(new_n840), .C2(new_n841), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n576), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT121), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n841), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n814), .B(new_n797), .C1(new_n826), .C2(new_n811), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n832), .A2(new_n576), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n650), .B1(new_n880), .B2(new_n837), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n831), .A3(new_n834), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n882), .B2(new_n606), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n871), .B1(new_n883), .B2(new_n496), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n842), .A2(KEYINPUT57), .A3(new_n497), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(KEYINPUT121), .A3(new_n869), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n877), .A2(new_n575), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n862), .B1(new_n888), .B2(G141gat), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n875), .B1(new_n889), .B2(new_n890), .ZN(G1344gat));
  AND2_X1   g690(.A1(new_n844), .A2(new_n861), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n892), .A2(new_n366), .A3(new_n672), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G148gat), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT121), .B1(new_n886), .B2(new_n869), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n876), .B(new_n868), .C1(new_n884), .C2(new_n885), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n895), .B1(new_n898), .B2(new_n672), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n885), .A2(KEYINPUT122), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT122), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n842), .A2(new_n901), .A3(KEYINPUT57), .A4(new_n497), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n704), .B1(new_n881), .B2(new_n829), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n497), .B1(new_n905), .B2(new_n878), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n906), .B2(new_n871), .ZN(new_n907));
  INV_X1    g706(.A(new_n829), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n606), .B1(new_n839), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n496), .B1(new_n909), .B2(new_n841), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n672), .B(new_n869), .C1(new_n903), .C2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n894), .B1(new_n913), .B2(G148gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n893), .B1(new_n899), .B2(new_n914), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n892), .A2(new_n360), .A3(new_n704), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n896), .A2(new_n897), .A3(new_n606), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n360), .ZN(G1346gat));
  AOI21_X1  g717(.A(G162gat), .B1(new_n892), .B2(new_n651), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n650), .A2(new_n361), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n898), .B2(new_n920), .ZN(G1347gat));
  NAND2_X1  g720(.A1(new_n680), .A2(new_n499), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n502), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n842), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g723(.A(new_n924), .B(KEYINPUT124), .Z(new_n925));
  AOI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n575), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n924), .B(KEYINPUT125), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(new_n222), .A3(new_n576), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n223), .A3(new_n672), .ZN(new_n930));
  OAI21_X1  g729(.A(G176gat), .B1(new_n927), .B2(new_n673), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1349gat));
  OAI21_X1  g731(.A(new_n704), .B1(new_n205), .B2(new_n204), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n934), .B(KEYINPUT126), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n257), .B1(new_n927), .B2(new_n606), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  INV_X1    g740(.A(G190gat), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n942), .A3(new_n651), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  INV_X1    g743(.A(new_n927), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n651), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n946), .B2(G190gat), .ZN(new_n947));
  AOI211_X1 g746(.A(KEYINPUT61), .B(new_n942), .C1(new_n945), .C2(new_n651), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n943), .B1(new_n947), .B2(new_n948), .ZN(G1351gat));
  NOR2_X1   g748(.A1(new_n883), .A2(new_n496), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n693), .A2(new_n922), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n575), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n903), .A2(new_n912), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(new_n951), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n575), .A2(G197gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1352gat));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n672), .A3(new_n951), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(G204gat), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n952), .A2(G204gat), .A3(new_n673), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT62), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1353gat));
  OAI211_X1 g762(.A(new_n704), .B(new_n951), .C1(new_n903), .C2(new_n912), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(G211gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT63), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT63), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n967), .A3(G211gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n952), .A2(G211gat), .A3(new_n606), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n968), .A3(new_n971), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n651), .A3(new_n951), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(G218gat), .ZN(new_n974));
  OR3_X1    g773(.A1(new_n952), .A2(G218gat), .A3(new_n650), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1355gat));
endmodule


