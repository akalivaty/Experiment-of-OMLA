//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT91), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT91), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT14), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n205), .B(new_n209), .C1(G29gat), .C2(G36gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT15), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(G50gat), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(G43gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT92), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n212), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n218), .A2(new_n208), .A3(new_n207), .A4(new_n210), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n214), .A3(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n207), .A2(new_n210), .ZN(new_n221));
  INV_X1    g020(.A(new_n214), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n221), .A2(new_n222), .A3(new_n218), .A4(new_n208), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(G1gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT16), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G1gat), .B2(new_n227), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n220), .A2(KEYINPUT17), .A3(new_n223), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n226), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n231), .B(G8gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n224), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n224), .B(new_n236), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n238), .B(KEYINPUT13), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n237), .A4(new_n238), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G141gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G169gat), .B(G197gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(KEYINPUT90), .B(KEYINPUT12), .Z(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n241), .A2(new_n254), .A3(new_n245), .A4(new_n246), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT93), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n257), .A2(new_n258), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  XNOR2_X1  g062(.A(G127gat), .B(G134gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT66), .ZN(new_n265));
  INV_X1    g064(.A(G113gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n265), .B1(new_n266), .B2(G120gat), .ZN(new_n267));
  INV_X1    g066(.A(G120gat), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(KEYINPUT66), .A3(G113gat), .ZN(new_n269));
  AOI22_X1  g068(.A1(new_n267), .A2(new_n269), .B1(new_n266), .B2(G120gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n263), .B(new_n264), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  AND2_X1   g071(.A1(new_n270), .A2(new_n271), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n264), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G127gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(G134gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(G113gat), .B(G120gat), .ZN(new_n279));
  OAI221_X1 g078(.A(new_n276), .B1(new_n275), .B2(new_n278), .C1(KEYINPUT1), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT76), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n280), .B(KEYINPUT76), .C1(new_n273), .C2(new_n272), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n286), .B1(new_n289), .B2(KEYINPUT2), .ZN(new_n290));
  XOR2_X1   g089(.A(G141gat), .B(G148gat), .Z(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT75), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n291), .ZN(new_n295));
  XOR2_X1   g094(.A(KEYINPUT74), .B(KEYINPUT2), .Z(new_n296));
  OAI211_X1 g095(.A(new_n286), .B(new_n289), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n285), .A2(KEYINPUT78), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT76), .B1(new_n274), .B2(new_n280), .ZN(new_n300));
  INV_X1    g099(.A(new_n284), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n281), .A2(new_n298), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n299), .A2(new_n304), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT84), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n298), .B(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n285), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n305), .A2(KEYINPUT4), .ZN(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n307), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT39), .B1(new_n310), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  XOR2_X1   g123(.A(G1gat), .B(G29gat), .Z(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n325), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G57gat), .B(G85gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n310), .A2(new_n322), .A3(KEYINPUT39), .A4(new_n319), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT40), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n318), .B1(new_n305), .B2(KEYINPUT4), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n313), .B(new_n335), .C1(new_n305), .C2(new_n315), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n299), .A2(new_n306), .A3(new_n304), .ZN(new_n337));
  OAI211_X1 g136(.A(KEYINPUT5), .B(new_n336), .C1(new_n337), .C2(new_n307), .ZN(new_n338));
  OR3_X1    g137(.A1(new_n317), .A2(KEYINPUT5), .A3(new_n318), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT86), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT86), .B1(new_n338), .B2(new_n339), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n329), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT30), .ZN(new_n344));
  NAND2_X1  g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT72), .Z(new_n346));
  INV_X1    g145(.A(KEYINPUT25), .ZN(new_n347));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT24), .ZN(new_n349));
  OR3_X1    g148(.A1(new_n348), .A2(new_n349), .A3(KEYINPUT64), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n348), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT64), .B1(new_n348), .B2(new_n349), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT23), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n347), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n352), .B1(new_n349), .B2(new_n348), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(new_n362), .A3(new_n347), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT27), .B(G183gat), .ZN(new_n367));
  INV_X1    g166(.A(G190gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT28), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n358), .A2(KEYINPUT26), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT28), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n367), .A2(new_n372), .A3(new_n368), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n370), .A2(new_n348), .A3(new_n371), .A4(new_n373), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n357), .A2(KEYINPUT26), .A3(new_n358), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n364), .B(new_n366), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT29), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n346), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT73), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G197gat), .B(G204gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT70), .B(G218gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n381), .B1(new_n382), .B2(KEYINPUT22), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G211gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(KEYINPUT22), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(G218gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AND2_X1   g188(.A1(new_n376), .A2(new_n346), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(new_n378), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n380), .B(new_n389), .C1(new_n391), .C2(KEYINPUT73), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(KEYINPUT71), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT71), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n396), .B1(new_n378), .B2(new_n390), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G8gat), .B(G36gat), .Z(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G64gat), .ZN(new_n400));
  INV_X1    g199(.A(G92gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n344), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n402), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n392), .A2(new_n397), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n344), .A3(new_n404), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT83), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n408), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n324), .A2(KEYINPUT40), .A3(new_n330), .A4(new_n331), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n334), .A2(new_n343), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n298), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n389), .A2(new_n377), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n419), .B2(new_n311), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n418), .B2(new_n311), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(new_n389), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n417), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT82), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(new_n417), .C1(new_n420), .C2(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(G22gat), .B(G50gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n421), .B1(new_n393), .B2(new_n395), .ZN(new_n432));
  OR3_X1    g231(.A1(new_n420), .A2(new_n432), .A3(new_n417), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n427), .B2(new_n433), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n416), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(new_n433), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n430), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n427), .A2(new_n431), .A3(new_n433), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n415), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n436), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT6), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n338), .A2(new_n339), .A3(new_n330), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n343), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT37), .ZN(new_n450));
  NOR2_X1   g249(.A1(new_n407), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n402), .B1(new_n398), .B2(KEYINPUT37), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT38), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n380), .B1(new_n391), .B2(KEYINPUT73), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n388), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n391), .A2(new_n393), .A3(new_n395), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n450), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OR3_X1    g256(.A1(new_n452), .A2(new_n457), .A3(KEYINPUT38), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(new_n405), .A3(new_n453), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n414), .A2(new_n441), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT80), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n447), .B2(new_n442), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n338), .A2(new_n339), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n329), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n464), .A2(KEYINPUT80), .A3(new_n446), .A4(new_n445), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n443), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n408), .ZN(new_n467));
  INV_X1    g266(.A(new_n406), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n436), .A2(new_n440), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  XOR2_X1   g270(.A(G71gat), .B(G99gat), .Z(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT68), .ZN(new_n473));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n376), .B(new_n281), .ZN(new_n477));
  NAND2_X1  g276(.A1(G227gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT33), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT34), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n477), .A2(new_n479), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT69), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n480), .A2(KEYINPUT32), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n486), .A3(new_n484), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n483), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n490), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT32), .B(new_n480), .C1(new_n494), .C2(new_n487), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(new_n482), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT36), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n460), .A2(new_n471), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n449), .B2(new_n412), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n408), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n409), .ZN(new_n504));
  INV_X1    g303(.A(new_n342), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n340), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n447), .B1(new_n506), .B2(new_n329), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n504), .B(KEYINPUT87), .C1(new_n507), .C2(new_n444), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  INV_X1    g308(.A(new_n498), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n510), .A2(new_n470), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n502), .A2(new_n508), .A3(new_n509), .A4(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n441), .A2(new_n498), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT35), .B1(new_n469), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT88), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n515), .A3(KEYINPUT88), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n262), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521));
  INV_X1    g320(.A(G85gat), .ZN(new_n522));
  AOI22_X1  g321(.A1(KEYINPUT8), .A2(new_n521), .B1(new_n522), .B2(new_n401), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(new_n522), .B2(new_n401), .ZN(new_n525));
  NAND3_X1  g324(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n523), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G99gat), .B(G106gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n226), .A2(new_n234), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n224), .A2(new_n529), .B1(KEYINPUT41), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G134gat), .B(G162gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n532), .A2(KEYINPUT41), .ZN(new_n537));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n536), .B(new_n539), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(G71gat), .A2(G78gat), .ZN(new_n542));
  XOR2_X1   g341(.A(G57gat), .B(G64gat), .Z(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT9), .ZN(new_n544));
  NOR2_X1   g343(.A1(G71gat), .A2(G78gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT94), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT95), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n545), .A2(KEYINPUT9), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n543), .B1(new_n549), .B2(new_n542), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(KEYINPUT10), .A3(new_n529), .ZN(new_n553));
  INV_X1    g352(.A(new_n528), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT97), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n548), .A2(new_n550), .A3(new_n529), .A4(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT95), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n558), .B1(new_n544), .B2(new_n546), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n550), .B(new_n555), .C1(new_n557), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n530), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT10), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n556), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G230gat), .A2(G233gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n565), .B1(new_n556), .B2(new_n561), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT98), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G120gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n571), .B(G148gat), .Z(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n568), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n565), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n553), .B2(new_n563), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n572), .B1(new_n576), .B2(new_n567), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n552), .A2(KEYINPUT21), .ZN(new_n579));
  XNOR2_X1  g378(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(G211gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n233), .B1(new_n551), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G183gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT96), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n589), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n592), .B1(new_n588), .B2(new_n589), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n583), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n582), .A3(new_n593), .ZN(new_n598));
  AOI211_X1 g397(.A(new_n541), .B(new_n578), .C1(new_n596), .C2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT99), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n520), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n466), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n228), .ZN(G1324gat));
  NOR2_X1   g402(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n601), .A2(new_n504), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT101), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(KEYINPUT42), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT42), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(KEYINPUT101), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(G8gat), .B1(new_n601), .B2(new_n504), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT100), .Z(new_n612));
  NAND4_X1  g411(.A1(new_n605), .A2(new_n607), .A3(KEYINPUT42), .A4(new_n606), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(new_n612), .A3(new_n613), .ZN(G1325gat));
  INV_X1    g413(.A(G15gat), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n601), .A2(new_n615), .A3(new_n499), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n520), .A2(new_n498), .A3(new_n600), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(G1326gat));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n441), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT43), .B(G22gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(G1327gat));
  NAND2_X1  g420(.A1(new_n596), .A2(new_n598), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n578), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n541), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n500), .A2(new_n515), .A3(KEYINPUT88), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT88), .B1(new_n500), .B2(new_n515), .ZN(new_n627));
  OAI221_X1 g426(.A(new_n261), .B1(KEYINPUT102), .B2(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(KEYINPUT102), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n466), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(new_n202), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT45), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n540), .B1(new_n500), .B2(new_n515), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n635), .A2(KEYINPUT44), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n540), .B1(new_n518), .B2(new_n519), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(KEYINPUT44), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n639), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n241), .A2(new_n246), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n642), .A2(KEYINPUT93), .A3(new_n254), .A4(new_n245), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n257), .A2(new_n258), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n639), .B1(new_n645), .B2(new_n256), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n622), .A2(new_n647), .A3(new_n578), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n638), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(G29gat), .B1(new_n649), .B2(new_n466), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n650), .ZN(G1328gat));
  NAND3_X1  g450(.A1(new_n631), .A2(new_n203), .A3(new_n412), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n652), .A2(KEYINPUT46), .ZN(new_n653));
  OAI21_X1  g452(.A(G36gat), .B1(new_n649), .B2(new_n504), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(KEYINPUT46), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(G1329gat));
  OAI21_X1  g455(.A(G43gat), .B1(new_n649), .B2(new_n499), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT104), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n510), .A2(G43gat), .ZN(new_n659));
  AND3_X1   g458(.A1(new_n631), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n658), .B1(new_n631), .B2(new_n659), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT47), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1330gat));
  NAND2_X1  g463(.A1(new_n470), .A2(new_n215), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT105), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n631), .A2(new_n666), .B1(KEYINPUT106), .B2(KEYINPUT48), .ZN(new_n667));
  OAI211_X1 g466(.A(KEYINPUT44), .B(new_n541), .C1(new_n626), .C2(new_n627), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n635), .A2(KEYINPUT44), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n668), .A2(new_n669), .A3(new_n470), .A4(new_n648), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT48), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n671), .A3(G50gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n631), .A2(KEYINPUT106), .A3(new_n666), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT107), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n670), .B(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(G50gat), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT108), .B(new_n673), .C1(new_n678), .C2(new_n671), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n638), .A2(new_n676), .A3(new_n470), .A4(new_n648), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n670), .A2(KEYINPUT107), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(G50gat), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n671), .B1(new_n683), .B2(new_n674), .ZN(new_n684));
  INV_X1    g483(.A(new_n673), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n679), .A2(new_n686), .ZN(G1331gat));
  AOI211_X1 g486(.A(new_n623), .B(new_n541), .C1(new_n500), .C2(new_n515), .ZN(new_n688));
  INV_X1    g487(.A(new_n647), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(new_n624), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n632), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g493(.A1(new_n691), .A2(new_n504), .ZN(new_n695));
  NOR2_X1   g494(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n696));
  AND2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n695), .B2(new_n696), .ZN(G1333gat));
  OR3_X1    g498(.A1(new_n691), .A2(G71gat), .A3(new_n510), .ZN(new_n700));
  OAI21_X1  g499(.A(G71gat), .B1(new_n691), .B2(new_n499), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT109), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g503(.A1(new_n691), .A2(new_n441), .ZN(new_n705));
  XOR2_X1   g504(.A(KEYINPUT110), .B(G78gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1335gat));
  NOR2_X1   g506(.A1(new_n689), .A2(new_n622), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n638), .A2(new_n578), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n522), .A3(new_n466), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n635), .A2(new_n708), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT51), .Z(new_n712));
  NAND3_X1  g511(.A1(new_n712), .A2(new_n632), .A3(new_n578), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n710), .B1(new_n522), .B2(new_n713), .ZN(G1336gat));
  OAI21_X1  g513(.A(G92gat), .B1(new_n709), .B2(new_n504), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n712), .A2(new_n401), .A3(new_n412), .A4(new_n578), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT52), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT111), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n717), .B(new_n720), .ZN(G1337gat));
  OAI21_X1  g520(.A(G99gat), .B1(new_n709), .B2(new_n499), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n510), .A2(G99gat), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n712), .A2(new_n578), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1338gat));
  OAI21_X1  g524(.A(G106gat), .B1(new_n709), .B2(new_n441), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n441), .A2(G106gat), .A3(new_n624), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT112), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n553), .A2(new_n563), .A3(new_n575), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n566), .A2(KEYINPUT54), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT54), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n573), .B1(new_n576), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT55), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n734), .A2(KEYINPUT55), .A3(new_n736), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n574), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n261), .A2(KEYINPUT103), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(new_n640), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n235), .A2(new_n237), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n744), .A2(new_n238), .B1(new_n242), .B2(new_n244), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n252), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT114), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(new_n645), .A3(new_n578), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n732), .B1(new_n743), .B2(new_n749), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n739), .A2(new_n574), .A3(new_n740), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n751), .B1(new_n641), .B2(new_n646), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(KEYINPUT115), .A3(new_n748), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n750), .A2(new_n753), .A3(new_n540), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n751), .A2(new_n645), .A3(new_n541), .A4(new_n747), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT116), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(KEYINPUT116), .A3(new_n755), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n623), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n599), .A2(new_n647), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT113), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n513), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n632), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(new_n504), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n266), .A3(new_n689), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n765), .A2(new_n412), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G113gat), .B1(new_n771), .B2(new_n262), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n772), .ZN(G1340gat));
  NAND3_X1  g572(.A1(new_n768), .A2(new_n268), .A3(new_n578), .ZN(new_n774));
  OAI21_X1  g573(.A(G120gat), .B1(new_n771), .B2(new_n624), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1341gat));
  NOR3_X1   g575(.A1(new_n771), .A2(new_n277), .A3(new_n623), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n768), .A2(new_n622), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n277), .ZN(G1342gat));
  NOR2_X1   g578(.A1(new_n540), .A2(G134gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n767), .A2(new_n504), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT56), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT118), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n781), .A2(KEYINPUT56), .ZN(new_n784));
  OAI21_X1  g583(.A(G134gat), .B1(new_n771), .B2(new_n540), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n781), .A2(new_n786), .A3(KEYINPUT56), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n783), .A2(new_n784), .A3(new_n785), .A4(new_n787), .ZN(G1343gat));
  NAND3_X1  g587(.A1(new_n499), .A2(new_n632), .A3(new_n504), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n749), .B1(new_n261), .B2(new_n751), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n755), .B1(new_n792), .B2(new_n541), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n793), .A2(new_n623), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT120), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n791), .B(new_n441), .C1(new_n795), .C2(new_n763), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n441), .B1(new_n760), .B2(new_n763), .ZN(new_n797));
  XNOR2_X1  g596(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n790), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(G141gat), .B1(new_n800), .B2(new_n262), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n797), .A2(new_n790), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n802), .A2(G141gat), .A3(new_n262), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(KEYINPUT58), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n689), .B(new_n790), .C1(new_n796), .C2(new_n799), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n803), .B1(new_n806), .B2(G141gat), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT121), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n807), .A2(new_n811), .A3(new_n808), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n810), .B2(new_n812), .ZN(G1344gat));
  INV_X1    g612(.A(KEYINPUT59), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n814), .B(G148gat), .C1(new_n800), .C2(new_n624), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n754), .A2(KEYINPUT116), .A3(new_n755), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT116), .B1(new_n754), .B2(new_n755), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n818), .A3(new_n622), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n470), .B(new_n798), .C1(new_n819), .C2(new_n762), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n794), .B1(new_n600), .B2(new_n262), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n791), .B1(new_n823), .B2(new_n441), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n797), .A2(KEYINPUT122), .A3(new_n798), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n578), .A3(new_n790), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G148gat), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n816), .B1(new_n828), .B2(KEYINPUT59), .ZN(new_n829));
  AOI211_X1 g628(.A(KEYINPUT123), .B(new_n814), .C1(new_n827), .C2(G148gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n815), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n802), .A2(G148gat), .A3(new_n624), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1345gat));
  NOR3_X1   g632(.A1(new_n800), .A2(new_n287), .A3(new_n623), .ZN(new_n834));
  INV_X1    g633(.A(new_n802), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n622), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT124), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n837), .B2(new_n287), .ZN(G1346gat));
  NOR3_X1   g637(.A1(new_n800), .A2(new_n288), .A3(new_n540), .ZN(new_n839));
  AOI21_X1  g638(.A(G162gat), .B1(new_n835), .B2(new_n541), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(G1347gat));
  NOR2_X1   g640(.A1(new_n632), .A2(new_n504), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n764), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n844), .A2(new_n355), .A3(new_n689), .ZN(new_n845));
  OAI21_X1  g644(.A(G169gat), .B1(new_n843), .B2(new_n262), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1348gat));
  NOR2_X1   g646(.A1(new_n843), .A2(new_n624), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n356), .ZN(G1349gat));
  NAND3_X1  g648(.A1(new_n844), .A2(new_n367), .A3(new_n622), .ZN(new_n850));
  OAI21_X1  g649(.A(G183gat), .B1(new_n843), .B2(new_n623), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n850), .B(new_n851), .C1(KEYINPUT125), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(KEYINPUT125), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n853), .B(new_n854), .ZN(G1350gat));
  NOR2_X1   g654(.A1(new_n843), .A2(new_n540), .ZN(new_n856));
  NAND2_X1  g655(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g657(.A(KEYINPUT61), .B(G190gat), .Z(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n856), .B2(new_n859), .ZN(G1351gat));
  AND2_X1   g659(.A1(new_n842), .A2(new_n499), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n797), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT126), .ZN(new_n863));
  INV_X1    g662(.A(G197gat), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n863), .A2(new_n864), .A3(new_n689), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(KEYINPUT127), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(KEYINPUT127), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n826), .A2(new_n261), .A3(new_n861), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n866), .A2(new_n867), .B1(new_n864), .B2(new_n868), .ZN(G1352gat));
  NOR3_X1   g668(.A1(new_n862), .A2(G204gat), .A3(new_n624), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT62), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n826), .A2(new_n578), .A3(new_n861), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G204gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(G1353gat));
  NAND3_X1  g673(.A1(new_n863), .A2(new_n385), .A3(new_n622), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n826), .A2(new_n622), .A3(new_n861), .ZN(new_n876));
  AND3_X1   g675(.A1(new_n876), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT63), .B1(new_n876), .B2(G211gat), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(G1354gat));
  AOI21_X1  g678(.A(G218gat), .B1(new_n863), .B2(new_n541), .ZN(new_n880));
  AND4_X1   g679(.A1(new_n382), .A2(new_n826), .A3(new_n541), .A4(new_n861), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(G1355gat));
endmodule


