

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728;

  BUF_X1 U365 ( .A(n686), .Z(n344) );
  NOR2_X1 U366 ( .A1(n725), .A2(n724), .ZN(n556) );
  NOR2_X1 U367 ( .A1(n674), .A2(n671), .ZN(n550) );
  NOR2_X1 U368 ( .A1(n570), .A2(n573), .ZN(n466) );
  BUF_X1 U369 ( .A(n481), .Z(n563) );
  XNOR2_X1 U370 ( .A(n346), .B(n345), .ZN(n441) );
  INV_X1 U371 ( .A(n415), .ZN(n345) );
  XOR2_X1 U372 ( .A(G101), .B(KEYINPUT4), .Z(n446) );
  AND2_X1 U373 ( .A1(n484), .A2(G234), .ZN(n392) );
  XNOR2_X2 U374 ( .A(n712), .B(G146), .ZN(n473) );
  NOR2_X2 U375 ( .A1(n520), .A2(n551), .ZN(n346) );
  BUF_X1 U376 ( .A(G143), .Z(n639) );
  XNOR2_X2 U377 ( .A(n362), .B(n494), .ZN(n523) );
  NOR2_X1 U378 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U379 ( .A(n364), .B(G122), .ZN(n448) );
  XNOR2_X1 U380 ( .A(G140), .B(G137), .ZN(n468) );
  XNOR2_X1 U381 ( .A(KEYINPUT104), .B(KEYINPUT30), .ZN(n543) );
  BUF_X1 U382 ( .A(n608), .Z(n618) );
  XNOR2_X2 U383 ( .A(n437), .B(n424), .ZN(n712) );
  XNOR2_X1 U384 ( .A(G146), .B(G125), .ZN(n453) );
  XNOR2_X1 U385 ( .A(n567), .B(n376), .ZN(n373) );
  INV_X1 U386 ( .A(KEYINPUT83), .ZN(n376) );
  XNOR2_X1 U387 ( .A(n566), .B(KEYINPUT77), .ZN(n372) );
  NOR2_X1 U388 ( .A1(n726), .A2(n504), .ZN(n506) );
  XNOR2_X1 U389 ( .A(G137), .B(G116), .ZN(n383) );
  XNOR2_X1 U390 ( .A(n349), .B(n382), .ZN(n450) );
  XNOR2_X1 U391 ( .A(KEYINPUT3), .B(KEYINPUT72), .ZN(n382) );
  XNOR2_X1 U392 ( .A(n453), .B(n452), .ZN(n454) );
  AND2_X1 U393 ( .A1(n358), .A2(n350), .ZN(n355) );
  NAND2_X1 U394 ( .A1(n509), .A2(n347), .ZN(n358) );
  OR2_X1 U395 ( .A1(n526), .A2(KEYINPUT101), .ZN(n356) );
  XNOR2_X1 U396 ( .A(n464), .B(n463), .ZN(n481) );
  AND2_X1 U397 ( .A1(n492), .A2(n508), .ZN(n363) );
  XNOR2_X1 U398 ( .A(n447), .B(G107), .ZN(n701) );
  XNOR2_X1 U399 ( .A(n450), .B(n449), .ZN(n702) );
  XNOR2_X1 U400 ( .A(n448), .B(KEYINPUT16), .ZN(n449) );
  XNOR2_X1 U401 ( .A(n701), .B(n360), .ZN(n472) );
  XNOR2_X1 U402 ( .A(n446), .B(KEYINPUT73), .ZN(n360) );
  XNOR2_X1 U403 ( .A(n378), .B(n377), .ZN(n569) );
  INV_X1 U404 ( .A(KEYINPUT39), .ZN(n377) );
  NOR2_X1 U405 ( .A1(n562), .A2(n379), .ZN(n378) );
  XNOR2_X1 U406 ( .A(n491), .B(KEYINPUT0), .ZN(n507) );
  NAND2_X1 U407 ( .A1(n370), .A2(n375), .ZN(n369) );
  INV_X1 U408 ( .A(G116), .ZN(n364) );
  XOR2_X1 U409 ( .A(G140), .B(G104), .Z(n426) );
  XNOR2_X1 U410 ( .A(n473), .B(n365), .ZN(n593) );
  XNOR2_X1 U411 ( .A(n366), .B(n387), .ZN(n365) );
  XNOR2_X1 U412 ( .A(n450), .B(n384), .ZN(n366) );
  INV_X2 U413 ( .A(G953), .ZN(n484) );
  XNOR2_X1 U414 ( .A(n389), .B(G110), .ZN(n391) );
  XNOR2_X1 U415 ( .A(G119), .B(KEYINPUT23), .ZN(n389) );
  XNOR2_X1 U416 ( .A(KEYINPUT24), .B(G128), .ZN(n390) );
  INV_X1 U417 ( .A(G134), .ZN(n381) );
  XNOR2_X1 U418 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U419 ( .A(n359), .B(n352), .ZN(n687) );
  NAND2_X1 U420 ( .A1(n355), .A2(n354), .ZN(n359) );
  OR2_X1 U421 ( .A1(n509), .A2(KEYINPUT101), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n493), .B(KEYINPUT76), .ZN(n494) );
  NAND2_X1 U423 ( .A1(n507), .A2(n363), .ZN(n362) );
  INV_X1 U424 ( .A(KEYINPUT22), .ZN(n493) );
  XNOR2_X1 U425 ( .A(n361), .B(n472), .ZN(n474) );
  XNOR2_X1 U426 ( .A(n471), .B(KEYINPUT78), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n470), .B(n469), .ZN(n471) );
  AND2_X1 U428 ( .A1(n569), .A2(n641), .ZN(n549) );
  NOR2_X2 U429 ( .A1(n558), .A2(n557), .ZN(n640) );
  AND2_X1 U430 ( .A1(n526), .A2(KEYINPUT101), .ZN(n347) );
  AND2_X1 U431 ( .A1(n372), .A2(n568), .ZN(n348) );
  XOR2_X1 U432 ( .A(G113), .B(G119), .Z(n349) );
  XNOR2_X1 U433 ( .A(n556), .B(KEYINPUT46), .ZN(n375) );
  AND2_X1 U434 ( .A1(n357), .A2(n356), .ZN(n350) );
  AND2_X1 U435 ( .A1(n373), .A2(n375), .ZN(n351) );
  XOR2_X1 U436 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n352) );
  XOR2_X1 U437 ( .A(KEYINPUT75), .B(KEYINPUT34), .Z(n353) );
  XNOR2_X2 U438 ( .A(n414), .B(n413), .ZN(n551) );
  XNOR2_X2 U439 ( .A(n542), .B(KEYINPUT6), .ZN(n520) );
  OR2_X2 U440 ( .A1(n610), .A2(G902), .ZN(n402) );
  NAND2_X1 U441 ( .A1(n509), .A2(n526), .ZN(n530) );
  INV_X1 U442 ( .A(n520), .ZN(n357) );
  XNOR2_X2 U443 ( .A(n457), .B(n381), .ZN(n437) );
  NAND2_X1 U444 ( .A1(n368), .A2(n367), .ZN(n577) );
  NAND2_X1 U445 ( .A1(n351), .A2(n348), .ZN(n367) );
  NAND2_X1 U446 ( .A1(n369), .A2(n374), .ZN(n368) );
  INV_X1 U447 ( .A(n371), .ZN(n370) );
  NAND2_X1 U448 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U449 ( .A(n568), .ZN(n374) );
  NAND2_X1 U450 ( .A1(n477), .A2(n509), .ZN(n567) );
  INV_X1 U451 ( .A(n669), .ZN(n379) );
  NAND2_X1 U452 ( .A1(n547), .A2(n548), .ZN(n562) );
  XNOR2_X1 U453 ( .A(n446), .B(n383), .ZN(n384) );
  XOR2_X1 U454 ( .A(n426), .B(n425), .Z(n380) );
  INV_X1 U455 ( .A(KEYINPUT90), .ZN(n469) );
  NOR2_X1 U456 ( .A1(n557), .A2(n490), .ZN(n491) );
  XNOR2_X1 U457 ( .A(n427), .B(n380), .ZN(n428) );
  INV_X1 U458 ( .A(KEYINPUT2), .ZN(n578) );
  XNOR2_X1 U459 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U460 ( .A(n429), .B(n428), .ZN(n602) );
  XNOR2_X1 U461 ( .A(n431), .B(KEYINPUT13), .ZN(n534) );
  XOR2_X2 U462 ( .A(G143), .B(G128), .Z(n457) );
  XOR2_X1 U463 ( .A(KEYINPUT69), .B(G131), .Z(n424) );
  XOR2_X1 U464 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n386) );
  NOR2_X1 U465 ( .A1(G953), .A2(G237), .ZN(n419) );
  NAND2_X1 U466 ( .A1(n419), .A2(G210), .ZN(n385) );
  XOR2_X1 U467 ( .A(n386), .B(n385), .Z(n387) );
  INV_X1 U468 ( .A(G902), .ZN(n444) );
  NAND2_X1 U469 ( .A1(n593), .A2(n444), .ZN(n388) );
  XNOR2_X2 U470 ( .A(n388), .B(G472), .ZN(n542) );
  XNOR2_X1 U471 ( .A(n453), .B(KEYINPUT10), .ZN(n422) );
  XNOR2_X1 U472 ( .A(n422), .B(n468), .ZN(n710) );
  XNOR2_X1 U473 ( .A(n391), .B(n390), .ZN(n395) );
  XNOR2_X1 U474 ( .A(KEYINPUT68), .B(KEYINPUT8), .ZN(n393) );
  XNOR2_X1 U475 ( .A(n393), .B(n392), .ZN(n434) );
  NAND2_X1 U476 ( .A1(n434), .A2(G221), .ZN(n394) );
  XNOR2_X1 U477 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U478 ( .A(n710), .B(n396), .ZN(n610) );
  XOR2_X1 U479 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n398) );
  XNOR2_X1 U480 ( .A(G902), .B(KEYINPUT15), .ZN(n580) );
  NAND2_X1 U481 ( .A1(n580), .A2(G234), .ZN(n397) );
  XNOR2_X1 U482 ( .A(n398), .B(n397), .ZN(n408) );
  AND2_X1 U483 ( .A1(n408), .A2(G217), .ZN(n400) );
  XNOR2_X1 U484 ( .A(KEYINPUT92), .B(KEYINPUT25), .ZN(n399) );
  XNOR2_X1 U485 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X2 U486 ( .A(n402), .B(n401), .ZN(n658) );
  NAND2_X1 U487 ( .A1(G234), .A2(G237), .ZN(n403) );
  XNOR2_X1 U488 ( .A(n403), .B(KEYINPUT14), .ZN(n488) );
  NOR2_X1 U489 ( .A1(n484), .A2(G900), .ZN(n404) );
  NAND2_X1 U490 ( .A1(n404), .A2(G902), .ZN(n405) );
  NAND2_X1 U491 ( .A1(n484), .A2(G952), .ZN(n486) );
  NAND2_X1 U492 ( .A1(n405), .A2(n486), .ZN(n406) );
  AND2_X1 U493 ( .A1(n488), .A2(n406), .ZN(n407) );
  XNOR2_X1 U494 ( .A(n407), .B(KEYINPUT81), .ZN(n546) );
  INV_X1 U495 ( .A(n546), .ZN(n411) );
  NAND2_X1 U496 ( .A1(n408), .A2(G221), .ZN(n410) );
  XNOR2_X1 U497 ( .A(KEYINPUT93), .B(KEYINPUT21), .ZN(n409) );
  XNOR2_X1 U498 ( .A(n410), .B(n409), .ZN(n657) );
  NAND2_X1 U499 ( .A1(n411), .A2(n657), .ZN(n412) );
  OR2_X2 U500 ( .A1(n658), .A2(n412), .ZN(n414) );
  INV_X1 U501 ( .A(KEYINPUT71), .ZN(n413) );
  INV_X1 U502 ( .A(KEYINPUT102), .ZN(n415) );
  XOR2_X1 U503 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n418) );
  XNOR2_X1 U504 ( .A(G122), .B(KEYINPUT97), .ZN(n417) );
  XNOR2_X1 U505 ( .A(n418), .B(n417), .ZN(n421) );
  NAND2_X1 U506 ( .A1(G214), .A2(n419), .ZN(n420) );
  XNOR2_X1 U507 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U508 ( .A(n423), .B(n422), .Z(n429) );
  XNOR2_X1 U509 ( .A(n424), .B(KEYINPUT11), .ZN(n427) );
  XNOR2_X1 U510 ( .A(n639), .B(G113), .ZN(n425) );
  NOR2_X1 U511 ( .A1(G902), .A2(n602), .ZN(n430) );
  XOR2_X1 U512 ( .A(G475), .B(n430), .Z(n431) );
  XNOR2_X1 U513 ( .A(KEYINPUT99), .B(G478), .ZN(n440) );
  XOR2_X1 U514 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n433) );
  XNOR2_X1 U515 ( .A(G107), .B(n448), .ZN(n432) );
  XNOR2_X1 U516 ( .A(n433), .B(n432), .ZN(n436) );
  NAND2_X1 U517 ( .A1(n434), .A2(G217), .ZN(n435) );
  XNOR2_X1 U518 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U519 ( .A(n438), .B(n437), .ZN(n615) );
  NOR2_X1 U520 ( .A1(G902), .A2(n615), .ZN(n439) );
  XNOR2_X1 U521 ( .A(n440), .B(n439), .ZN(n533) );
  NOR2_X1 U522 ( .A1(n534), .A2(n533), .ZN(n641) );
  NAND2_X1 U523 ( .A1(n441), .A2(n641), .ZN(n442) );
  XNOR2_X1 U524 ( .A(n442), .B(KEYINPUT103), .ZN(n445) );
  INV_X1 U525 ( .A(G237), .ZN(n443) );
  NAND2_X1 U526 ( .A1(n444), .A2(n443), .ZN(n460) );
  NAND2_X1 U527 ( .A1(n460), .A2(G214), .ZN(n668) );
  NAND2_X1 U528 ( .A1(n445), .A2(n668), .ZN(n570) );
  XNOR2_X1 U529 ( .A(G104), .B(G110), .ZN(n447) );
  XNOR2_X1 U530 ( .A(n472), .B(n702), .ZN(n459) );
  NAND2_X1 U531 ( .A1(n484), .A2(G224), .ZN(n451) );
  XNOR2_X1 U532 ( .A(n451), .B(KEYINPUT87), .ZN(n455) );
  XOR2_X1 U533 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n452) );
  XNOR2_X1 U534 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U535 ( .A(n459), .B(n458), .ZN(n585) );
  NAND2_X1 U536 ( .A1(n585), .A2(n580), .ZN(n464) );
  XOR2_X1 U537 ( .A(KEYINPUT80), .B(KEYINPUT88), .Z(n462) );
  NAND2_X1 U538 ( .A1(n460), .A2(G210), .ZN(n461) );
  XNOR2_X1 U539 ( .A(n462), .B(n461), .ZN(n463) );
  INV_X1 U540 ( .A(n563), .ZN(n573) );
  XOR2_X1 U541 ( .A(KEYINPUT105), .B(KEYINPUT36), .Z(n465) );
  XNOR2_X1 U542 ( .A(n466), .B(n465), .ZN(n477) );
  NAND2_X1 U543 ( .A1(n484), .A2(G227), .ZN(n467) );
  XNOR2_X1 U544 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U545 ( .A(n474), .B(n473), .ZN(n622) );
  NOR2_X1 U546 ( .A1(G902), .A2(n622), .ZN(n476) );
  INV_X1 U547 ( .A(G469), .ZN(n475) );
  XNOR2_X2 U548 ( .A(n476), .B(n475), .ZN(n553) );
  XNOR2_X2 U549 ( .A(n553), .B(KEYINPUT1), .ZN(n509) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(KEYINPUT111), .Z(n478) );
  XOR2_X1 U551 ( .A(n478), .B(G125), .Z(n479) );
  XNOR2_X1 U552 ( .A(n567), .B(n479), .ZN(G27) );
  INV_X1 U553 ( .A(n533), .ZN(n480) );
  NAND2_X1 U554 ( .A1(n480), .A2(n534), .ZN(n671) );
  INV_X1 U555 ( .A(n671), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n657), .B(KEYINPUT94), .ZN(n508) );
  NAND2_X1 U557 ( .A1(n481), .A2(n668), .ZN(n483) );
  XOR2_X1 U558 ( .A(KEYINPUT19), .B(KEYINPUT66), .Z(n482) );
  XNOR2_X1 U559 ( .A(n483), .B(n482), .ZN(n557) );
  NOR2_X1 U560 ( .A1(n484), .A2(G898), .ZN(n485) );
  XOR2_X1 U561 ( .A(KEYINPUT89), .B(n485), .Z(n705) );
  NAND2_X1 U562 ( .A1(n705), .A2(G902), .ZN(n487) );
  AND2_X1 U563 ( .A1(n487), .A2(n486), .ZN(n489) );
  INV_X1 U564 ( .A(n488), .ZN(n683) );
  OR2_X1 U565 ( .A1(n489), .A2(n683), .ZN(n490) );
  OR2_X1 U566 ( .A1(n542), .A2(n658), .ZN(n495) );
  NOR2_X1 U567 ( .A1(n509), .A2(n495), .ZN(n496) );
  NAND2_X1 U568 ( .A1(n523), .A2(n496), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(G110), .ZN(G12) );
  INV_X1 U570 ( .A(n658), .ZN(n497) );
  NAND2_X1 U571 ( .A1(n509), .A2(n497), .ZN(n499) );
  XNOR2_X1 U572 ( .A(n520), .B(KEYINPUT79), .ZN(n498) );
  NOR2_X1 U573 ( .A1(n499), .A2(n498), .ZN(n500) );
  NAND2_X1 U574 ( .A1(n523), .A2(n500), .ZN(n502) );
  INV_X1 U575 ( .A(KEYINPUT32), .ZN(n501) );
  XNOR2_X1 U576 ( .A(n502), .B(n501), .ZN(n726) );
  INV_X1 U577 ( .A(n503), .ZN(n504) );
  INV_X1 U578 ( .A(KEYINPUT44), .ZN(n517) );
  NAND2_X1 U579 ( .A1(n517), .A2(KEYINPUT84), .ZN(n505) );
  XNOR2_X1 U580 ( .A(n506), .B(n505), .ZN(n515) );
  INV_X1 U581 ( .A(n507), .ZN(n528) );
  AND2_X1 U582 ( .A1(n658), .A2(n508), .ZN(n526) );
  NOR2_X1 U583 ( .A1(n528), .A2(n687), .ZN(n510) );
  XNOR2_X1 U584 ( .A(n510), .B(n353), .ZN(n513) );
  INV_X1 U585 ( .A(n534), .ZN(n511) );
  NAND2_X1 U586 ( .A1(n533), .A2(n511), .ZN(n561) );
  INV_X1 U587 ( .A(n561), .ZN(n512) );
  NAND2_X1 U588 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U589 ( .A(n514), .B(KEYINPUT35), .ZN(n516) );
  INV_X1 U590 ( .A(n516), .ZN(n723) );
  NAND2_X1 U591 ( .A1(n515), .A2(n723), .ZN(n519) );
  NAND2_X1 U592 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U593 ( .A1(n519), .A2(n518), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n520), .A2(n658), .ZN(n521) );
  NOR2_X1 U595 ( .A1(n509), .A2(n521), .ZN(n522) );
  NAND2_X1 U596 ( .A1(n523), .A2(n522), .ZN(n525) );
  INV_X1 U597 ( .A(KEYINPUT100), .ZN(n524) );
  XNOR2_X1 U598 ( .A(n525), .B(n524), .ZN(n727) );
  INV_X1 U599 ( .A(n727), .ZN(n537) );
  INV_X1 U600 ( .A(n553), .ZN(n527) );
  INV_X1 U601 ( .A(n526), .ZN(n652) );
  NOR2_X1 U602 ( .A1(n527), .A2(n652), .ZN(n548) );
  NOR2_X1 U603 ( .A1(n542), .A2(n528), .ZN(n529) );
  NAND2_X1 U604 ( .A1(n548), .A2(n529), .ZN(n629) );
  XOR2_X1 U605 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n532) );
  INV_X1 U606 ( .A(n542), .ZN(n655) );
  NOR2_X1 U607 ( .A1(n530), .A2(n655), .ZN(n665) );
  NAND2_X1 U608 ( .A1(n665), .A2(n507), .ZN(n531) );
  XNOR2_X1 U609 ( .A(n532), .B(n531), .ZN(n646) );
  NAND2_X1 U610 ( .A1(n629), .A2(n646), .ZN(n535) );
  INV_X1 U611 ( .A(n641), .ZN(n643) );
  AND2_X1 U612 ( .A1(n534), .A2(n533), .ZN(n635) );
  INV_X1 U613 ( .A(n635), .ZN(n645) );
  NAND2_X1 U614 ( .A1(n643), .A2(n645), .ZN(n673) );
  NAND2_X1 U615 ( .A1(n535), .A2(n673), .ZN(n536) );
  AND2_X1 U616 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U617 ( .A1(n539), .A2(n538), .ZN(n541) );
  INV_X1 U618 ( .A(KEYINPUT45), .ZN(n540) );
  XNOR2_X1 U619 ( .A(n541), .B(n540), .ZN(n698) );
  NAND2_X1 U620 ( .A1(n668), .A2(n542), .ZN(n544) );
  XOR2_X2 U621 ( .A(n563), .B(KEYINPUT38), .Z(n669) );
  XNOR2_X1 U622 ( .A(n549), .B(KEYINPUT40), .ZN(n725) );
  NAND2_X1 U623 ( .A1(n669), .A2(n668), .ZN(n674) );
  XNOR2_X1 U624 ( .A(n550), .B(KEYINPUT41), .ZN(n686) );
  NOR2_X1 U625 ( .A1(n551), .A2(n655), .ZN(n552) );
  XNOR2_X1 U626 ( .A(n552), .B(KEYINPUT28), .ZN(n554) );
  NAND2_X1 U627 ( .A1(n554), .A2(n553), .ZN(n558) );
  NOR2_X1 U628 ( .A1(n686), .A2(n558), .ZN(n555) );
  XNOR2_X1 U629 ( .A(n555), .B(KEYINPUT42), .ZN(n724) );
  NAND2_X1 U630 ( .A1(n640), .A2(n673), .ZN(n559) );
  NOR2_X1 U631 ( .A1(KEYINPUT67), .A2(n559), .ZN(n560) );
  XNOR2_X1 U632 ( .A(KEYINPUT47), .B(n560), .ZN(n565) );
  NOR2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n564) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n638) );
  NAND2_X1 U635 ( .A1(n565), .A2(n638), .ZN(n566) );
  XNOR2_X1 U636 ( .A(KEYINPUT70), .B(KEYINPUT48), .ZN(n568) );
  NAND2_X1 U637 ( .A1(n569), .A2(n635), .ZN(n648) );
  INV_X1 U638 ( .A(n648), .ZN(n575) );
  INV_X1 U639 ( .A(n570), .ZN(n571) );
  INV_X1 U640 ( .A(n509), .ZN(n653) );
  NAND2_X1 U641 ( .A1(n571), .A2(n653), .ZN(n572) );
  XNOR2_X1 U642 ( .A(n572), .B(KEYINPUT43), .ZN(n574) );
  AND2_X1 U643 ( .A1(n574), .A2(n573), .ZN(n649) );
  NOR2_X1 U644 ( .A1(n575), .A2(n649), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n713) );
  NOR2_X2 U646 ( .A1(n698), .A2(n713), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n579), .B(n578), .ZN(n651) );
  INV_X1 U648 ( .A(n580), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n651), .A2(n581), .ZN(n583) );
  INV_X1 U650 ( .A(KEYINPUT64), .ZN(n582) );
  XNOR2_X2 U651 ( .A(n583), .B(n582), .ZN(n608) );
  NAND2_X1 U652 ( .A1(n608), .A2(G210), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n584) );
  XNOR2_X1 U654 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n587), .B(n586), .ZN(n589) );
  INV_X1 U656 ( .A(G952), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n588), .A2(G953), .ZN(n613) );
  NAND2_X1 U658 ( .A1(n589), .A2(n613), .ZN(n591) );
  XOR2_X1 U659 ( .A(KEYINPUT82), .B(KEYINPUT56), .Z(n590) );
  XNOR2_X1 U660 ( .A(n591), .B(n590), .ZN(G51) );
  NAND2_X1 U661 ( .A1(n608), .A2(G472), .ZN(n595) );
  XOR2_X1 U662 ( .A(KEYINPUT85), .B(KEYINPUT62), .Z(n592) );
  XNOR2_X1 U663 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n595), .B(n594), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n596), .A2(n613), .ZN(n599) );
  XNOR2_X1 U666 ( .A(KEYINPUT106), .B(KEYINPUT63), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n597), .B(KEYINPUT86), .ZN(n598) );
  XNOR2_X1 U668 ( .A(n599), .B(n598), .ZN(G57) );
  NAND2_X1 U669 ( .A1(n608), .A2(G475), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT65), .B(KEYINPUT120), .ZN(n600) );
  XOR2_X1 U671 ( .A(n600), .B(KEYINPUT59), .Z(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U673 ( .A(n604), .B(n603), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n605), .A2(n613), .ZN(n607) );
  INV_X1 U675 ( .A(KEYINPUT60), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(G60) );
  NAND2_X1 U677 ( .A1(n618), .A2(G217), .ZN(n612) );
  XOR2_X1 U678 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n609) );
  XNOR2_X1 U679 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U681 ( .A(n613), .ZN(n625) );
  NOR2_X1 U682 ( .A1(n614), .A2(n625), .ZN(G66) );
  NAND2_X1 U683 ( .A1(n618), .A2(G478), .ZN(n616) );
  XNOR2_X1 U684 ( .A(n616), .B(n615), .ZN(n617) );
  NOR2_X1 U685 ( .A1(n617), .A2(n625), .ZN(G63) );
  NAND2_X1 U686 ( .A1(n618), .A2(G469), .ZN(n624) );
  XOR2_X1 U687 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n620) );
  XNOR2_X1 U688 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(n621) );
  XOR2_X1 U690 ( .A(n622), .B(n621), .Z(n623) );
  XNOR2_X1 U691 ( .A(n624), .B(n623), .ZN(n626) );
  NOR2_X1 U692 ( .A1(n626), .A2(n625), .ZN(G54) );
  NOR2_X1 U693 ( .A1(n643), .A2(n629), .ZN(n627) );
  XOR2_X1 U694 ( .A(KEYINPUT108), .B(n627), .Z(n628) );
  XNOR2_X1 U695 ( .A(G104), .B(n628), .ZN(G6) );
  NOR2_X1 U696 ( .A1(n645), .A2(n629), .ZN(n634) );
  XOR2_X1 U697 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n631) );
  XNOR2_X1 U698 ( .A(G107), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U700 ( .A(KEYINPUT27), .B(n632), .ZN(n633) );
  XNOR2_X1 U701 ( .A(n634), .B(n633), .ZN(G9) );
  XOR2_X1 U702 ( .A(G128), .B(KEYINPUT29), .Z(n637) );
  NAND2_X1 U703 ( .A1(n635), .A2(n640), .ZN(n636) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(G30) );
  XNOR2_X1 U705 ( .A(n639), .B(n638), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U707 ( .A(n642), .B(G146), .ZN(G48) );
  NOR2_X1 U708 ( .A1(n646), .A2(n643), .ZN(n644) );
  XOR2_X1 U709 ( .A(G113), .B(n644), .Z(G15) );
  NOR2_X1 U710 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U711 ( .A(G116), .B(n647), .Z(G18) );
  XNOR2_X1 U712 ( .A(G134), .B(n648), .ZN(G36) );
  XOR2_X1 U713 ( .A(G140), .B(n649), .Z(n650) );
  XNOR2_X1 U714 ( .A(KEYINPUT112), .B(n650), .ZN(G42) );
  BUF_X1 U715 ( .A(n651), .Z(n692) );
  NAND2_X1 U716 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U717 ( .A(n654), .B(KEYINPUT50), .ZN(n656) );
  NAND2_X1 U718 ( .A1(n656), .A2(n655), .ZN(n663) );
  XOR2_X1 U719 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n660) );
  NOR2_X1 U720 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U721 ( .A(n660), .B(n659), .Z(n661) );
  XNOR2_X1 U722 ( .A(n661), .B(KEYINPUT114), .ZN(n662) );
  NOR2_X1 U723 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U724 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U725 ( .A(KEYINPUT51), .B(n666), .Z(n667) );
  NOR2_X1 U726 ( .A1(n344), .A2(n667), .ZN(n680) );
  NOR2_X1 U727 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U728 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U729 ( .A(KEYINPUT115), .B(n672), .Z(n677) );
  INV_X1 U730 ( .A(n673), .ZN(n675) );
  NOR2_X1 U731 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U732 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U733 ( .A1(n687), .A2(n678), .ZN(n679) );
  NOR2_X1 U734 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U735 ( .A(n681), .B(KEYINPUT116), .ZN(n682) );
  XNOR2_X1 U736 ( .A(n682), .B(KEYINPUT52), .ZN(n684) );
  NOR2_X1 U737 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U738 ( .A1(G952), .A2(n685), .ZN(n690) );
  NOR2_X1 U739 ( .A1(n687), .A2(n344), .ZN(n688) );
  NOR2_X1 U740 ( .A1(n688), .A2(G953), .ZN(n689) );
  NAND2_X1 U741 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U742 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U743 ( .A(n693), .B(KEYINPUT117), .Z(n694) );
  XNOR2_X1 U744 ( .A(KEYINPUT53), .B(n694), .ZN(G75) );
  NAND2_X1 U745 ( .A1(G953), .A2(G224), .ZN(n695) );
  XNOR2_X1 U746 ( .A(KEYINPUT61), .B(n695), .ZN(n696) );
  NAND2_X1 U747 ( .A1(n696), .A2(G898), .ZN(n697) );
  XNOR2_X1 U748 ( .A(n697), .B(KEYINPUT123), .ZN(n700) );
  NOR2_X1 U749 ( .A1(n698), .A2(G953), .ZN(n699) );
  NOR2_X1 U750 ( .A1(n700), .A2(n699), .ZN(n707) );
  XNOR2_X1 U751 ( .A(G101), .B(n701), .ZN(n703) );
  XNOR2_X1 U752 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U753 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U754 ( .A(n707), .B(n706), .Z(n708) );
  XNOR2_X1 U755 ( .A(KEYINPUT124), .B(n708), .ZN(G69) );
  XOR2_X1 U756 ( .A(KEYINPUT4), .B(KEYINPUT90), .Z(n709) );
  XNOR2_X1 U757 ( .A(n710), .B(n709), .ZN(n711) );
  XNOR2_X1 U758 ( .A(n712), .B(n711), .ZN(n716) );
  XOR2_X1 U759 ( .A(n716), .B(n713), .Z(n714) );
  NOR2_X1 U760 ( .A1(n714), .A2(G953), .ZN(n715) );
  XNOR2_X1 U761 ( .A(n715), .B(KEYINPUT125), .ZN(n722) );
  XNOR2_X1 U762 ( .A(n716), .B(G227), .ZN(n717) );
  XNOR2_X1 U763 ( .A(n717), .B(KEYINPUT126), .ZN(n718) );
  NAND2_X1 U764 ( .A1(n718), .A2(G900), .ZN(n719) );
  XOR2_X1 U765 ( .A(KEYINPUT127), .B(n719), .Z(n720) );
  NAND2_X1 U766 ( .A1(n720), .A2(G953), .ZN(n721) );
  NAND2_X1 U767 ( .A1(n722), .A2(n721), .ZN(G72) );
  XNOR2_X1 U768 ( .A(n723), .B(G122), .ZN(G24) );
  XOR2_X1 U769 ( .A(n724), .B(G137), .Z(G39) );
  XOR2_X1 U770 ( .A(n725), .B(G131), .Z(G33) );
  XOR2_X1 U771 ( .A(G119), .B(n726), .Z(G21) );
  XNOR2_X1 U772 ( .A(G101), .B(KEYINPUT107), .ZN(n728) );
  XNOR2_X1 U773 ( .A(n728), .B(n727), .ZN(G3) );
endmodule

