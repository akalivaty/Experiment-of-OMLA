

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XOR2_X1 U319 ( .A(G99GAT), .B(G85GAT), .Z(n380) );
  XNOR2_X1 U320 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U321 ( .A(n419), .B(KEYINPUT36), .ZN(n578) );
  XNOR2_X1 U322 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U323 ( .A(n454), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U324 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U325 ( .A(KEYINPUT0), .B(KEYINPUT77), .Z(n288) );
  XNOR2_X1 U326 ( .A(G120GAT), .B(G127GAT), .ZN(n287) );
  XNOR2_X1 U327 ( .A(n288), .B(n287), .ZN(n289) );
  XOR2_X1 U328 ( .A(n289), .B(G134GAT), .Z(n291) );
  XNOR2_X1 U329 ( .A(G113GAT), .B(KEYINPUT76), .ZN(n290) );
  XNOR2_X1 U330 ( .A(n291), .B(n290), .ZN(n318) );
  XOR2_X1 U331 ( .A(G190GAT), .B(G99GAT), .Z(n293) );
  XNOR2_X1 U332 ( .A(KEYINPUT83), .B(KEYINPUT20), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U334 ( .A(n318), .B(n294), .Z(n296) );
  NAND2_X1 U335 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U336 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U337 ( .A(G176GAT), .B(G43GAT), .Z(n298) );
  XNOR2_X1 U338 ( .A(G169GAT), .B(G15GAT), .ZN(n297) );
  XNOR2_X1 U339 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U340 ( .A(n300), .B(n299), .Z(n309) );
  XNOR2_X1 U341 ( .A(KEYINPUT18), .B(KEYINPUT80), .ZN(n301) );
  XNOR2_X1 U342 ( .A(n301), .B(G183GAT), .ZN(n302) );
  XOR2_X1 U343 ( .A(n302), .B(KEYINPUT81), .Z(n304) );
  XNOR2_X1 U344 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n303) );
  XNOR2_X1 U345 ( .A(n304), .B(n303), .ZN(n341) );
  XOR2_X1 U346 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n306) );
  XNOR2_X1 U347 ( .A(G71GAT), .B(KEYINPUT82), .ZN(n305) );
  XNOR2_X1 U348 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U349 ( .A(n341), .B(n307), .ZN(n308) );
  XOR2_X1 U350 ( .A(n309), .B(n308), .Z(n495) );
  INV_X1 U351 ( .A(n495), .ZN(n527) );
  XOR2_X1 U352 ( .A(G162GAT), .B(G85GAT), .Z(n311) );
  NAND2_X1 U353 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n314) );
  XOR2_X1 U355 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n313) );
  XNOR2_X1 U356 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n441) );
  XOR2_X1 U358 ( .A(n314), .B(n441), .Z(n320) );
  XOR2_X1 U359 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n316) );
  XNOR2_X1 U360 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n315) );
  XNOR2_X1 U361 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U362 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U363 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U364 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n322) );
  XNOR2_X1 U365 ( .A(G57GAT), .B(KEYINPUT93), .ZN(n321) );
  XNOR2_X1 U366 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U367 ( .A(G148GAT), .B(G29GAT), .Z(n324) );
  XNOR2_X1 U368 ( .A(G1GAT), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U369 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U370 ( .A(n326), .B(n325), .Z(n327) );
  XOR2_X1 U371 ( .A(n328), .B(n327), .Z(n514) );
  INV_X1 U372 ( .A(n514), .ZN(n489) );
  XOR2_X1 U373 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n330) );
  XNOR2_X1 U374 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U375 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U376 ( .A(G197GAT), .B(n331), .Z(n450) );
  XOR2_X1 U377 ( .A(G169GAT), .B(G8GAT), .Z(n349) );
  XOR2_X1 U378 ( .A(KEYINPUT95), .B(KEYINPUT98), .Z(n333) );
  XNOR2_X1 U379 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n332) );
  XNOR2_X1 U380 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U381 ( .A(n349), .B(n334), .Z(n336) );
  NAND2_X1 U382 ( .A1(G226GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U383 ( .A(n336), .B(n335), .ZN(n339) );
  XOR2_X1 U384 ( .A(G64GAT), .B(G204GAT), .Z(n338) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G92GAT), .ZN(n337) );
  XNOR2_X1 U386 ( .A(n338), .B(n337), .ZN(n370) );
  XOR2_X1 U387 ( .A(n339), .B(n370), .Z(n343) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(G190GAT), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n340), .B(G218GAT), .ZN(n391) );
  XNOR2_X1 U390 ( .A(n341), .B(n391), .ZN(n342) );
  XNOR2_X1 U391 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U392 ( .A(n450), .B(n344), .Z(n517) );
  INV_X1 U393 ( .A(n517), .ZN(n493) );
  INV_X1 U394 ( .A(KEYINPUT113), .ZN(n376) );
  XOR2_X1 U395 ( .A(KEYINPUT65), .B(G197GAT), .Z(n346) );
  XNOR2_X1 U396 ( .A(G50GAT), .B(G36GAT), .ZN(n345) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n359) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G43GAT), .Z(n348) );
  XNOR2_X1 U399 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n392) );
  XOR2_X1 U401 ( .A(n392), .B(n349), .Z(n351) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U404 ( .A(G113GAT), .B(KEYINPUT66), .Z(n353) );
  XNOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n352) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U407 ( .A(n355), .B(n354), .Z(n357) );
  XOR2_X1 U408 ( .A(G15GAT), .B(G1GAT), .Z(n402) );
  XOR2_X1 U409 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XNOR2_X1 U410 ( .A(n402), .B(n432), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U412 ( .A(n359), .B(n358), .ZN(n552) );
  XOR2_X1 U413 ( .A(G78GAT), .B(G148GAT), .Z(n361) );
  XNOR2_X1 U414 ( .A(G106GAT), .B(KEYINPUT68), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n442) );
  XNOR2_X1 U416 ( .A(G71GAT), .B(G57GAT), .ZN(n362) );
  XNOR2_X1 U417 ( .A(n362), .B(KEYINPUT13), .ZN(n401) );
  XNOR2_X1 U418 ( .A(n442), .B(n401), .ZN(n374) );
  XNOR2_X1 U419 ( .A(KEYINPUT67), .B(KEYINPUT69), .ZN(n364) );
  XNOR2_X1 U420 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n380), .B(n365), .ZN(n367) );
  NAND2_X1 U423 ( .A1(G230GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n369) );
  INV_X1 U425 ( .A(KEYINPUT33), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n370), .B(KEYINPUT32), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n569) );
  XOR2_X1 U430 ( .A(n569), .B(KEYINPUT41), .Z(n557) );
  NAND2_X1 U431 ( .A1(n552), .A2(n557), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n377), .B(KEYINPUT46), .ZN(n417) );
  XOR2_X1 U434 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n379) );
  XNOR2_X1 U435 ( .A(G134GAT), .B(KEYINPUT70), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n398) );
  XNOR2_X1 U437 ( .A(n380), .B(G92GAT), .ZN(n386) );
  XNOR2_X1 U438 ( .A(G50GAT), .B(G162GAT), .ZN(n431) );
  NAND2_X1 U439 ( .A1(KEYINPUT10), .A2(n431), .ZN(n384) );
  INV_X1 U440 ( .A(KEYINPUT10), .ZN(n382) );
  XOR2_X1 U441 ( .A(G50GAT), .B(G162GAT), .Z(n381) );
  NAND2_X1 U442 ( .A1(n382), .A2(n381), .ZN(n383) );
  NAND2_X1 U443 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U445 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n388) );
  XNOR2_X1 U446 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n387) );
  XOR2_X1 U447 ( .A(n388), .B(n387), .Z(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n392), .B(n391), .ZN(n394) );
  NAND2_X1 U450 ( .A1(G232GAT), .A2(G233GAT), .ZN(n393) );
  XOR2_X1 U451 ( .A(n398), .B(n397), .Z(n549) );
  INV_X1 U452 ( .A(n549), .ZN(n419) );
  XOR2_X1 U453 ( .A(G78GAT), .B(G211GAT), .Z(n400) );
  XNOR2_X1 U454 ( .A(G22GAT), .B(G183GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n415) );
  XOR2_X1 U456 ( .A(n401), .B(G64GAT), .Z(n404) );
  XNOR2_X1 U457 ( .A(n402), .B(G8GAT), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U459 ( .A(KEYINPUT14), .B(G155GAT), .Z(n406) );
  NAND2_X1 U460 ( .A1(G231GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U461 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U462 ( .A(n408), .B(n407), .Z(n413) );
  XOR2_X1 U463 ( .A(KEYINPUT15), .B(KEYINPUT75), .Z(n410) );
  XNOR2_X1 U464 ( .A(KEYINPUT12), .B(KEYINPUT74), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U466 ( .A(G127GAT), .B(n411), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U468 ( .A(n415), .B(n414), .Z(n534) );
  AND2_X1 U469 ( .A1(n419), .A2(n534), .ZN(n416) );
  AND2_X1 U470 ( .A1(n417), .A2(n416), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n418), .B(KEYINPUT47), .ZN(n425) );
  NOR2_X1 U472 ( .A1(n578), .A2(n534), .ZN(n420) );
  XOR2_X1 U473 ( .A(n420), .B(KEYINPUT45), .Z(n421) );
  NOR2_X1 U474 ( .A1(n569), .A2(n421), .ZN(n422) );
  XNOR2_X1 U475 ( .A(KEYINPUT114), .B(n422), .ZN(n423) );
  INV_X1 U476 ( .A(n552), .ZN(n566) );
  NAND2_X1 U477 ( .A1(n423), .A2(n566), .ZN(n424) );
  NAND2_X1 U478 ( .A1(n425), .A2(n424), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n426), .B(KEYINPUT48), .ZN(n541) );
  NAND2_X1 U480 ( .A1(n493), .A2(n541), .ZN(n428) );
  XNOR2_X1 U481 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n427) );
  XOR2_X1 U482 ( .A(n428), .B(n427), .Z(n429) );
  NOR2_X1 U483 ( .A1(n489), .A2(n429), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n430), .B(KEYINPUT64), .ZN(n565) );
  XOR2_X1 U485 ( .A(n381), .B(G204GAT), .Z(n434) );
  XNOR2_X1 U486 ( .A(n432), .B(G218GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n446) );
  XOR2_X1 U488 ( .A(KEYINPUT86), .B(KEYINPUT90), .Z(n436) );
  XNOR2_X1 U489 ( .A(KEYINPUT84), .B(KEYINPUT91), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U491 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n438) );
  XNOR2_X1 U492 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U494 ( .A(n440), .B(n439), .Z(n444) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U497 ( .A(n446), .B(n445), .Z(n448) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U500 ( .A(n450), .B(n449), .ZN(n462) );
  NAND2_X1 U501 ( .A1(n565), .A2(n462), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X2 U504 ( .A1(n527), .A2(n453), .ZN(n560) );
  NAND2_X1 U505 ( .A1(n560), .A2(n549), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n454) );
  XOR2_X1 U507 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n474) );
  NOR2_X1 U508 ( .A1(n549), .A2(n534), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT16), .ZN(n470) );
  XOR2_X1 U510 ( .A(KEYINPUT27), .B(n517), .Z(n464) );
  NAND2_X1 U511 ( .A1(n464), .A2(n489), .ZN(n543) );
  XNOR2_X1 U512 ( .A(KEYINPUT28), .B(n462), .ZN(n521) );
  INV_X1 U513 ( .A(n521), .ZN(n500) );
  NOR2_X1 U514 ( .A1(n543), .A2(n500), .ZN(n525) );
  NAND2_X1 U515 ( .A1(n527), .A2(n525), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT99), .B(n458), .Z(n469) );
  NAND2_X1 U517 ( .A1(n495), .A2(n493), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n459), .A2(n462), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n460), .Z(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT100), .ZN(n466) );
  NOR2_X1 U521 ( .A1(n462), .A2(n495), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n463), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U523 ( .A1(n464), .A2(n564), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U525 ( .A1(n514), .A2(n467), .ZN(n468) );
  NAND2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n482) );
  NAND2_X1 U527 ( .A1(n470), .A2(n482), .ZN(n471) );
  XNOR2_X1 U528 ( .A(KEYINPUT101), .B(n471), .ZN(n503) );
  NOR2_X1 U529 ( .A1(n566), .A2(n569), .ZN(n486) );
  NAND2_X1 U530 ( .A1(n503), .A2(n486), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT102), .B(n472), .Z(n480) );
  NAND2_X1 U532 ( .A1(n480), .A2(n489), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U534 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n480), .A2(n493), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U538 ( .A1(n480), .A2(n495), .ZN(n477) );
  XNOR2_X1 U539 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n479), .ZN(G1326GAT) );
  NAND2_X1 U541 ( .A1(n480), .A2(n500), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n481), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT107), .B(KEYINPUT39), .Z(n491) );
  XOR2_X1 U544 ( .A(KEYINPUT106), .B(KEYINPUT38), .Z(n488) );
  NAND2_X1 U545 ( .A1(n534), .A2(n482), .ZN(n483) );
  NOR2_X1 U546 ( .A1(n578), .A2(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(KEYINPUT105), .B(KEYINPUT37), .ZN(n484) );
  XNOR2_X1 U548 ( .A(n485), .B(n484), .ZN(n513) );
  NAND2_X1 U549 ( .A1(n513), .A2(n486), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n499) );
  NAND2_X1 U551 ( .A1(n499), .A2(n489), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U553 ( .A(G29GAT), .B(n492), .Z(G1328GAT) );
  NAND2_X1 U554 ( .A1(n493), .A2(n499), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n497) );
  NAND2_X1 U557 ( .A1(n499), .A2(n495), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U559 ( .A(G43GAT), .B(n498), .Z(G1330GAT) );
  NAND2_X1 U560 ( .A1(n500), .A2(n499), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(G50GAT), .ZN(G1331GAT) );
  NAND2_X1 U562 ( .A1(n557), .A2(n566), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT109), .ZN(n512) );
  NAND2_X1 U564 ( .A1(n503), .A2(n512), .ZN(n508) );
  NOR2_X1 U565 ( .A1(n514), .A2(n508), .ZN(n504) );
  XOR2_X1 U566 ( .A(n504), .B(KEYINPUT42), .Z(n505) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(n505), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n517), .A2(n508), .ZN(n506) );
  XOR2_X1 U569 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U570 ( .A1(n527), .A2(n508), .ZN(n507) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n521), .A2(n508), .ZN(n510) );
  XNOR2_X1 U573 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n513), .A2(n512), .ZN(n520) );
  NOR2_X1 U577 ( .A1(n514), .A2(n520), .ZN(n516) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n517), .A2(n520), .ZN(n518) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n518), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n527), .A2(n520), .ZN(n519) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n519), .Z(G1338GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U585 ( .A(KEYINPUT112), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  NAND2_X1 U588 ( .A1(n541), .A2(n525), .ZN(n526) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U590 ( .A(KEYINPUT115), .B(n528), .Z(n538) );
  NAND2_X1 U591 ( .A1(n538), .A2(n552), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n531) );
  NAND2_X1 U594 ( .A1(n538), .A2(n557), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT116), .Z(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n536) );
  INV_X1 U599 ( .A(n534), .ZN(n574) );
  NAND2_X1 U600 ( .A1(n538), .A2(n574), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(G127GAT), .B(n537), .Z(G1342GAT) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U604 ( .A1(n538), .A2(n549), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n541), .A2(n564), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n552), .A2(n550), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n544), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U611 ( .A1(n550), .A2(n557), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n574), .A2(n550), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U618 ( .A1(n552), .A2(n560), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U623 ( .A(KEYINPUT121), .B(n556), .Z(n559) );
  NAND2_X1 U624 ( .A1(n560), .A2(n557), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U626 ( .A1(n574), .A2(n560), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n563) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n577) );
  NOR2_X1 U632 ( .A1(n566), .A2(n577), .ZN(n567) );
  XOR2_X1 U633 ( .A(n568), .B(n567), .Z(G1352GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n571) );
  INV_X1 U635 ( .A(n577), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n573), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G211GAT), .B(n576), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

