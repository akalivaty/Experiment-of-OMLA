//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT66), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT68), .B(KEYINPUT69), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  XOR2_X1   g041(.A(KEYINPUT3), .B(G2104), .Z(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n462), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT71), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G2105), .B1(new_n471), .B2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n461), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n477), .B(new_n480), .C1(G124), .C2(new_n482), .ZN(G162));
  INV_X1    g058(.A(G126), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n486));
  OAI22_X1  g061(.A1(new_n481), .A2(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n462), .A2(G138), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(KEYINPUT72), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n461), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n461), .A2(new_n488), .ZN(new_n492));
  INV_X1    g067(.A(new_n490), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n487), .B1(new_n491), .B2(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n499), .A2(KEYINPUT76), .A3(G543), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT76), .B1(new_n499), .B2(G543), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G62), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT73), .B(G651), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT73), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT6), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n509), .B2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT74), .A4(KEYINPUT6), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n502), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G88), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  NAND2_X1  g097(.A1(G50), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n521), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AOI211_X1 g100(.A(KEYINPUT75), .B(new_n523), .C1(new_n517), .C2(new_n518), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n520), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n520), .B(new_n529), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n508), .B1(new_n528), .B2(new_n530), .ZN(G166));
  AOI21_X1  g106(.A(new_n515), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n532));
  AND4_X1   g107(.A1(KEYINPUT74), .A2(new_n510), .A3(new_n512), .A4(KEYINPUT6), .ZN(new_n533));
  OAI21_X1  g108(.A(KEYINPUT78), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT78), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n517), .A2(new_n535), .A3(new_n518), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(G543), .A3(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G51), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT7), .Z(new_n541));
  NOR2_X1   g116(.A1(new_n499), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n543), .B1(new_n497), .B2(KEYINPUT5), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n499), .A2(KEYINPUT76), .A3(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g121(.A1(new_n546), .A2(G63), .A3(G651), .ZN(new_n547));
  AOI211_X1 g122(.A(new_n541), .B(new_n547), .C1(G89), .C2(new_n519), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n539), .A2(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  AOI21_X1  g125(.A(new_n497), .B1(new_n522), .B2(KEYINPUT78), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n551), .A2(G52), .A3(new_n536), .ZN(new_n552));
  NAND2_X1  g127(.A1(G77), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G64), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n502), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n519), .A2(G90), .B1(new_n555), .B2(new_n506), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G301));
  INV_X1    g132(.A(G301), .ZN(G171));
  OAI211_X1 g133(.A(G56), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n505), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(G81), .B2(new_n519), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n534), .A2(G43), .A3(G543), .A4(new_n536), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT80), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND4_X1  g147(.A1(new_n534), .A2(G53), .A3(G543), .A4(new_n536), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n551), .A2(new_n575), .A3(G53), .A4(new_n536), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n546), .A2(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(G78), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n509), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n522), .A2(new_n546), .ZN(new_n581));
  INV_X1    g156(.A(G91), .ZN(new_n582));
  OAI21_X1  g157(.A(KEYINPUT81), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT81), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n519), .A2(new_n584), .A3(G91), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n580), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n577), .A2(new_n586), .ZN(G299));
  OAI21_X1  g162(.A(new_n524), .B1(new_n532), .B2(new_n533), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT75), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n522), .A2(new_n521), .A3(new_n524), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n529), .B1(new_n591), .B2(new_n520), .ZN(new_n592));
  INV_X1    g167(.A(new_n530), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n507), .B1(new_n592), .B2(new_n593), .ZN(G303));
  NAND4_X1  g169(.A1(new_n534), .A2(G49), .A3(G543), .A4(new_n536), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n546), .B2(G74), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT82), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  OAI211_X1 g173(.A(new_n598), .B(G651), .C1(new_n546), .C2(G74), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n519), .A2(G87), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n595), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT83), .ZN(G288));
  NAND2_X1  g178(.A1(new_n546), .A2(G61), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n604), .A2(new_n605), .B1(G73), .B2(G543), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n546), .A2(KEYINPUT84), .A3(G61), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(new_n506), .ZN(new_n609));
  NAND2_X1  g184(.A1(G48), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G86), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n502), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(new_n522), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(G305));
  NAND2_X1  g189(.A1(new_n519), .A2(G85), .ZN(new_n615));
  AOI22_X1  g190(.A1(new_n546), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G47), .ZN(new_n617));
  OAI221_X1 g192(.A(new_n615), .B1(new_n505), .B2(new_n616), .C1(new_n537), .C2(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n522), .A2(G92), .A3(new_n546), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n519), .A2(KEYINPUT10), .A3(G92), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n502), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n622), .A2(new_n623), .B1(G651), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n538), .A2(G54), .ZN(new_n628));
  AND2_X1   g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n619), .B1(new_n629), .B2(G868), .ZN(G284));
  OAI21_X1  g205(.A(new_n619), .B1(new_n629), .B2(G868), .ZN(G321));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(G299), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n632), .B2(G168), .ZN(G280));
  XNOR2_X1  g209(.A(G280), .B(KEYINPUT85), .ZN(G297));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g215(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g216(.A1(new_n471), .A2(new_n461), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT12), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n482), .A2(G123), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n478), .A2(G135), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n462), .A2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n646), .A2(new_n647), .A3(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(KEYINPUT14), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT15), .B(G2435), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2438), .ZN(new_n657));
  XOR2_X1   g232(.A(G2427), .B(G2430), .Z(new_n658));
  AOI21_X1  g233(.A(new_n655), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n657), .B2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2451), .B(G2454), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n660), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(G14), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2084), .B(G2090), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT87), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n671), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(new_n645), .ZN(new_n679));
  NOR2_X1   g254(.A1(G2072), .A2(G2078), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n442), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G2096), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n679), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1961), .B(G1966), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n686), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT20), .Z(new_n693));
  AOI211_X1 g268(.A(new_n691), .B(new_n693), .C1(new_n686), .C2(new_n690), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT88), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n695), .B(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(G229));
  AOI22_X1  g277(.A1(new_n478), .A2(G141), .B1(new_n471), .B2(G105), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT26), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n482), .B2(G129), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G29), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n709), .B2(G32), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT27), .B(G1996), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT89), .B(G29), .ZN(new_n714));
  NOR2_X1   g289(.A1(G164), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G27), .B2(new_n714), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n713), .B1(G2078), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(G286), .A2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G21), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n709), .A2(G33), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT25), .ZN(new_n728));
  NAND2_X1  g303(.A1(G115), .A2(G2104), .ZN(new_n729));
  INV_X1    g304(.A(G127), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n467), .B2(new_n730), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n731), .A2(G2105), .B1(new_n478), .B2(G139), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT95), .B(G2072), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n736), .A2(G34), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(G34), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n714), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n473), .B2(new_n709), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  OAI22_X1  g316(.A1(new_n734), .A2(new_n735), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n741), .B2(new_n740), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT31), .B(G11), .Z(new_n744));
  INV_X1    g319(.A(G28), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n745), .A2(KEYINPUT30), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT96), .ZN(new_n747));
  AOI21_X1  g322(.A(G29), .B1(new_n745), .B2(KEYINPUT30), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n749), .B1(new_n652), .B2(new_n714), .C1(new_n717), .C2(G2078), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n734), .B2(new_n735), .ZN(new_n751));
  NAND4_X1  g326(.A1(new_n718), .A2(new_n724), .A3(new_n743), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G171), .A2(new_n720), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G5), .B2(new_n720), .ZN(new_n754));
  INV_X1    g329(.A(G1961), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n722), .A2(new_n723), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n754), .A2(new_n755), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n756), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  OR3_X1    g334(.A1(new_n752), .A2(KEYINPUT97), .A3(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(KEYINPUT97), .B1(new_n752), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n720), .A2(G20), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT23), .Z(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G299), .B2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1956), .ZN(new_n765));
  NOR2_X1   g340(.A1(G4), .A2(G16), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n629), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n714), .A2(G35), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT98), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G162), .B2(new_n714), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT29), .B(G2090), .Z(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n565), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G16), .B2(G19), .ZN(new_n775));
  INV_X1    g350(.A(G1341), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n714), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n482), .A2(G128), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n478), .A2(G140), .ZN(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n779), .B1(new_n785), .B2(new_n709), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n773), .A2(new_n777), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n775), .A2(new_n776), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n768), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n760), .A2(new_n761), .A3(new_n765), .A4(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n505), .B1(new_n606), .B2(new_n607), .ZN(new_n793));
  INV_X1    g368(.A(new_n613), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n795), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G6), .B2(G16), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT32), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(KEYINPUT32), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G1981), .ZN(new_n801));
  INV_X1    g376(.A(G1981), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n798), .A2(new_n802), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G23), .ZN(new_n805));
  AND4_X1   g380(.A1(KEYINPUT92), .A2(new_n595), .A3(new_n600), .A4(new_n601), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n597), .A2(new_n599), .B1(new_n519), .B2(G87), .ZN(new_n807));
  AOI21_X1  g382(.A(KEYINPUT92), .B1(new_n807), .B2(new_n595), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n805), .B1(new_n809), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n804), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n720), .A2(G22), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G166), .B2(new_n720), .ZN(new_n816));
  INV_X1    g391(.A(G1971), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n813), .A2(new_n814), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n812), .A4(new_n804), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  INV_X1    g399(.A(new_n714), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(G25), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n482), .A2(G119), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n478), .A2(G131), .ZN(new_n828));
  OR2_X1    g403(.A1(G95), .A2(G2105), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n829), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n826), .B1(new_n832), .B2(new_n825), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT90), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT91), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n720), .B1(G290), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n837), .B2(G290), .ZN(new_n839));
  INV_X1    g414(.A(G24), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(G16), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n836), .B1(new_n841), .B2(G1986), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G1986), .B2(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n822), .A2(new_n824), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT36), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT36), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n822), .A2(new_n824), .A3(new_n846), .A4(new_n843), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n792), .B1(new_n845), .B2(new_n847), .ZN(G311));
  INV_X1    g423(.A(G311), .ZN(G150));
  OAI211_X1 g424(.A(G67), .B(new_n498), .C1(new_n500), .C2(new_n501), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n519), .A2(G93), .B1(new_n852), .B2(new_n506), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n534), .A2(G55), .A3(G543), .A4(new_n536), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(G860), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT37), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n629), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT38), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n564), .A2(new_n855), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n562), .A2(new_n853), .A3(new_n563), .A4(new_n854), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n859), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  AOI21_X1  g443(.A(G860), .B1(new_n863), .B2(new_n864), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n857), .B1(new_n870), .B2(new_n871), .ZN(G145));
  XNOR2_X1  g447(.A(new_n733), .B(new_n707), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n643), .B(new_n831), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n876));
  INV_X1    g451(.A(new_n491), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n490), .B1(new_n461), .B2(new_n488), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n494), .A2(KEYINPUT101), .A3(new_n491), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n487), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n784), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n478), .A2(G142), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n462), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n482), .A2(new_n886), .A3(G130), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n482), .B2(G130), .ZN(new_n888));
  OAI221_X1 g463(.A(new_n883), .B1(new_n884), .B2(new_n885), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n882), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n875), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(G162), .B(new_n652), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n473), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(KEYINPUT103), .Z(new_n895));
  AOI21_X1  g470(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g473(.A(G868), .B1(new_n853), .B2(new_n854), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(KEYINPUT105), .ZN(new_n900));
  XOR2_X1   g475(.A(new_n638), .B(new_n862), .Z(new_n901));
  NAND2_X1  g476(.A1(new_n627), .A2(new_n628), .ZN(new_n902));
  NAND2_X1  g477(.A1(G299), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n577), .A2(new_n586), .A3(new_n627), .A4(new_n628), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT104), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  AND4_X1   g486(.A1(new_n577), .A2(new_n586), .A3(new_n627), .A4(new_n628), .ZN(new_n912));
  AOI22_X1  g487(.A1(new_n577), .A2(new_n586), .B1(new_n627), .B2(new_n628), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n903), .A2(KEYINPUT41), .A3(new_n904), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n901), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n910), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n910), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(G290), .B(new_n795), .ZN(new_n922));
  NOR2_X1   g497(.A1(G303), .A2(new_n809), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT92), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n602), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n807), .A2(KEYINPUT92), .A3(new_n595), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(G166), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n922), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(G290), .B(G305), .ZN(new_n930));
  NAND2_X1  g505(.A1(G303), .A2(new_n809), .ZN(new_n931));
  NAND2_X1  g506(.A1(G166), .A2(new_n927), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n632), .B1(new_n921), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n918), .A2(new_n936), .A3(new_n920), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n900), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n920), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n919), .B1(new_n910), .B2(new_n916), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  AND4_X1   g516(.A1(KEYINPUT105), .A2(new_n941), .A3(new_n937), .A4(G868), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n938), .A2(new_n942), .ZN(G295));
  NOR2_X1   g518(.A1(new_n938), .A2(new_n942), .ZN(G331));
  AND3_X1   g519(.A1(new_n860), .A2(G301), .A3(new_n861), .ZN(new_n945));
  AOI21_X1  g520(.A(G301), .B1(new_n860), .B2(new_n861), .ZN(new_n946));
  OAI21_X1  g521(.A(G286), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND4_X1   g522(.A1(new_n563), .A2(new_n562), .A3(new_n853), .A4(new_n854), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n563), .A2(new_n562), .B1(new_n853), .B2(new_n854), .ZN(new_n949));
  OAI21_X1  g524(.A(G171), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n860), .A2(G301), .A3(new_n861), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(G168), .A3(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n947), .A2(new_n914), .A3(new_n915), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n905), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n945), .A2(new_n946), .A3(G286), .ZN(new_n955));
  AOI21_X1  g530(.A(G168), .B1(new_n950), .B2(new_n951), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n934), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n934), .A2(new_n957), .A3(new_n953), .A4(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n957), .A2(new_n953), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n936), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G37), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n962), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT43), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n955), .A2(new_n956), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n953), .B1(new_n909), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(G37), .B1(new_n973), .B2(new_n936), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n962), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT108), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n962), .A2(new_n977), .A3(new_n974), .A4(new_n971), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n970), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n962), .A2(new_n974), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n980), .B1(new_n983), .B2(KEYINPUT43), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n962), .A2(new_n967), .A3(new_n971), .A4(new_n968), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n982), .A2(new_n987), .A3(KEYINPUT44), .A4(new_n985), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n981), .B1(new_n986), .B2(new_n988), .ZN(G397));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n707), .B(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n784), .B(new_n787), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n832), .A2(new_n834), .ZN(new_n994));
  OAI22_X1  g569(.A1(new_n993), .A2(new_n994), .B1(G2067), .B2(new_n784), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n881), .B2(G1384), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n465), .A2(new_n472), .A3(G40), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n999), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n1001), .A2(G1986), .A3(G290), .ZN(new_n1002));
  XOR2_X1   g577(.A(new_n1002), .B(KEYINPUT127), .Z(new_n1003));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n831), .B(new_n834), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n1006), .B(KEYINPUT110), .Z(new_n1007));
  OAI21_X1  g582(.A(new_n999), .B1(new_n1007), .B2(new_n993), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1000), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1001), .B1(new_n708), .B2(new_n992), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT125), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT46), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n1001), .B2(G1996), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n999), .A2(KEYINPUT46), .A3(new_n990), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT126), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1018), .A2(KEYINPUT47), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(KEYINPUT47), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1011), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G8), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(new_n881), .B2(G1384), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n485), .A2(new_n486), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1025), .B1(new_n482), .B2(G126), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n877), .A2(new_n876), .A3(new_n878), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT101), .B1(new_n494), .B2(new_n491), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(KEYINPUT112), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT45), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n494), .A2(new_n491), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n1026), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n998), .B1(KEYINPUT45), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n723), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1024), .A2(new_n1031), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1034), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n998), .B1(new_n1040), .B2(KEYINPUT50), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n741), .A3(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1022), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(G286), .A2(G8), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OR3_X1    g621(.A1(new_n1043), .A2(KEYINPUT122), .A3(new_n1046), .ZN(new_n1047));
  XOR2_X1   g622(.A(new_n1044), .B(KEYINPUT121), .Z(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT51), .B1(new_n1048), .B2(new_n1043), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT122), .B1(new_n1043), .B2(new_n1046), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1047), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1042), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT112), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n881), .A2(new_n1023), .A3(G1384), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n996), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G1966), .B1(new_n1055), .B2(new_n1035), .ZN(new_n1056));
  OAI211_X1 g631(.A(G8), .B(G286), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1051), .A2(new_n1060), .A3(new_n1057), .ZN(new_n1061));
  INV_X1    g636(.A(new_n998), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1024), .A2(new_n1031), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1976), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(G8), .C1(new_n927), .C2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT52), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT114), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(KEYINPUT114), .A3(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1065), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT52), .B1(G288), .B2(new_n1064), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n1068), .A2(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n609), .A2(new_n802), .A3(new_n613), .ZN(new_n1074));
  OAI21_X1  g649(.A(G1981), .B1(new_n793), .B2(new_n794), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n802), .B1(new_n609), .B2(new_n613), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n793), .A2(G1981), .A3(new_n794), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1077), .A2(G8), .A3(new_n1063), .A4(new_n1081), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1076), .A2(KEYINPUT115), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1073), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1081), .A2(G8), .A3(new_n1063), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1083), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1085), .A2(new_n1086), .A3(KEYINPUT116), .A4(new_n1077), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n881), .A2(G1384), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT45), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n998), .B1(new_n1040), .B2(new_n996), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n817), .ZN(new_n1093));
  INV_X1    g668(.A(G2090), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1039), .A2(new_n1094), .A3(new_n1041), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1022), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT55), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(G166), .B2(new_n1022), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n1100));
  AND3_X1   g675(.A1(new_n1097), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1100), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1096), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1038), .B1(new_n1024), .B2(new_n1031), .ZN(new_n1104));
  NOR4_X1   g679(.A1(G164), .A2(KEYINPUT117), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT117), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1062), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1104), .A2(new_n1108), .A3(G2090), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1093), .ZN(new_n1110));
  OAI21_X1  g685(.A(G8), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1072), .A2(new_n1088), .A3(new_n1103), .A4(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n755), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n1092), .B2(G2078), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(G2078), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1055), .A2(new_n1035), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(G171), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1114), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1059), .A2(new_n1061), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1063), .A2(G8), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OR2_X1    g701(.A1(G288), .A2(G1976), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1126), .B1(new_n1128), .B2(new_n1080), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1103), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(new_n1088), .A3(new_n1072), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1043), .A2(G168), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1114), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1043), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1096), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1136), .B1(new_n1112), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(new_n1088), .A3(new_n1072), .A4(new_n1103), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1132), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT56), .B(G2072), .ZN(new_n1141));
  AND3_X1   g716(.A1(new_n1090), .A2(new_n1091), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n577), .A2(new_n586), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1144), .B1(new_n577), .B2(new_n586), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(G1956), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1143), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1063), .A2(G2067), .ZN(new_n1152));
  AOI21_X1  g727(.A(G1348), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1151), .B(new_n629), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT119), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1147), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1145), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1107), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1034), .A2(new_n1106), .A3(new_n1038), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n998), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT50), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1162));
  AOI21_X1  g737(.A(G1956), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1155), .B(new_n1158), .C1(new_n1163), .C2(new_n1142), .ZN(new_n1164));
  AND2_X1   g739(.A1(new_n1154), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(G1348), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1115), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1152), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT60), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT120), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1153), .A2(new_n1152), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT60), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT60), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1174), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1170), .A2(new_n1173), .A3(new_n629), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n629), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1172), .B1(new_n1171), .B2(KEYINPUT60), .ZN(new_n1178));
  NOR4_X1   g753(.A1(new_n1153), .A2(new_n1152), .A3(KEYINPUT120), .A4(new_n1174), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1143), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1148), .B1(new_n1150), .B2(new_n1143), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1164), .A2(KEYINPUT61), .A3(new_n1151), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT58), .B(G1341), .Z(new_n1188));
  AOI22_X1  g763(.A1(new_n1187), .A2(new_n990), .B1(new_n1063), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g764(.A(KEYINPUT59), .B1(new_n1189), .B2(new_n564), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1063), .A2(new_n1188), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1191), .B1(G1996), .B2(new_n1092), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1192), .A2(new_n1193), .A3(new_n565), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1185), .A2(new_n1186), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1165), .B1(new_n1181), .B2(new_n1196), .ZN(new_n1197));
  AND3_X1   g772(.A1(new_n997), .A2(KEYINPUT123), .A3(new_n1062), .ZN(new_n1198));
  AOI21_X1  g773(.A(KEYINPUT123), .B1(new_n997), .B2(new_n1062), .ZN(new_n1199));
  OAI211_X1 g774(.A(new_n1090), .B(new_n1119), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1200), .A2(new_n1116), .A3(new_n1118), .A4(G301), .ZN(new_n1201));
  AOI21_X1  g776(.A(KEYINPUT54), .B1(new_n1122), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1114), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1116), .A2(new_n1118), .A3(new_n1120), .A4(G301), .ZN(new_n1204));
  OR2_X1    g779(.A1(new_n1204), .A2(KEYINPUT124), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1204), .A2(KEYINPUT124), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1200), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(G171), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1205), .A2(KEYINPUT54), .A3(new_n1206), .A4(new_n1208), .ZN(new_n1209));
  NAND4_X1  g784(.A1(new_n1197), .A2(new_n1058), .A3(new_n1203), .A4(new_n1209), .ZN(new_n1210));
  AND3_X1   g785(.A1(new_n1124), .A2(new_n1140), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g786(.A(G290), .B(G1986), .Z(new_n1212));
  OAI21_X1  g787(.A(new_n1008), .B1(new_n1001), .B2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT111), .ZN(new_n1214));
  OAI21_X1  g789(.A(new_n1021), .B1(new_n1211), .B2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g790(.A(G319), .B1(new_n668), .B2(new_n669), .ZN(new_n1217));
  NOR3_X1   g791(.A1(G229), .A2(G227), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n979), .A2(new_n897), .A3(new_n1218), .ZN(G225));
  INV_X1    g793(.A(G225), .ZN(G308));
endmodule


