//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n798, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(KEYINPUT73), .A2(KEYINPUT1), .ZN(new_n206));
  NOR2_X1   g005(.A1(G127gat), .A2(G134gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G127gat), .A2(G134gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI221_X1 g008(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(KEYINPUT1), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n206), .B1(new_n208), .B2(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT27), .B(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n216), .B(new_n217), .C1(KEYINPUT70), .C2(KEYINPUT28), .ZN(new_n221));
  NAND2_X1  g020(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT71), .ZN(new_n225));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(KEYINPUT26), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n232), .A2(KEYINPUT71), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n224), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n215), .B1(new_n223), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n232), .A2(KEYINPUT71), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n237), .B(new_n229), .C1(KEYINPUT26), .C2(new_n230), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n236), .A2(KEYINPUT72), .A3(new_n224), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n224), .B1(KEYINPUT68), .B2(KEYINPUT24), .ZN(new_n242));
  AND2_X1   g041(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n243));
  OAI221_X1 g042(.A(new_n241), .B1(G183gat), .B2(G190gat), .C1(new_n242), .C2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n245), .B1(new_n230), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n226), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n227), .A2(KEYINPUT23), .B1(new_n226), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n244), .A2(new_n247), .A3(new_n249), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n224), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT64), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n256), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n241), .A2(KEYINPUT64), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n260));
  INV_X1    g059(.A(G176gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n260), .A2(KEYINPUT23), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n248), .B1(new_n230), .B2(new_n246), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n245), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT66), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n268), .A3(new_n245), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n253), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n240), .B1(new_n270), .B2(KEYINPUT69), .ZN(new_n271));
  INV_X1    g070(.A(new_n269), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n265), .B2(new_n245), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n252), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n214), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G227gat), .ZN(new_n278));
  INV_X1    g077(.A(G233gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n275), .ZN(new_n282));
  INV_X1    g081(.A(new_n214), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .A4(new_n240), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n277), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n205), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT34), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n277), .A2(new_n284), .ZN(new_n289));
  INV_X1    g088(.A(new_n280), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g090(.A(KEYINPUT34), .B(new_n280), .C1(new_n277), .C2(new_n284), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n287), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n287), .A2(new_n291), .A3(new_n292), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n296));
  INV_X1    g095(.A(new_n285), .ZN(new_n297));
  OAI22_X1  g096(.A1(new_n294), .A2(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(G228gat), .A2(G233gat), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G141gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n305), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(KEYINPUT79), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT79), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(G155gat), .B2(G162gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n308), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT80), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT80), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n307), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  NOR2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n304), .B(new_n306), .C1(new_n308), .C2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327));
  INV_X1    g126(.A(KEYINPUT22), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n328), .A2(KEYINPUT74), .B1(G211gat), .B2(G218gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT22), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(KEYINPUT75), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G197gat), .B(G204gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT75), .B1(new_n329), .B2(new_n331), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n335), .ZN(new_n337));
  INV_X1    g136(.A(new_n327), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(new_n338), .A3(new_n332), .A4(new_n333), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n336), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n326), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n318), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n317), .B1(new_n307), .B2(new_n314), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n322), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n324), .B1(new_n336), .B2(new_n339), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT3), .B1(new_n346), .B2(KEYINPUT84), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT84), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n348), .B1(new_n340), .B2(new_n324), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n345), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n341), .B1(new_n350), .B2(KEYINPUT85), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT85), .ZN(new_n352));
  AOI211_X1 g151(.A(new_n352), .B(new_n345), .C1(new_n347), .C2(new_n349), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n299), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G22gat), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n320), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(new_n344), .ZN(new_n357));
  OR2_X1    g156(.A1(new_n357), .A2(KEYINPUT86), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(KEYINPUT86), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n299), .B1(new_n326), .B2(new_n340), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n355), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(KEYINPUT31), .B(G50gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n354), .A2(KEYINPUT88), .A3(new_n361), .A4(new_n355), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n367), .A2(KEYINPUT87), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n361), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(G22gat), .ZN(new_n373));
  AOI211_X1 g172(.A(new_n355), .B(new_n370), .C1(new_n354), .C2(new_n361), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n362), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n291), .A2(new_n292), .ZN(new_n376));
  INV_X1    g175(.A(new_n287), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n297), .A2(new_n296), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n379), .A3(new_n293), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n298), .A2(new_n369), .A3(new_n375), .A4(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n214), .B(new_n322), .C1(new_n342), .C2(new_n343), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n319), .A2(new_n384), .A3(new_n322), .A4(new_n214), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n323), .A3(new_n283), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n344), .A2(new_n283), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n382), .ZN(new_n393));
  INV_X1    g192(.A(new_n389), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  INV_X1    g199(.A(KEYINPUT81), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n385), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n383), .A2(new_n401), .A3(new_n385), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n394), .A2(KEYINPUT5), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n402), .A2(new_n403), .A3(new_n388), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n396), .A2(new_n400), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT6), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n396), .A2(new_n405), .ZN(new_n411));
  INV_X1    g210(.A(new_n400), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n406), .A2(KEYINPUT82), .A3(new_n407), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n413), .A2(new_n407), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n410), .A2(KEYINPUT83), .A3(new_n413), .A4(new_n414), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n281), .A2(new_n282), .A3(new_n240), .ZN(new_n422));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n423), .B(KEYINPUT76), .Z(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n340), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n236), .A2(new_n224), .A3(new_n238), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n274), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n423), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n425), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n423), .B1(new_n274), .B2(new_n427), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n325), .B1(new_n271), .B2(new_n276), .ZN(new_n434));
  INV_X1    g233(.A(new_n424), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n432), .B1(new_n436), .B2(new_n426), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT78), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n437), .A2(KEYINPUT78), .A3(new_n441), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n432), .B(new_n440), .C1(new_n436), .C2(new_n426), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT30), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n424), .B1(new_n422), .B2(new_n325), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n340), .B1(new_n448), .B2(new_n433), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n432), .A4(new_n440), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n444), .A2(new_n445), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n421), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT35), .B1(new_n381), .B2(new_n453), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n443), .B(new_n440), .C1(new_n449), .C2(new_n432), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT78), .B1(new_n437), .B2(new_n441), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g256(.A1(new_n447), .A2(new_n451), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT35), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n378), .A2(new_n379), .A3(new_n293), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n379), .B1(new_n378), .B2(new_n293), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n375), .A2(new_n369), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT89), .B1(new_n411), .B2(new_n412), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT89), .ZN(new_n465));
  AOI211_X1 g264(.A(new_n465), .B(new_n400), .C1(new_n396), .C2(new_n405), .ZN(new_n466));
  NOR3_X1   g265(.A1(new_n464), .A2(new_n466), .A3(new_n408), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT90), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n418), .B1(new_n467), .B2(KEYINPUT90), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n459), .A2(new_n462), .A3(new_n463), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n402), .A2(new_n403), .A3(new_n388), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n394), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n400), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT39), .B1(new_n393), .B2(new_n394), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n473), .B2(new_n394), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT40), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n400), .A4(new_n475), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n464), .B(new_n466), .C1(new_n479), .C2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n457), .B2(new_n458), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n441), .B1(new_n437), .B2(KEYINPUT37), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n449), .B2(new_n432), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT38), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n441), .A2(KEYINPUT37), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n442), .A2(new_n489), .ZN(new_n490));
  AND2_X1   g289(.A1(new_n425), .A2(new_n431), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n486), .B1(new_n491), .B2(new_n340), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n426), .B1(new_n448), .B2(new_n433), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n488), .A2(new_n495), .A3(new_n446), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n463), .B(new_n484), .C1(new_n496), .C2(new_n470), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n375), .A2(new_n369), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n453), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n460), .B2(new_n461), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n298), .A2(KEYINPUT36), .A3(new_n380), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n472), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(G1gat), .ZN(new_n506));
  INV_X1    g305(.A(G15gat), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(G22gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n355), .A2(G15gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(G8gat), .B1(new_n510), .B2(KEYINPUT94), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n506), .A2(KEYINPUT93), .A3(KEYINPUT16), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT16), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(G1gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n512), .A2(new_n513), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n510), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n517), .B(new_n510), .C1(KEYINPUT94), .C2(G8gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT95), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  INV_X1    g322(.A(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G36gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(new_n525), .A3(KEYINPUT14), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n527), .B1(G29gat), .B2(G36gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT15), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT15), .A4(new_n529), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n526), .A2(new_n529), .ZN(new_n536));
  XOR2_X1   g335(.A(G43gat), .B(G50gat), .Z(new_n537));
  NAND4_X1  g336(.A1(new_n536), .A2(KEYINPUT15), .A3(new_n528), .A4(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(new_n522), .B(new_n523), .C1(new_n535), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n523), .ZN(new_n540));
  NAND2_X1  g339(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n541));
  AND4_X1   g340(.A1(new_n535), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n521), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n530), .A2(new_n531), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n533), .A2(new_n534), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n520), .A3(new_n519), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n543), .A2(KEYINPUT18), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(new_n544), .B(KEYINPUT13), .Z(new_n550));
  INV_X1    g349(.A(new_n548), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n520), .B2(new_n519), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n547), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n535), .A2(new_n538), .A3(new_n540), .A4(new_n541), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n551), .B1(new_n557), .B2(new_n521), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT18), .B1(new_n558), .B2(new_n544), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561));
  INV_X1    g360(.A(G197gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT11), .B(G169gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n560), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(KEYINPUT92), .B(new_n567), .C1(new_n554), .C2(new_n559), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n505), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G231gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n573), .A2(new_n279), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G57gat), .B(G64gat), .Z(new_n576));
  INV_X1    g375(.A(KEYINPUT9), .ZN(new_n577));
  INV_X1    g376(.A(G71gat), .ZN(new_n578));
  INV_X1    g377(.A(G78gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n576), .A2(new_n582), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n575), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AOI211_X1 g388(.A(new_n574), .B(new_n587), .C1(new_n584), .C2(new_n585), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G127gat), .B(G155gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT20), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n593), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n589), .B2(new_n590), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n521), .B1(new_n600), .B2(new_n586), .ZN(new_n601));
  XNOR2_X1  g400(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n598), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n594), .A2(new_n605), .A3(new_n596), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n599), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n604), .B1(new_n599), .B2(new_n606), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(G134gat), .B(G162gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G99gat), .B(G106gat), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n617));
  AND2_X1   g416(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n618), .A2(new_n619), .A3(G92gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT8), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n621), .B1(G99gat), .B2(G106gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n617), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  OR2_X1    g422(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n624));
  INV_X1    g423(.A(G92gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(KEYINPUT98), .A2(G85gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(G99gat), .ZN(new_n628));
  INV_X1    g427(.A(G106gat), .ZN(new_n629));
  OAI21_X1  g428(.A(KEYINPUT8), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G85gat), .A2(G92gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT7), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n616), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  AOI211_X1 g435(.A(new_n615), .B(new_n634), .C1(new_n623), .C2(new_n631), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n638), .A2(new_n547), .B1(KEYINPUT41), .B2(new_n610), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n627), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n640));
  AOI21_X1  g439(.A(KEYINPUT99), .B1(new_n627), .B2(new_n630), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n635), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n615), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n632), .A2(new_n616), .A3(new_n635), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n557), .A2(KEYINPUT100), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT100), .B1(new_n557), .B2(new_n645), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G190gat), .B(G218gat), .Z(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n650), .ZN(new_n652));
  INV_X1    g451(.A(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n646), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n654), .B2(new_n639), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n614), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n649), .A2(new_n650), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n652), .A3(new_n639), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n613), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n609), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n586), .B1(new_n636), .B2(new_n637), .ZN(new_n664));
  INV_X1    g463(.A(new_n586), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n643), .A2(new_n665), .A3(new_n644), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n664), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n638), .A2(KEYINPUT10), .A3(new_n665), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n663), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n661), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(G120gat), .B(G148gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT102), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n661), .B(new_n676), .C1(new_n670), .C2(new_n671), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n660), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n421), .A2(KEYINPUT104), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n421), .A2(KEYINPUT104), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n572), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(new_n506), .ZN(G1324gat));
  NOR3_X1   g487(.A1(new_n572), .A2(new_n452), .A3(new_n682), .ZN(new_n689));
  INV_X1    g488(.A(G8gat), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  XOR2_X1   g491(.A(KEYINPUT16), .B(G8gat), .Z(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n692), .A2(KEYINPUT105), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n693), .B2(new_n697), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n691), .A2(new_n694), .B1(new_n689), .B2(new_n698), .ZN(G1325gat));
  NOR2_X1   g498(.A1(new_n572), .A2(new_n682), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(new_n507), .A3(new_n462), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n572), .A2(new_n503), .A3(new_n682), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n701), .B1(new_n507), .B2(new_n702), .ZN(G1326gat));
  INV_X1    g502(.A(new_n682), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n505), .A2(new_n498), .A3(new_n571), .A4(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(KEYINPUT106), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n708), .B(new_n710), .ZN(G1327gat));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712));
  INV_X1    g511(.A(new_n571), .ZN(new_n713));
  INV_X1    g512(.A(new_n609), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n713), .A2(new_n714), .A3(new_n680), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716));
  INV_X1    g515(.A(new_n659), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n613), .B1(new_n657), .B2(new_n658), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n716), .B1(new_n505), .B2(new_n719), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n502), .A2(new_n501), .B1(new_n453), .B2(new_n498), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(new_n497), .B1(new_n454), .B2(new_n471), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n717), .B2(new_n718), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n656), .A2(KEYINPUT107), .A3(new_n659), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n716), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n722), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n715), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n712), .B1(new_n729), .B2(new_n686), .ZN(new_n730));
  INV_X1    g529(.A(new_n715), .ZN(new_n731));
  INV_X1    g530(.A(new_n719), .ZN(new_n732));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n722), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n505), .A2(new_n716), .A3(new_n726), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n731), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n735), .A2(KEYINPUT108), .A3(new_n685), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n730), .A2(G29gat), .A3(new_n736), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n722), .A2(new_n732), .A3(new_n731), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n738), .A2(new_n524), .A3(new_n685), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n740), .ZN(G1328gat));
  OAI21_X1  g540(.A(G36gat), .B1(new_n729), .B2(new_n452), .ZN(new_n742));
  INV_X1    g541(.A(new_n452), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n525), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(KEYINPUT109), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n742), .B(new_n748), .C1(new_n746), .C2(new_n744), .ZN(G1329gat));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  INV_X1    g549(.A(G43gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n503), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n735), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n462), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(G43gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n750), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G43gat), .B1(new_n729), .B2(new_n503), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(KEYINPUT47), .A3(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1330gat));
  INV_X1    g560(.A(KEYINPUT48), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(KEYINPUT110), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n498), .B(new_n715), .C1(new_n720), .C2(new_n728), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G50gat), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n463), .A2(G50gat), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n505), .A2(new_n719), .A3(new_n715), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(KEYINPUT110), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n764), .B1(new_n766), .B2(new_n771), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n763), .B(new_n770), .C1(new_n765), .C2(G50gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(G1331gat));
  NAND3_X1  g573(.A1(new_n660), .A2(new_n713), .A3(new_n680), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n722), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n685), .A2(KEYINPUT111), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT111), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n683), .B2(new_n684), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g582(.A(new_n452), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n785), .A2(KEYINPUT112), .ZN(new_n788));
  OAI22_X1  g587(.A1(new_n787), .A2(new_n788), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  INV_X1    g588(.A(new_n788), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n791), .A3(new_n786), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1333gat));
  NAND3_X1  g592(.A1(new_n776), .A2(new_n578), .A3(new_n462), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n722), .A2(new_n503), .A3(new_n775), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n578), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g596(.A1(new_n776), .A2(new_n498), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g598(.A1(new_n714), .A2(new_n571), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n681), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n803), .B1(new_n733), .B2(new_n734), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n685), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n624), .A2(new_n626), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n505), .A2(new_n719), .A3(new_n800), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n505), .A2(KEYINPUT51), .A3(new_n719), .A4(new_n800), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n686), .A2(new_n806), .A3(new_n681), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n807), .A2(new_n814), .ZN(G1336gat));
  NOR3_X1   g614(.A1(new_n452), .A2(G92gat), .A3(new_n681), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n743), .B(new_n802), .C1(new_n720), .C2(new_n728), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G92gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n816), .B(KEYINPUT113), .Z(new_n822));
  AOI22_X1  g621(.A1(new_n812), .A2(new_n822), .B1(new_n818), .B2(G92gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n823), .B2(new_n820), .ZN(G1337gat));
  XOR2_X1   g623(.A(KEYINPUT114), .B(G99gat), .Z(new_n825));
  NAND4_X1  g624(.A1(new_n812), .A2(new_n462), .A3(new_n680), .A4(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n804), .A2(new_n752), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n827), .B2(new_n825), .ZN(G1338gat));
  AOI21_X1  g627(.A(new_n629), .B1(new_n804), .B2(new_n498), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n498), .A2(new_n629), .A3(new_n680), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT115), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n810), .B2(new_n811), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT53), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n833), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n802), .B1(new_n720), .B2(new_n728), .ZN(new_n836));
  OAI21_X1  g635(.A(G106gat), .B1(new_n836), .B2(new_n463), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n834), .A2(new_n839), .ZN(G1339gat));
  NAND3_X1  g639(.A1(new_n660), .A2(new_n713), .A3(new_n681), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n841), .B(KEYINPUT116), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n668), .A2(new_n663), .A3(new_n669), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n844), .A2(new_n670), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n668), .A2(new_n669), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(new_n845), .A3(new_n662), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n676), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n843), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  OR3_X1    g649(.A1(new_n670), .A2(new_n671), .A3(new_n676), .ZN(new_n851));
  INV_X1    g650(.A(new_n670), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n668), .A2(new_n663), .A3(new_n669), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n677), .B1(new_n670), .B2(new_n845), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(KEYINPUT55), .A3(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n571), .A2(new_n850), .A3(new_n851), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n554), .A2(new_n559), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n551), .A2(new_n552), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n544), .A2(new_n558), .B1(new_n859), .B2(new_n550), .ZN(new_n860));
  AOI22_X1  g659(.A1(new_n858), .A2(new_n568), .B1(new_n565), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n680), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n725), .A3(new_n724), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n861), .A2(new_n850), .A3(new_n851), .A4(new_n856), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n726), .A2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n842), .B1(new_n867), .B2(new_n714), .ZN(new_n868));
  INV_X1    g667(.A(new_n381), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n452), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(new_n780), .ZN(new_n871));
  AOI21_X1  g670(.A(G113gat), .B1(new_n871), .B2(new_n571), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n870), .B2(new_n686), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n714), .B1(new_n864), .B2(new_n866), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n841), .B(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n381), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n879), .A2(KEYINPUT117), .A3(new_n452), .A4(new_n685), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n874), .A2(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n571), .A2(G113gat), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n872), .B1(new_n881), .B2(new_n882), .ZN(G1340gat));
  NAND3_X1  g682(.A1(new_n874), .A2(new_n880), .A3(new_n680), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G120gat), .ZN(new_n885));
  INV_X1    g684(.A(G120gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n886), .A3(new_n680), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT118), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n885), .A2(new_n890), .A3(new_n887), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(G1341gat));
  INV_X1    g691(.A(G127gat), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n871), .A2(new_n893), .A3(new_n714), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n881), .A2(new_n714), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n893), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n874), .A2(new_n880), .A3(new_n719), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G134gat), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n452), .A2(new_n719), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n900), .A2(G134gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n781), .A2(new_n879), .A3(new_n901), .ZN(new_n902));
  XOR2_X1   g701(.A(new_n902), .B(KEYINPUT56), .Z(new_n903));
  NAND2_X1  g702(.A1(new_n898), .A2(KEYINPUT119), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(G1343gat));
  NAND3_X1  g704(.A1(new_n685), .A2(new_n452), .A3(new_n503), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n463), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n862), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n680), .A2(KEYINPUT120), .A3(new_n861), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n912), .A2(new_n857), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n732), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n714), .B1(new_n915), .B2(new_n866), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n877), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n914), .A2(new_n732), .B1(new_n726), .B2(new_n865), .ZN(new_n919));
  OAI21_X1  g718(.A(KEYINPUT121), .B1(new_n919), .B2(new_n714), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n910), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n868), .B2(new_n498), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(G141gat), .B1(new_n923), .B2(new_n713), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n777), .A2(new_n503), .A3(new_n779), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n498), .B1(new_n875), .B2(new_n877), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n925), .A2(new_n743), .A3(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n713), .A2(G141gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT58), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n866), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n932), .A2(new_n917), .A3(new_n609), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n933), .A2(new_n920), .A3(new_n842), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n934), .A2(new_n909), .B1(new_n908), .B2(new_n926), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n906), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n907), .B(KEYINPUT122), .C1(new_n921), .C2(new_n922), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n571), .A3(new_n937), .ZN(new_n938));
  AOI22_X1  g737(.A1(new_n938), .A2(G141gat), .B1(new_n927), .B2(new_n928), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n930), .B1(new_n939), .B2(new_n940), .ZN(G1344gat));
  NOR2_X1   g740(.A1(new_n302), .A2(KEYINPUT59), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n936), .A2(new_n937), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n681), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n868), .A2(new_n945), .A3(new_n909), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT123), .B1(new_n878), .B2(new_n910), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n865), .A2(new_n719), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n915), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n841), .B1(new_n950), .B2(new_n714), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT57), .B1(new_n951), .B2(new_n498), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n680), .B(new_n907), .C1(new_n948), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(G148gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(KEYINPUT59), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n944), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n927), .A2(new_n302), .A3(new_n680), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(G1345gat));
  OAI21_X1  g757(.A(G155gat), .B1(new_n943), .B2(new_n609), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n927), .A2(new_n309), .A3(new_n714), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1346gat));
  NAND3_X1  g760(.A1(new_n936), .A2(new_n726), .A3(new_n937), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT124), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n936), .A2(new_n937), .A3(new_n964), .A4(new_n726), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(G162gat), .A3(new_n965), .ZN(new_n966));
  OR4_X1    g765(.A1(G162gat), .A2(new_n925), .A3(new_n900), .A4(new_n926), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1347gat));
  NAND3_X1  g767(.A1(new_n780), .A2(new_n743), .A3(new_n879), .ZN(new_n969));
  OAI21_X1  g768(.A(G169gat), .B1(new_n969), .B2(new_n713), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n878), .A2(new_n685), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n743), .A3(new_n869), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n571), .A2(new_n260), .A3(new_n262), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1348gat));
  INV_X1    g773(.A(new_n972), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n261), .A3(new_n680), .ZN(new_n976));
  OAI21_X1  g775(.A(G176gat), .B1(new_n969), .B2(new_n681), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1349gat));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n216), .A3(new_n714), .ZN(new_n979));
  OAI21_X1  g778(.A(G183gat), .B1(new_n969), .B2(new_n609), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n981), .B(new_n982), .ZN(G1350gat));
  NAND3_X1  g782(.A1(new_n975), .A2(new_n217), .A3(new_n726), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n969), .A2(new_n732), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n985), .A2(new_n986), .A3(G190gat), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n985), .B2(G190gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n984), .B1(new_n987), .B2(new_n988), .ZN(G1351gat));
  AOI211_X1 g788(.A(new_n452), .B(new_n752), .C1(new_n777), .C2(new_n779), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n990), .B(new_n571), .C1(new_n948), .C2(new_n952), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT126), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n562), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n993), .B1(new_n992), .B2(new_n991), .ZN(new_n994));
  AND4_X1   g793(.A1(new_n498), .A2(new_n971), .A3(new_n743), .A4(new_n503), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(new_n562), .A3(new_n571), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1352gat));
  XNOR2_X1  g796(.A(KEYINPUT127), .B(G204gat), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n681), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  OR2_X1    g801(.A1(new_n948), .A2(new_n952), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1003), .A2(new_n680), .A3(new_n990), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1004), .A2(new_n998), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1002), .A2(new_n1005), .ZN(G1353gat));
  INV_X1    g805(.A(G211gat), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n995), .A2(new_n1007), .A3(new_n714), .ZN(new_n1008));
  OAI211_X1 g807(.A(new_n990), .B(new_n714), .C1(new_n948), .C2(new_n952), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1009), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(KEYINPUT63), .B1(new_n1009), .B2(G211gat), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(G1354gat));
  INV_X1    g811(.A(G218gat), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n995), .A2(new_n1013), .A3(new_n726), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1003), .A2(new_n719), .A3(new_n990), .ZN(new_n1015));
  INV_X1    g814(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1014), .B1(new_n1016), .B2(new_n1013), .ZN(G1355gat));
endmodule


