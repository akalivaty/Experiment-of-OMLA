//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0002(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AND2_X1   g0018(.A1(G107), .A2(G264), .ZN(new_n219));
  NOR4_X1   g0019(.A1(new_n212), .A2(new_n215), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n204), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(G58), .A2(G68), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n207), .B(new_n230), .C1(new_n233), .C2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(G226), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n214), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n213), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n231), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT66), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n256), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n259), .B1(new_n265), .B2(G226), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n266), .B(KEYINPUT67), .ZN(new_n267));
  AND2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT68), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT68), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G222), .ZN(new_n279));
  INV_X1    g0079(.A(G223), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n277), .B(new_n279), .C1(new_n280), .C2(new_n278), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n260), .A2(KEYINPUT69), .A3(new_n231), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT69), .ZN(new_n283));
  AND2_X1   g0083(.A1(G1), .A2(G13), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n281), .B(new_n287), .C1(G77), .C2(new_n277), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n267), .A2(G190), .A3(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(G20), .B1(new_n235), .B2(G50), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G150), .ZN(new_n292));
  XOR2_X1   g0092(.A(KEYINPUT8), .B(G58), .Z(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n232), .A2(G33), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n290), .B(new_n292), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n231), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT70), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n297), .A2(KEYINPUT70), .A3(new_n231), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G13), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G20), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n296), .A2(new_n303), .B1(new_n221), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n256), .A2(G20), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n302), .A2(G50), .A3(new_n306), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(KEYINPUT9), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n310), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT9), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n289), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n267), .B2(new_n288), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n289), .A2(KEYINPUT73), .A3(new_n311), .A4(new_n314), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n318), .A2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n259), .B1(new_n265), .B2(G244), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n277), .B1(new_n217), .B2(new_n278), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n227), .A2(G1698), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT71), .B(G107), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI22_X1  g0129(.A1(new_n326), .A2(new_n327), .B1(new_n277), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n287), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(G179), .ZN(new_n335));
  INV_X1    g0135(.A(new_n298), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n309), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n223), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n306), .A2(G77), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n293), .A2(new_n291), .B1(G20), .B2(G77), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT72), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n341), .B(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n340), .B1(new_n343), .B2(new_n295), .ZN(new_n344));
  AOI211_X1 g0144(.A(new_n338), .B(new_n339), .C1(new_n344), .C2(new_n298), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n334), .A2(new_n335), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n324), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n222), .A2(new_n278), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n227), .A2(G1698), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n277), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(G33), .A2(G97), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n331), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n259), .B1(new_n265), .B2(G238), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(KEYINPUT13), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n270), .A2(new_n276), .B1(new_n227), .B2(G1698), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n349), .B1(G33), .B2(G97), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n357), .B(new_n354), .C1(new_n359), .C2(new_n331), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n356), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n348), .B1(new_n361), .B2(G169), .ZN(new_n362));
  AOI211_X1 g0162(.A(KEYINPUT14), .B(new_n333), .C1(new_n356), .C2(new_n360), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G179), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n356), .A2(new_n360), .A3(KEYINPUT74), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n367), .B(KEYINPUT13), .C1(new_n353), .C2(new_n355), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n365), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n364), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n232), .A2(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n305), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n373), .A2(KEYINPUT12), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(KEYINPUT12), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n374), .A2(new_n375), .B1(new_n337), .B2(new_n216), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n372), .B1(G50), .B2(new_n291), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n223), .B2(new_n295), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n303), .A2(new_n378), .ZN(new_n379));
  XOR2_X1   g0179(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n303), .A2(new_n378), .A3(new_n380), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n376), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT76), .B(new_n376), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n371), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G190), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n366), .B2(new_n368), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n388), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n316), .B1(new_n356), .B2(new_n360), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n392), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n347), .A2(new_n389), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n293), .A2(new_n309), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT77), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n302), .A2(new_n306), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n399), .A2(new_n400), .B1(new_n306), .B2(new_n293), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NOR4_X1   g0203(.A1(new_n268), .A2(new_n269), .A3(new_n403), .A4(G20), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n270), .A2(new_n276), .A3(new_n232), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n403), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n216), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n226), .A2(new_n216), .ZN(new_n408));
  OAI21_X1  g0208(.A(G20), .B1(new_n408), .B2(new_n234), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n291), .A2(G159), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n407), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n273), .A2(new_n275), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n403), .B1(new_n413), .B2(G20), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n268), .A2(new_n269), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n411), .B1(new_n417), .B2(G68), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n336), .B1(new_n418), .B2(KEYINPUT16), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n401), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(KEYINPUT80), .A2(KEYINPUT17), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n280), .A2(new_n278), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n222), .A2(G1698), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n423), .C1(new_n268), .C2(new_n269), .ZN(new_n424));
  NAND2_X1  g0224(.A1(G33), .A2(G87), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(KEYINPUT78), .A3(new_n425), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n287), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n259), .B1(new_n265), .B2(G232), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n430), .A2(G190), .A3(new_n431), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n420), .A2(new_n421), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT80), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n435), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n430), .A2(new_n365), .A3(new_n431), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT79), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n432), .A2(new_n333), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT79), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n430), .A2(new_n443), .A3(new_n365), .A4(new_n431), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n412), .A2(new_n419), .ZN(new_n446));
  INV_X1    g0246(.A(new_n401), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(new_n420), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n332), .A2(G200), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n454), .B(new_n345), .C1(new_n390), .C2(new_n332), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n267), .A2(new_n288), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n333), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n267), .A2(new_n365), .A3(new_n288), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n312), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n439), .A2(new_n453), .A3(new_n455), .A4(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n397), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n306), .A2(G97), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n256), .A2(G33), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n302), .A2(new_n306), .A3(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n210), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n291), .A2(G77), .ZN(new_n467));
  NOR2_X1   g0267(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n210), .A2(new_n249), .ZN(new_n469));
  NOR2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(G97), .B(G107), .ZN(new_n472));
  NAND2_X1  g0272(.A1(KEYINPUT6), .A2(G107), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G20), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n467), .B(new_n476), .C1(new_n406), .C2(new_n328), .ZN(new_n477));
  AOI211_X1 g0277(.A(new_n463), .B(new_n466), .C1(new_n477), .C2(new_n298), .ZN(new_n478));
  NAND2_X1  g0278(.A1(G33), .A2(G283), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n224), .B1(new_n273), .B2(new_n275), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(KEYINPUT4), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n482), .A2(G1698), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n224), .B1(new_n270), .B2(new_n276), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n209), .B1(new_n270), .B2(new_n276), .ZN(new_n486));
  OAI21_X1  g0286(.A(G1698), .B1(new_n486), .B2(new_n482), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n331), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G45), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT5), .B(G41), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n261), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G257), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(G274), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n488), .A2(G190), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n277), .A2(G250), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n278), .B1(new_n497), .B2(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n277), .A2(G244), .A3(new_n483), .ZN(new_n499));
  INV_X1    g0299(.A(new_n479), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n413), .A2(G244), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n501), .B2(new_n482), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n287), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n495), .ZN(new_n505));
  AOI21_X1  g0305(.A(G200), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n478), .B1(new_n496), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n217), .A2(new_n278), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n224), .A2(G1698), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n509), .C1(new_n268), .C2(new_n269), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G116), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n287), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n256), .A2(G45), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(G250), .C1(new_n260), .C2(new_n231), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT82), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n284), .A2(new_n285), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n518), .A2(KEYINPUT82), .A3(G250), .A4(new_n514), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n490), .A2(G274), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n513), .A2(new_n520), .A3(G190), .A4(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT83), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n287), .A2(new_n512), .B1(G274), .B2(new_n490), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n524), .A2(new_n525), .A3(G190), .A4(new_n520), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n413), .A2(new_n232), .A3(G68), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n295), .A2(new_n210), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(KEYINPUT19), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G87), .A2(G97), .ZN(new_n533));
  NAND3_X1  g0333(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n328), .A2(new_n533), .B1(new_n232), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n298), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n343), .A2(new_n307), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n302), .A2(G87), .A3(new_n306), .A4(new_n464), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n316), .B1(new_n524), .B2(new_n520), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n526), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n529), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n477), .A2(new_n298), .ZN(new_n544));
  INV_X1    g0344(.A(new_n463), .ZN(new_n545));
  INV_X1    g0345(.A(new_n466), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n504), .A2(new_n365), .A3(new_n505), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n333), .B1(new_n488), .B2(new_n495), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n524), .A2(new_n520), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n365), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n551), .A2(new_n333), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n536), .B(new_n537), .C1(new_n343), .C2(new_n465), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AND4_X1   g0356(.A1(new_n507), .A2(new_n543), .A3(new_n550), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n211), .A2(G1698), .ZN(new_n558));
  OAI221_X1 g0358(.A(new_n558), .B1(G250), .B2(G1698), .C1(new_n268), .C2(new_n269), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G33), .A2(G294), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n287), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n492), .A2(G264), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n494), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G169), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n365), .B2(new_n564), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n232), .A2(G33), .A3(G116), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(new_n249), .A3(G20), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n232), .A2(KEYINPUT22), .A3(G87), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n568), .B(new_n570), .C1(new_n415), .C2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n569), .B1(new_n328), .B2(G20), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n208), .A2(G20), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n277), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n567), .B(new_n574), .C1(new_n576), .C2(KEYINPUT22), .ZN(new_n577));
  AOI21_X1  g0377(.A(KEYINPUT22), .B1(new_n277), .B2(new_n575), .ZN(new_n578));
  AND2_X1   g0378(.A1(KEYINPUT71), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(KEYINPUT71), .A2(G107), .ZN(new_n580));
  OAI21_X1  g0380(.A(G20), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT23), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n575), .B(KEYINPUT22), .C1(new_n269), .C2(new_n268), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n568), .A4(new_n570), .ZN(new_n584));
  OAI21_X1  g0384(.A(KEYINPUT86), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n577), .A2(new_n585), .A3(KEYINPUT24), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  OAI211_X1 g0387(.A(KEYINPUT86), .B(new_n587), .C1(new_n578), .C2(new_n584), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n298), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n307), .B2(new_n249), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n307), .A2(new_n249), .A3(new_n590), .ZN(new_n592));
  NOR2_X1   g0392(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n465), .ZN(new_n595));
  AOI211_X1 g0395(.A(new_n591), .B(new_n594), .C1(G107), .C2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n589), .A2(KEYINPUT88), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT88), .B1(new_n589), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n566), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n562), .A2(new_n390), .A3(new_n563), .A4(new_n494), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT89), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n564), .A2(new_n316), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n561), .A2(new_n287), .B1(new_n492), .B2(G264), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT89), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n390), .A4(new_n494), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n589), .A2(new_n596), .A3(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT90), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n589), .A2(KEYINPUT90), .A3(new_n596), .A4(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g0411(.A1(KEYINPUT5), .A2(G41), .ZN(new_n612));
  NOR2_X1   g0412(.A1(KEYINPUT5), .A2(G41), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n490), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(G270), .A3(new_n518), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n494), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT85), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT85), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n615), .A2(new_n618), .A3(new_n494), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n270), .A2(new_n276), .A3(G303), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n211), .A2(new_n278), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n413), .B(new_n621), .C1(G264), .C2(new_n278), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n617), .A2(new_n619), .B1(new_n287), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(G190), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n305), .A2(G20), .A3(new_n213), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n336), .A2(new_n306), .A3(G116), .A4(new_n464), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n479), .B(new_n232), .C1(G33), .C2(new_n210), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n628), .B(new_n298), .C1(new_n232), .C2(G116), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT20), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n626), .B(new_n627), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n625), .B(new_n634), .C1(new_n624), .C2(new_n316), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n623), .A2(new_n287), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n615), .A2(new_n618), .A3(new_n494), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n618), .B1(new_n615), .B2(new_n494), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n639), .A2(G169), .A3(new_n633), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n639), .A2(new_n633), .A3(KEYINPUT21), .A4(G169), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n636), .B(G179), .C1(new_n637), .C2(new_n638), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n633), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n635), .A2(new_n642), .A3(new_n643), .A4(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n557), .A2(new_n599), .A3(new_n611), .A4(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n462), .A2(new_n649), .ZN(G372));
  NAND2_X1  g0450(.A1(new_n589), .A2(new_n596), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n566), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n642), .A2(new_n643), .A3(new_n646), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n507), .A2(new_n550), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n541), .A2(new_n527), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n611), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n556), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n659));
  XOR2_X1   g0459(.A(KEYINPUT91), .B(KEYINPUT26), .Z(new_n660));
  NAND4_X1  g0460(.A1(new_n659), .A2(new_n556), .A3(new_n543), .A4(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n656), .A2(new_n556), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n550), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n461), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n459), .ZN(new_n668));
  INV_X1    g0468(.A(new_n389), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n396), .B1(new_n669), .B2(new_n346), .ZN(new_n670));
  INV_X1    g0470(.A(new_n439), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n453), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n322), .A2(KEYINPUT92), .A3(new_n323), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT92), .B1(new_n322), .B2(new_n323), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n668), .B1(new_n672), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n667), .A2(new_n676), .ZN(G369));
  INV_X1    g0477(.A(new_n305), .ZN(new_n678));
  OR3_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .A3(G20), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT27), .B1(new_n678), .B2(G20), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n597), .B2(new_n598), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n599), .A2(new_n684), .A3(new_n611), .ZN(new_n685));
  INV_X1    g0485(.A(new_n683), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n685), .B1(new_n599), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n642), .A2(new_n646), .A3(new_n643), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n634), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n647), .B2(new_n689), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G330), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n653), .A2(new_n683), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n599), .A2(new_n611), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n683), .B(KEYINPUT93), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n651), .A2(new_n566), .A3(new_n700), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n696), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n205), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n328), .A2(new_n213), .A3(new_n533), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n236), .B2(new_n706), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NOR3_X1   g0511(.A1(new_n644), .A2(new_n488), .A3(new_n495), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n552), .A2(new_n603), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n504), .A2(new_n624), .A3(G179), .A4(new_n505), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT30), .B1(new_n717), .B2(new_n714), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n564), .B(new_n551), .C1(new_n488), .C2(new_n495), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G179), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n716), .A2(new_n718), .B1(new_n720), .B2(new_n639), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n722), .A2(KEYINPUT31), .A3(new_n699), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n721), .B2(new_n686), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n723), .B(new_n725), .C1(new_n649), .C2(new_n699), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G330), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  INV_X1    g0529(.A(new_n663), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT26), .A3(new_n659), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n659), .A2(new_n556), .A3(new_n543), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(new_n660), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n611), .A2(new_n655), .A3(new_n656), .ZN(new_n734));
  INV_X1    g0534(.A(new_n598), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n589), .A2(KEYINPUT88), .A3(new_n596), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n688), .B1(new_n737), .B2(new_n566), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n733), .B(new_n556), .C1(new_n734), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n729), .B1(new_n739), .B2(new_n686), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n666), .A2(new_n700), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(KEYINPUT29), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n728), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n711), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n304), .A2(G20), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G45), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n706), .A2(G1), .A3(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n232), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT98), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n747), .B1(new_n692), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(G20), .B1(KEYINPUT94), .B2(G169), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(KEYINPUT94), .A2(G169), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n231), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n390), .A2(G20), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT96), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(G179), .A3(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G159), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT32), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n232), .A2(new_n365), .A3(G190), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G200), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G68), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n232), .A2(new_n365), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G190), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n232), .B1(new_n769), .B2(G190), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n768), .A2(G50), .B1(new_n771), .B2(G97), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n761), .A2(new_n277), .A3(new_n765), .A4(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n758), .A2(G179), .A3(new_n316), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G107), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT95), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n762), .A2(new_n776), .A3(new_n316), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n776), .B1(new_n762), .B2(new_n316), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n775), .B1(new_n779), .B2(new_n223), .C1(new_n760), .C2(KEYINPUT32), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n316), .A2(G179), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(G20), .A3(G190), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n208), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n766), .A2(G190), .A3(new_n316), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n226), .ZN(new_n785));
  NOR4_X1   g0585(.A1(new_n773), .A2(new_n780), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n277), .B1(new_n759), .B2(G329), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  INV_X1    g0588(.A(G303), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n782), .B(KEYINPUT97), .Z(new_n790));
  OAI221_X1 g0590(.A(new_n787), .B1(new_n788), .B2(new_n779), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G317), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n792), .A2(KEYINPUT33), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n764), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G326), .ZN(new_n796));
  INV_X1    g0596(.A(new_n774), .ZN(new_n797));
  INV_X1    g0597(.A(G283), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n795), .B1(new_n796), .B2(new_n767), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n784), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(G322), .ZN(new_n801));
  INV_X1    g0601(.A(G294), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n770), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g0603(.A1(new_n791), .A2(new_n799), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n755), .B1(new_n786), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n254), .A2(G45), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n704), .A2(new_n413), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G45), .C2(new_n236), .ZN(new_n808));
  INV_X1    g0608(.A(G355), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n277), .A2(new_n205), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n808), .B1(G116), .B2(new_n205), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n749), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n755), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n751), .A2(new_n805), .A3(new_n814), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n815), .B(KEYINPUT99), .Z(new_n816));
  INV_X1    g0616(.A(new_n747), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n694), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G330), .B2(new_n691), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n816), .A2(new_n819), .ZN(G396));
  OAI21_X1  g0620(.A(new_n455), .B1(new_n345), .B2(new_n686), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n334), .A2(new_n335), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n345), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n346), .A2(new_n686), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n741), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n666), .A2(new_n700), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n829), .B(new_n728), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n747), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n825), .A2(new_n748), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n755), .A2(new_n748), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n223), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n784), .A2(new_n802), .B1(new_n770), .B2(new_n210), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n779), .A2(new_n213), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n763), .A2(KEYINPUT100), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n763), .A2(KEYINPUT100), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n835), .B(new_n836), .C1(G283), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n774), .A2(G87), .ZN(new_n842));
  INV_X1    g0642(.A(new_n790), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n843), .A2(G107), .B1(new_n759), .B2(G311), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n277), .B1(new_n768), .B2(G303), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n841), .A2(new_n842), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n764), .A2(G150), .B1(new_n800), .B2(G143), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  INV_X1    g0648(.A(G159), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(new_n848), .B2(new_n767), .C1(new_n779), .C2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT34), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n797), .A2(new_n216), .B1(new_n790), .B2(new_n221), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G58), .B2(new_n771), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n413), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n759), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n846), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(new_n755), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n832), .A2(new_n817), .A3(new_n834), .A4(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n831), .A2(new_n860), .ZN(G384));
  NOR3_X1   g0661(.A1(new_n391), .A2(new_n388), .A3(new_n394), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n388), .B(new_n683), .C1(new_n371), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n388), .A2(new_n683), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n369), .A2(new_n362), .A3(new_n363), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n396), .B(new_n864), .C1(new_n865), .C2(new_n393), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  OR2_X1    g0667(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n418), .A2(KEYINPUT16), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n303), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n447), .ZN(new_n871));
  INV_X1    g0671(.A(new_n681), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n445), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n420), .A2(new_n433), .A3(new_n434), .ZN(new_n874));
  AND3_X1   g0674(.A1(new_n873), .A2(KEYINPUT37), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n446), .A2(new_n447), .A3(new_n434), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n876), .A2(new_n421), .A3(new_n433), .A4(new_n438), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n436), .A3(new_n437), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n453), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n681), .B1(new_n870), .B2(new_n447), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  INV_X1    g0682(.A(new_n874), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n420), .B1(new_n451), .B2(new_n681), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n881), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT101), .ZN(new_n891));
  INV_X1    g0691(.A(new_n824), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n699), .B1(new_n657), .B2(new_n665), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n891), .B(new_n892), .C1(new_n893), .C2(new_n827), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT101), .B1(new_n828), .B2(new_n824), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n867), .B(new_n890), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n449), .A2(new_n452), .A3(new_n681), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT102), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n448), .A2(new_n872), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n439), .B2(new_n453), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n882), .B1(new_n901), .B2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g0703(.A(new_n884), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n903), .A2(new_n904), .A3(new_n874), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n420), .A2(new_n681), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT103), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT37), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n883), .B2(new_n884), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n887), .B1(new_n902), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n889), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT39), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n890), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n389), .A2(new_n683), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n896), .A2(KEYINPUT102), .A3(new_n897), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n900), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n461), .B1(new_n740), .B2(new_n742), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n676), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n920), .B(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n911), .A2(new_n889), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n507), .A2(new_n543), .A3(new_n550), .A4(new_n556), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n925), .A2(new_n647), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n926), .A2(new_n599), .A3(new_n611), .A4(new_n700), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT104), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n716), .A2(new_n718), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n720), .A2(new_n639), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n686), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n928), .B1(new_n931), .B2(KEYINPUT31), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n721), .A2(KEYINPUT104), .A3(new_n724), .A4(new_n686), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n927), .B(new_n725), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n825), .B1(new_n863), .B2(new_n866), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT40), .B1(new_n924), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n867), .A2(new_n827), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n927), .A2(new_n725), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n932), .A2(new_n933), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n890), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n937), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n461), .A2(new_n934), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n946), .A2(new_n693), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n923), .B(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n256), .B2(new_n745), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n213), .B1(new_n475), .B2(KEYINPUT35), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n233), .C1(KEYINPUT35), .C2(new_n475), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI21_X1  g0752(.A(G77), .B1(new_n226), .B2(new_n216), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n236), .A2(new_n953), .B1(G50), .B2(new_n216), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n304), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n949), .A2(new_n952), .A3(new_n955), .ZN(G367));
  INV_X1    g0756(.A(KEYINPUT108), .ZN(new_n957));
  INV_X1    g0757(.A(new_n807), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n813), .B1(new_n205), .B2(new_n343), .C1(new_n246), .C2(new_n958), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n840), .A2(G159), .B1(G143), .B2(new_n768), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n216), .B2(new_n770), .ZN(new_n961));
  INV_X1    g0761(.A(new_n277), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n797), .A2(new_n223), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n782), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G150), .A2(new_n800), .B1(new_n965), .B2(G58), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n966), .C1(new_n848), .C2(new_n855), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n779), .A2(new_n221), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n797), .A2(new_n210), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n415), .B1(new_n779), .B2(new_n798), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G317), .B2(new_n759), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n771), .A2(new_n329), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n782), .B2(new_n213), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n789), .B2(new_n784), .C1(new_n788), .C2(new_n767), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n840), .B2(G294), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n843), .A2(KEYINPUT46), .A3(G116), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n971), .A2(new_n972), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n967), .A2(new_n968), .B1(new_n969), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n755), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n959), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n539), .A2(new_n683), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n730), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n556), .B2(new_n984), .ZN(new_n986));
  INV_X1    g0786(.A(new_n750), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n983), .A2(new_n747), .A3(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT107), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n746), .A2(G1), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT45), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n547), .A2(new_n699), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n507), .A2(new_n550), .A3(new_n993), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n547), .A2(new_n699), .A3(new_n548), .A4(new_n549), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT105), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n996), .B1(new_n994), .B2(new_n995), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n698), .A2(new_n701), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n994), .A2(new_n995), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(KEYINPUT105), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n994), .A2(new_n996), .A3(new_n995), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1005), .A2(KEYINPUT45), .A3(new_n701), .A4(new_n698), .ZN(new_n1006));
  AND2_X1   g0806(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT44), .B1(new_n702), .B2(new_n1005), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n999), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n695), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n698), .B1(new_n687), .B2(new_n697), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n694), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n999), .A2(new_n1000), .A3(new_n1009), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1009), .B1(new_n999), .B2(new_n1000), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1017), .A2(new_n696), .A3(new_n1018), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1012), .A2(new_n743), .A3(new_n1014), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n743), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n705), .B(KEYINPUT41), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n991), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n599), .A2(new_n684), .A3(new_n611), .A4(new_n697), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT42), .B1(new_n999), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1024), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT42), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1026), .A2(new_n1005), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n599), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n659), .B1(new_n1005), .B2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1025), .B(new_n1028), .C1(new_n1030), .C2(new_n699), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1033), .A2(new_n695), .A3(new_n1005), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n695), .A2(new_n1005), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1031), .A2(new_n1036), .A3(new_n1032), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1035), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1037), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1036), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n957), .B(new_n990), .C1(new_n1023), .C2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1022), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n1020), .B2(new_n743), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1038), .B(new_n1042), .C1(new_n1047), .C2(new_n991), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n957), .B1(new_n1048), .B2(new_n990), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G387));
  OR2_X1    g0851(.A1(new_n743), .A2(new_n1014), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n743), .A2(new_n1014), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n705), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1014), .A2(new_n991), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n779), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1056), .A2(G303), .B1(G317), .B2(new_n800), .ZN(new_n1057));
  XOR2_X1   g0857(.A(KEYINPUT110), .B(G322), .Z(new_n1058));
  NAND2_X1  g0858(.A1(new_n768), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1057), .B(new_n1059), .C1(new_n788), .C2(new_n839), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT48), .Z(new_n1061));
  NOR2_X1   g0861(.A1(new_n770), .A2(new_n798), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n782), .A2(new_n802), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1064), .A2(KEYINPUT49), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n415), .B1(new_n855), .B2(new_n796), .C1(new_n213), .C2(new_n797), .ZN(new_n1067));
  OR3_X1    g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n969), .B1(G150), .B2(new_n759), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1056), .A2(G68), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n343), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n771), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n294), .A2(new_n763), .B1(new_n221), .B2(new_n784), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n767), .A2(new_n849), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n782), .A2(new_n223), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n415), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .A4(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n982), .B1(new_n1068), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n243), .A2(G45), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n293), .A2(new_n221), .ZN(new_n1080));
  XOR2_X1   g0880(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n1081));
  XNOR2_X1  g0881(.A(new_n1080), .B(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n708), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1079), .A2(new_n807), .A3(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(G107), .B2(new_n205), .C1(new_n708), .C2(new_n810), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1086), .A2(new_n813), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1078), .A2(new_n747), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n687), .B2(new_n987), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1054), .A2(new_n1055), .A3(new_n1089), .ZN(G393));
  NAND2_X1  g0890(.A1(new_n1012), .A2(new_n1019), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n706), .B1(new_n1091), .B2(new_n1053), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1020), .ZN(new_n1093));
  AND4_X1   g0893(.A1(new_n696), .A2(new_n1018), .A3(new_n1008), .A4(new_n1010), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n696), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1095));
  OAI21_X1  g0895(.A(KEYINPUT111), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT111), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1012), .A2(new_n1097), .A3(new_n1019), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n991), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n747), .B1(new_n999), .B2(new_n812), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n251), .A2(new_n807), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1101), .B(new_n813), .C1(new_n210), .C2(new_n205), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n415), .B1(new_n759), .B2(G143), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n842), .C1(new_n216), .C2(new_n782), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n768), .B1(new_n800), .B2(G159), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(KEYINPUT51), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n293), .B2(new_n1056), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n221), .B2(new_n839), .C1(new_n223), .C2(new_n770), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1104), .B(new_n1108), .C1(KEYINPUT51), .C2(new_n1105), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1056), .A2(G294), .B1(new_n774), .B2(G107), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n962), .B1(new_n798), .B2(new_n782), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n759), .B2(new_n1058), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n771), .A2(G116), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n784), .A2(new_n788), .B1(new_n767), .B2(new_n792), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT52), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .A4(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(G303), .B2(new_n840), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n755), .B1(new_n1109), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1100), .A2(new_n1102), .A3(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1099), .A2(KEYINPUT112), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT112), .B1(new_n1099), .B2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1093), .B1(new_n1120), .B2(new_n1121), .ZN(G390));
  INV_X1    g0922(.A(new_n867), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n895), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n828), .A2(KEYINPUT101), .A3(new_n824), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n915), .B1(new_n1126), .B2(new_n916), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n739), .A2(new_n686), .A3(new_n823), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1128), .A2(new_n824), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n912), .B(new_n917), .C1(new_n1129), .C2(new_n1123), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n934), .A2(G330), .A3(new_n935), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n727), .A2(new_n938), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1127), .A2(new_n1130), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n991), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n915), .A2(new_n748), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n833), .A2(new_n294), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n768), .A2(G283), .B1(new_n771), .B2(G77), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1140), .B1(new_n839), .B2(new_n328), .C1(new_n802), .C2(new_n855), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n962), .B1(new_n790), .B2(new_n208), .C1(new_n797), .C2(new_n216), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n784), .A2(new_n213), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n779), .A2(new_n210), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n768), .A2(G128), .B1(new_n771), .B2(G159), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT116), .Z(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1146), .B1(new_n839), .B2(new_n848), .C1(new_n779), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n759), .A2(G125), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1151), .B(new_n277), .C1(new_n797), .C2(new_n221), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n784), .A2(new_n856), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n965), .A2(G150), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT53), .ZN(new_n1155));
  NOR4_X1   g0955(.A1(new_n1150), .A2(new_n1152), .A3(new_n1153), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n755), .B1(new_n1145), .B2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1138), .A2(new_n817), .A3(new_n1139), .A4(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1137), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT117), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT115), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n934), .A2(G330), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(KEYINPUT114), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT114), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n934), .A2(new_n1165), .A3(G330), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1164), .A2(new_n827), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1134), .B1(new_n1167), .B2(new_n1123), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n726), .A2(G330), .A3(new_n827), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1123), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT113), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(KEYINPUT113), .A3(new_n1123), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(new_n1132), .A3(new_n1174), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1168), .A2(new_n1129), .B1(new_n1169), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n461), .A2(G330), .A3(new_n934), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n921), .A2(new_n1177), .A3(new_n676), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1162), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1134), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n934), .A2(new_n1165), .A3(G330), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1165), .B1(new_n934), .B2(G330), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n825), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1129), .B(new_n1180), .C1(new_n1183), .C2(new_n867), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1175), .A2(new_n1169), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1178), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(KEYINPUT115), .A3(new_n1187), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1179), .A2(new_n1133), .A3(new_n1188), .A4(new_n1135), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT115), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1162), .B(new_n1178), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1136), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1189), .A2(new_n1192), .A3(new_n705), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n1158), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1161), .A2(new_n1193), .A3(new_n1194), .ZN(G378));
  AND3_X1   g0995(.A1(new_n896), .A2(KEYINPUT102), .A3(new_n897), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT102), .B1(new_n896), .B2(new_n897), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n312), .A2(new_n872), .ZN(new_n1199));
  XOR2_X1   g0999(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(new_n675), .B2(new_n459), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n673), .A2(new_n674), .A3(new_n668), .A4(new_n1201), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n944), .A2(G330), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n942), .B1(new_n941), .B2(new_n912), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n879), .A2(new_n880), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n875), .ZN(new_n1210));
  AND4_X1   g1010(.A1(KEYINPUT38), .A2(new_n1209), .A3(new_n885), .A4(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT38), .B1(new_n881), .B2(new_n885), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n934), .A2(new_n942), .A3(new_n935), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(G330), .B1(new_n1208), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(new_n1205), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1198), .A2(new_n918), .A3(new_n1207), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1217), .A2(new_n1207), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n920), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1220), .A3(KEYINPUT57), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1192), .B2(new_n1187), .ZN(new_n1222));
  OAI21_X1  g1022(.A(KEYINPUT119), .B1(new_n1222), .B2(new_n706), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT57), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1179), .A2(new_n1188), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1178), .B1(new_n1225), .B2(new_n1136), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT119), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n705), .C1(new_n1226), .C2(new_n1221), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1223), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1227), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n991), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1206), .A2(new_n748), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n221), .B1(new_n268), .B2(G41), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n763), .A2(new_n856), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n768), .A2(G125), .B1(new_n771), .B2(G150), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT118), .Z(new_n1238));
  AOI211_X1 g1038(.A(new_n1236), .B(new_n1238), .C1(G128), .C2(new_n800), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n848), .B2(new_n779), .C1(new_n782), .C2(new_n1149), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n774), .A2(G159), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G41), .B1(new_n759), .B2(G124), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1241), .A2(new_n272), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1240), .A2(KEYINPUT59), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1235), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(G41), .B1(new_n1056), .B2(new_n1071), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n800), .A2(G107), .B1(new_n771), .B2(G68), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1247), .B(new_n1248), .C1(new_n226), .C2(new_n797), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n1075), .B(new_n1249), .C1(G283), .C2(new_n759), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n413), .B1(new_n764), .B2(G97), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n213), .C2(new_n767), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT58), .Z(new_n1253));
  OAI21_X1  g1053(.A(new_n755), .B1(new_n1246), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n833), .A2(new_n221), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1234), .A2(new_n817), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1233), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1231), .A2(new_n1258), .ZN(G375));
  AOI21_X1  g1059(.A(new_n415), .B1(new_n774), .B2(G58), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT121), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1056), .A2(G150), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n839), .C2(new_n1149), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G137), .B2(new_n800), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n771), .A2(G50), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n759), .A2(G128), .B1(G132), .B2(new_n768), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G159), .B2(new_n843), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n843), .A2(G97), .B1(new_n759), .B2(G303), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(new_n1269), .B(KEYINPUT120), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n840), .A2(G116), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1056), .A2(new_n329), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1270), .A2(new_n1072), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n962), .B1(new_n802), .B2(new_n767), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n784), .A2(new_n798), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1273), .A2(new_n963), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n755), .B1(new_n1268), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1123), .A2(new_n748), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1278), .A3(new_n817), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1279), .B1(new_n216), .B2(new_n833), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1186), .B2(new_n991), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1179), .A2(new_n1188), .A3(new_n1282), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1281), .B1(new_n1283), .B2(new_n1046), .ZN(G381));
  NOR3_X1   g1084(.A1(G381), .A2(G396), .A3(G393), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1099), .A2(new_n1119), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT112), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1099), .A2(KEYINPUT112), .A3(new_n1119), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n1289), .A2(new_n1290), .B1(new_n1020), .B2(new_n1092), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1285), .A2(new_n1286), .A3(new_n1050), .A4(new_n1291), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1292), .A2(KEYINPUT122), .ZN(new_n1293));
  INV_X1    g1093(.A(G378), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1231), .A2(new_n1294), .A3(new_n1258), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(KEYINPUT122), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1295), .A3(new_n1296), .ZN(G407));
  NAND3_X1  g1097(.A1(new_n1231), .A2(new_n1294), .A3(new_n1258), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G407), .B(G213), .C1(G343), .C2(new_n1298), .ZN(G409));
  NAND2_X1  g1099(.A1(G375), .A2(G378), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n682), .A2(G213), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1192), .A2(new_n1187), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1022), .A3(new_n1232), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT123), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT123), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1302), .A2(new_n1305), .A3(new_n1022), .A4(new_n1232), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1294), .A3(new_n1258), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1300), .A2(new_n1301), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT60), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1283), .B2(KEYINPUT60), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n705), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1281), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1286), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1312), .A2(G384), .A3(new_n1281), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1301), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(G2897), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1314), .A2(new_n1315), .A3(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1317), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1320), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1300), .A2(new_n1301), .A3(new_n1308), .A4(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1294), .B1(new_n1231), .B2(new_n1258), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(new_n1316), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT62), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1326), .A2(new_n1327), .A3(new_n1308), .A4(new_n1322), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1321), .A2(new_n1324), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1330), .A2(new_n1048), .A3(new_n990), .A4(new_n1093), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n990), .B1(new_n1023), .B2(new_n1043), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(G390), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(G396), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(G393), .B(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1331), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1336));
  AOI22_X1  g1136(.A1(new_n1330), .A2(new_n1093), .B1(new_n1048), .B2(new_n990), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1337), .B1(new_n1050), .B2(new_n1291), .ZN(new_n1338));
  OAI211_X1 g1138(.A(KEYINPUT126), .B(new_n1336), .C1(new_n1338), .C2(new_n1335), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT126), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1332), .A2(KEYINPUT108), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1291), .A2(new_n1341), .A3(new_n1044), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1335), .B1(new_n1342), .B2(new_n1333), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1331), .A2(new_n1333), .A3(new_n1335), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1340), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1339), .A2(new_n1345), .ZN(new_n1346));
  AND3_X1   g1146(.A1(new_n1300), .A2(new_n1301), .A3(new_n1308), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT125), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1347), .A2(new_n1348), .A3(KEYINPUT63), .A4(new_n1322), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT63), .ZN(new_n1350));
  OAI21_X1  g1150(.A(KEYINPUT125), .B1(new_n1323), .B2(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1336), .B1(new_n1338), .B2(new_n1335), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1323), .A2(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1321), .A2(new_n1353), .A3(new_n1355), .ZN(new_n1356));
  OAI22_X1  g1156(.A1(new_n1329), .A2(new_n1346), .B1(new_n1352), .B2(new_n1356), .ZN(G405));
  OAI21_X1  g1157(.A(new_n1346), .B1(new_n1295), .B2(new_n1325), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT127), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1339), .A2(new_n1345), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1300), .A2(new_n1298), .A3(new_n1360), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1358), .A2(new_n1359), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1359), .B1(new_n1358), .B2(new_n1361), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1322), .ZN(new_n1364));
  NOR3_X1   g1164(.A1(new_n1362), .A2(new_n1363), .A3(new_n1364), .ZN(new_n1365));
  AND3_X1   g1165(.A1(new_n1300), .A2(new_n1298), .A3(new_n1360), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1360), .B1(new_n1300), .B2(new_n1298), .ZN(new_n1367));
  OAI21_X1  g1167(.A(KEYINPUT127), .B1(new_n1366), .B2(new_n1367), .ZN(new_n1368));
  NAND3_X1  g1168(.A1(new_n1358), .A2(new_n1361), .A3(new_n1359), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1322), .B1(new_n1368), .B2(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1365), .A2(new_n1370), .ZN(G402));
endmodule


