

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U554 ( .A1(n725), .A2(n724), .ZN(n730) );
  NAND2_X1 U555 ( .A1(n616), .A2(n615), .ZN(n986) );
  AND2_X1 U556 ( .A1(n813), .A2(n707), .ZN(n709) );
  XNOR2_X1 U557 ( .A(n555), .B(KEYINPUT23), .ZN(n556) );
  XNOR2_X1 U558 ( .A(n539), .B(n538), .ZN(n585) );
  AND2_X2 U559 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U560 ( .A(n737), .B(KEYINPUT94), .ZN(n741) );
  INV_X1 U561 ( .A(n755), .ZN(n732) );
  NOR2_X1 U562 ( .A1(G1966), .A2(n810), .ZN(n776) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n606) );
  NOR2_X2 U564 ( .A1(n719), .A2(n986), .ZN(n720) );
  XNOR2_X2 U565 ( .A(n525), .B(KEYINPUT0), .ZN(n655) );
  OR2_X1 U566 ( .A1(n542), .A2(KEYINPUT67), .ZN(n543) );
  BUF_X1 U567 ( .A(n617), .Z(n532) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n531), .Z(n617) );
  NOR2_X2 U569 ( .A1(n655), .A2(G651), .ZN(n676) );
  NOR2_X1 U570 ( .A1(G543), .A2(n530), .ZN(n531) );
  NOR2_X2 U571 ( .A1(n557), .A2(n556), .ZN(n520) );
  NOR2_X1 U572 ( .A1(n557), .A2(n556), .ZN(n716) );
  AND2_X1 U573 ( .A1(n545), .A2(G2105), .ZN(n589) );
  NOR2_X2 U574 ( .A1(n741), .A2(n740), .ZN(n744) );
  AND2_X1 U575 ( .A1(n786), .A2(n785), .ZN(n787) );
  INV_X1 U576 ( .A(n1000), .ZN(n785) );
  NAND2_X1 U577 ( .A1(n770), .A2(n769), .ZN(n771) );
  OR2_X1 U578 ( .A1(n768), .A2(n767), .ZN(n769) );
  BUF_X1 U579 ( .A(n589), .Z(n916) );
  AND2_X1 U580 ( .A1(n551), .A2(G101), .ZN(n552) );
  NOR2_X1 U581 ( .A1(n723), .A2(n522), .ZN(n724) );
  XNOR2_X1 U582 ( .A(n742), .B(KEYINPUT29), .ZN(n743) );
  INV_X1 U583 ( .A(KEYINPUT95), .ZN(n742) );
  AND2_X1 U584 ( .A1(n781), .A2(n521), .ZN(n782) );
  XNOR2_X1 U585 ( .A(n771), .B(KEYINPUT32), .ZN(n783) );
  NAND2_X1 U586 ( .A1(G8), .A2(n755), .ZN(n810) );
  INV_X1 U587 ( .A(G2104), .ZN(n545) );
  INV_X1 U588 ( .A(KEYINPUT17), .ZN(n538) );
  NOR2_X2 U589 ( .A1(G2104), .A2(G2105), .ZN(n539) );
  INV_X1 U590 ( .A(KEYINPUT13), .ZN(n611) );
  INV_X1 U591 ( .A(KEYINPUT83), .ZN(n593) );
  NOR2_X1 U592 ( .A1(n623), .A2(n622), .ZN(n624) );
  BUF_X1 U593 ( .A(n606), .Z(n669) );
  NAND2_X1 U594 ( .A1(n547), .A2(n546), .ZN(n557) );
  BUF_X1 U595 ( .A(n520), .Z(G160) );
  BUF_X1 U596 ( .A(n585), .Z(n913) );
  NAND2_X1 U597 ( .A1(n548), .A2(G2104), .ZN(n549) );
  AND2_X1 U598 ( .A1(n780), .A2(n779), .ZN(n521) );
  AND2_X1 U599 ( .A1(n732), .A2(n1007), .ZN(n522) );
  XOR2_X1 U600 ( .A(KEYINPUT6), .B(n535), .Z(n523) );
  INV_X1 U601 ( .A(KEYINPUT93), .ZN(n727) );
  XNOR2_X1 U602 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U603 ( .A1(n755), .A2(G2084), .ZN(n756) );
  INV_X1 U604 ( .A(G168), .ZN(n759) );
  AND2_X1 U605 ( .A1(G8), .A2(n752), .ZN(n754) );
  INV_X1 U606 ( .A(KEYINPUT31), .ZN(n764) );
  INV_X1 U607 ( .A(n993), .ZN(n789) );
  NOR2_X1 U608 ( .A1(n810), .A2(n789), .ZN(n790) );
  NOR2_X1 U609 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U610 ( .A(n607), .B(KEYINPUT12), .ZN(n608) );
  INV_X1 U611 ( .A(G2105), .ZN(n548) );
  INV_X1 U612 ( .A(KEYINPUT101), .ZN(n847) );
  INV_X1 U613 ( .A(G543), .ZN(n525) );
  XNOR2_X1 U614 ( .A(KEYINPUT7), .B(n537), .ZN(G168) );
  NAND2_X1 U615 ( .A1(n669), .A2(G89), .ZN(n524) );
  XNOR2_X1 U616 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  INV_X1 U617 ( .A(G651), .ZN(n530) );
  NOR2_X2 U618 ( .A1(n655), .A2(n530), .ZN(n672) );
  NAND2_X1 U619 ( .A1(G76), .A2(n672), .ZN(n526) );
  NAND2_X1 U620 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U621 ( .A(KEYINPUT5), .B(n528), .ZN(n536) );
  NAND2_X1 U622 ( .A1(n676), .A2(G51), .ZN(n529) );
  XOR2_X1 U623 ( .A(KEYINPUT73), .B(n529), .Z(n534) );
  NAND2_X1 U624 ( .A1(n532), .A2(G63), .ZN(n533) );
  NAND2_X1 U625 ( .A1(n534), .A2(n533), .ZN(n535) );
  NAND2_X1 U626 ( .A1(n536), .A2(n523), .ZN(n537) );
  NAND2_X1 U627 ( .A1(n585), .A2(G137), .ZN(n541) );
  AND2_X4 U628 ( .A1(G2105), .A2(G2104), .ZN(n590) );
  NAND2_X1 U629 ( .A1(G113), .A2(n590), .ZN(n540) );
  NAND2_X1 U630 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n542), .A2(KEYINPUT67), .ZN(n544) );
  NAND2_X1 U632 ( .A1(n544), .A2(n543), .ZN(n547) );
  NAND2_X1 U633 ( .A1(G125), .A2(n916), .ZN(n546) );
  XNOR2_X2 U634 ( .A(n549), .B(KEYINPUT65), .ZN(n586) );
  NAND2_X1 U635 ( .A1(n586), .A2(G101), .ZN(n550) );
  NAND2_X1 U636 ( .A1(n550), .A2(KEYINPUT66), .ZN(n554) );
  INV_X1 U637 ( .A(KEYINPUT66), .ZN(n551) );
  NAND2_X1 U638 ( .A1(n586), .A2(n552), .ZN(n553) );
  NAND2_X1 U639 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U640 ( .A(G2435), .B(G2427), .Z(n559) );
  XNOR2_X1 U641 ( .A(G2446), .B(G2454), .ZN(n558) );
  XNOR2_X1 U642 ( .A(n559), .B(n558), .ZN(n565) );
  XOR2_X1 U643 ( .A(G2451), .B(G2430), .Z(n561) );
  XNOR2_X1 U644 ( .A(G1348), .B(G1341), .ZN(n560) );
  XNOR2_X1 U645 ( .A(n561), .B(n560), .ZN(n563) );
  XOR2_X1 U646 ( .A(G2438), .B(G2443), .Z(n562) );
  XNOR2_X1 U647 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U648 ( .A(n565), .B(n564), .Z(n566) );
  AND2_X1 U649 ( .A1(G14), .A2(n566), .ZN(G401) );
  NAND2_X1 U650 ( .A1(G52), .A2(n676), .ZN(n568) );
  NAND2_X1 U651 ( .A1(G64), .A2(n532), .ZN(n567) );
  NAND2_X1 U652 ( .A1(n568), .A2(n567), .ZN(n574) );
  NAND2_X1 U653 ( .A1(G77), .A2(n672), .ZN(n570) );
  NAND2_X1 U654 ( .A1(G90), .A2(n669), .ZN(n569) );
  NAND2_X1 U655 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U656 ( .A(KEYINPUT69), .B(n571), .ZN(n572) );
  XNOR2_X1 U657 ( .A(KEYINPUT9), .B(n572), .ZN(n573) );
  NOR2_X1 U658 ( .A1(n574), .A2(n573), .ZN(G171) );
  AND2_X1 U659 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U660 ( .A1(G123), .A2(n916), .ZN(n575) );
  XNOR2_X1 U661 ( .A(n575), .B(KEYINPUT18), .ZN(n583) );
  NAND2_X1 U662 ( .A1(G135), .A2(n913), .ZN(n578) );
  BUF_X1 U663 ( .A(n586), .Z(n576) );
  NAND2_X1 U664 ( .A1(G99), .A2(n576), .ZN(n577) );
  NAND2_X1 U665 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U666 ( .A1(n590), .A2(G111), .ZN(n579) );
  XOR2_X1 U667 ( .A(KEYINPUT74), .B(n579), .Z(n580) );
  NOR2_X1 U668 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n583), .A2(n582), .ZN(n954) );
  XNOR2_X1 U670 ( .A(G2096), .B(n954), .ZN(n584) );
  OR2_X1 U671 ( .A1(G2100), .A2(n584), .ZN(G156) );
  INV_X1 U672 ( .A(G57), .ZN(G237) );
  INV_X1 U673 ( .A(G132), .ZN(G219) );
  INV_X1 U674 ( .A(G82), .ZN(G220) );
  NAND2_X1 U675 ( .A1(G138), .A2(n585), .ZN(n588) );
  NAND2_X1 U676 ( .A1(G102), .A2(n586), .ZN(n587) );
  NAND2_X1 U677 ( .A1(n588), .A2(n587), .ZN(n596) );
  NAND2_X1 U678 ( .A1(G126), .A2(n589), .ZN(n592) );
  NAND2_X1 U679 ( .A1(G114), .A2(n590), .ZN(n591) );
  NAND2_X1 U680 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U681 ( .A(n594), .B(n593), .ZN(n595) );
  NOR2_X1 U682 ( .A1(n596), .A2(n595), .ZN(n706) );
  BUF_X1 U683 ( .A(n706), .Z(G164) );
  NAND2_X1 U684 ( .A1(G75), .A2(n672), .ZN(n598) );
  NAND2_X1 U685 ( .A1(G88), .A2(n669), .ZN(n597) );
  NAND2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U687 ( .A1(G50), .A2(n676), .ZN(n600) );
  NAND2_X1 U688 ( .A1(G62), .A2(n532), .ZN(n599) );
  NAND2_X1 U689 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U690 ( .A1(n602), .A2(n601), .ZN(G166) );
  XOR2_X1 U691 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U692 ( .A1(G7), .A2(G661), .ZN(n603) );
  XNOR2_X1 U693 ( .A(n603), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U694 ( .A(G223), .ZN(n867) );
  NAND2_X1 U695 ( .A1(n867), .A2(G567), .ZN(n604) );
  XOR2_X1 U696 ( .A(KEYINPUT11), .B(n604), .Z(G234) );
  NAND2_X1 U697 ( .A1(G56), .A2(n617), .ZN(n605) );
  XOR2_X1 U698 ( .A(KEYINPUT14), .B(n605), .Z(n614) );
  NAND2_X1 U699 ( .A1(G68), .A2(n672), .ZN(n610) );
  NAND2_X1 U700 ( .A1(G81), .A2(n606), .ZN(n607) );
  XNOR2_X1 U701 ( .A(n608), .B(KEYINPUT72), .ZN(n609) );
  NAND2_X1 U702 ( .A1(n610), .A2(n609), .ZN(n612) );
  XNOR2_X1 U703 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X2 U704 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U705 ( .A1(n676), .A2(G43), .ZN(n615) );
  INV_X1 U706 ( .A(G860), .ZN(n644) );
  OR2_X1 U707 ( .A1(n986), .A2(n644), .ZN(G153) );
  INV_X1 U708 ( .A(G171), .ZN(G301) );
  NAND2_X1 U709 ( .A1(G868), .A2(G301), .ZN(n626) );
  NAND2_X1 U710 ( .A1(G92), .A2(n669), .ZN(n619) );
  NAND2_X1 U711 ( .A1(G66), .A2(n617), .ZN(n618) );
  NAND2_X1 U712 ( .A1(n619), .A2(n618), .ZN(n623) );
  NAND2_X1 U713 ( .A1(G79), .A2(n672), .ZN(n621) );
  NAND2_X1 U714 ( .A1(G54), .A2(n676), .ZN(n620) );
  NAND2_X1 U715 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U716 ( .A(KEYINPUT15), .B(n624), .Z(n977) );
  OR2_X1 U717 ( .A1(n977), .A2(G868), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n626), .A2(n625), .ZN(G284) );
  NAND2_X1 U719 ( .A1(G78), .A2(n672), .ZN(n627) );
  XNOR2_X1 U720 ( .A(n627), .B(KEYINPUT70), .ZN(n634) );
  NAND2_X1 U721 ( .A1(G91), .A2(n669), .ZN(n629) );
  NAND2_X1 U722 ( .A1(G53), .A2(n676), .ZN(n628) );
  NAND2_X1 U723 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U724 ( .A1(G65), .A2(n532), .ZN(n630) );
  XNOR2_X1 U725 ( .A(KEYINPUT71), .B(n630), .ZN(n631) );
  NOR2_X1 U726 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U727 ( .A1(n634), .A2(n633), .ZN(G299) );
  INV_X1 U728 ( .A(G868), .ZN(n688) );
  NOR2_X1 U729 ( .A1(G286), .A2(n688), .ZN(n636) );
  NOR2_X1 U730 ( .A1(G868), .A2(G299), .ZN(n635) );
  NOR2_X1 U731 ( .A1(n636), .A2(n635), .ZN(G297) );
  NAND2_X1 U732 ( .A1(n644), .A2(G559), .ZN(n637) );
  NAND2_X1 U733 ( .A1(n637), .A2(n977), .ZN(n638) );
  XNOR2_X1 U734 ( .A(n638), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U735 ( .A1(G868), .A2(n986), .ZN(n641) );
  NAND2_X1 U736 ( .A1(G868), .A2(n977), .ZN(n639) );
  NOR2_X1 U737 ( .A1(G559), .A2(n639), .ZN(n640) );
  NOR2_X1 U738 ( .A1(n641), .A2(n640), .ZN(G282) );
  XNOR2_X1 U739 ( .A(n986), .B(KEYINPUT75), .ZN(n643) );
  NAND2_X1 U740 ( .A1(n977), .A2(G559), .ZN(n642) );
  XNOR2_X1 U741 ( .A(n643), .B(n642), .ZN(n685) );
  NAND2_X1 U742 ( .A1(n644), .A2(n685), .ZN(n654) );
  NAND2_X1 U743 ( .A1(G55), .A2(n676), .ZN(n646) );
  NAND2_X1 U744 ( .A1(G67), .A2(n532), .ZN(n645) );
  NAND2_X1 U745 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U746 ( .A(KEYINPUT78), .B(n647), .ZN(n653) );
  NAND2_X1 U747 ( .A1(n669), .A2(G93), .ZN(n648) );
  XNOR2_X1 U748 ( .A(n648), .B(KEYINPUT76), .ZN(n650) );
  NAND2_X1 U749 ( .A1(G80), .A2(n672), .ZN(n649) );
  NAND2_X1 U750 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U751 ( .A(KEYINPUT77), .B(n651), .Z(n652) );
  NOR2_X1 U752 ( .A1(n653), .A2(n652), .ZN(n687) );
  XOR2_X1 U753 ( .A(n654), .B(n687), .Z(G145) );
  NAND2_X1 U754 ( .A1(G49), .A2(n676), .ZN(n657) );
  NAND2_X1 U755 ( .A1(G87), .A2(n655), .ZN(n656) );
  NAND2_X1 U756 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U757 ( .A1(n532), .A2(n658), .ZN(n661) );
  NAND2_X1 U758 ( .A1(G74), .A2(G651), .ZN(n659) );
  XOR2_X1 U759 ( .A(KEYINPUT79), .B(n659), .Z(n660) );
  NAND2_X1 U760 ( .A1(n661), .A2(n660), .ZN(G288) );
  NAND2_X1 U761 ( .A1(G72), .A2(n672), .ZN(n663) );
  NAND2_X1 U762 ( .A1(G85), .A2(n669), .ZN(n662) );
  NAND2_X1 U763 ( .A1(n663), .A2(n662), .ZN(n666) );
  NAND2_X1 U764 ( .A1(G60), .A2(n532), .ZN(n664) );
  XOR2_X1 U765 ( .A(KEYINPUT68), .B(n664), .Z(n665) );
  NOR2_X1 U766 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U767 ( .A1(n676), .A2(G47), .ZN(n667) );
  NAND2_X1 U768 ( .A1(n668), .A2(n667), .ZN(G290) );
  NAND2_X1 U769 ( .A1(G86), .A2(n669), .ZN(n671) );
  NAND2_X1 U770 ( .A1(G61), .A2(n532), .ZN(n670) );
  NAND2_X1 U771 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U772 ( .A1(n672), .A2(G73), .ZN(n673) );
  XOR2_X1 U773 ( .A(KEYINPUT2), .B(n673), .Z(n674) );
  NOR2_X1 U774 ( .A1(n675), .A2(n674), .ZN(n678) );
  NAND2_X1 U775 ( .A1(n676), .A2(G48), .ZN(n677) );
  NAND2_X1 U776 ( .A1(n678), .A2(n677), .ZN(G305) );
  XOR2_X1 U777 ( .A(KEYINPUT80), .B(KEYINPUT19), .Z(n679) );
  XNOR2_X1 U778 ( .A(G288), .B(n679), .ZN(n680) );
  XNOR2_X1 U779 ( .A(n680), .B(G290), .ZN(n681) );
  XNOR2_X1 U780 ( .A(n681), .B(G299), .ZN(n682) );
  XNOR2_X1 U781 ( .A(n687), .B(n682), .ZN(n684) );
  XNOR2_X1 U782 ( .A(G305), .B(G166), .ZN(n683) );
  XNOR2_X1 U783 ( .A(n684), .B(n683), .ZN(n938) );
  XOR2_X1 U784 ( .A(n938), .B(n685), .Z(n686) );
  NOR2_X1 U785 ( .A1(n688), .A2(n686), .ZN(n690) );
  AND2_X1 U786 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U787 ( .A1(n690), .A2(n689), .ZN(G295) );
  NAND2_X1 U788 ( .A1(G2078), .A2(G2084), .ZN(n691) );
  XOR2_X1 U789 ( .A(KEYINPUT20), .B(n691), .Z(n692) );
  NAND2_X1 U790 ( .A1(G2090), .A2(n692), .ZN(n693) );
  XNOR2_X1 U791 ( .A(KEYINPUT21), .B(n693), .ZN(n694) );
  NAND2_X1 U792 ( .A1(n694), .A2(G2072), .ZN(n695) );
  XOR2_X1 U793 ( .A(KEYINPUT81), .B(n695), .Z(G158) );
  XNOR2_X1 U794 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  INV_X1 U795 ( .A(G661), .ZN(n705) );
  NOR2_X1 U796 ( .A1(G220), .A2(G219), .ZN(n696) );
  XOR2_X1 U797 ( .A(KEYINPUT22), .B(n696), .Z(n697) );
  NOR2_X1 U798 ( .A1(G218), .A2(n697), .ZN(n698) );
  NAND2_X1 U799 ( .A1(G96), .A2(n698), .ZN(n871) );
  NAND2_X1 U800 ( .A1(G2106), .A2(n871), .ZN(n702) );
  NAND2_X1 U801 ( .A1(G69), .A2(G120), .ZN(n699) );
  NOR2_X1 U802 ( .A1(G237), .A2(n699), .ZN(n700) );
  NAND2_X1 U803 ( .A1(G108), .A2(n700), .ZN(n872) );
  NAND2_X1 U804 ( .A1(G567), .A2(n872), .ZN(n701) );
  NAND2_X1 U805 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U806 ( .A(KEYINPUT82), .B(n703), .Z(n873) );
  NAND2_X1 U807 ( .A1(G483), .A2(n873), .ZN(n704) );
  NOR2_X1 U808 ( .A1(n705), .A2(n704), .ZN(n870) );
  NAND2_X1 U809 ( .A1(n870), .A2(G36), .ZN(G176) );
  INV_X1 U810 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U811 ( .A(KEYINPUT26), .B(KEYINPUT91), .ZN(n710) );
  NOR2_X2 U812 ( .A1(n706), .A2(G1384), .ZN(n813) );
  AND2_X1 U813 ( .A1(G1996), .A2(G40), .ZN(n707) );
  AND2_X1 U814 ( .A1(n710), .A2(n709), .ZN(n708) );
  NAND2_X1 U815 ( .A1(n708), .A2(n520), .ZN(n714) );
  NAND2_X1 U816 ( .A1(n716), .A2(n709), .ZN(n712) );
  INV_X1 U817 ( .A(n710), .ZN(n711) );
  NAND2_X1 U818 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U819 ( .A1(n714), .A2(n713), .ZN(n718) );
  AND2_X1 U820 ( .A1(n813), .A2(G40), .ZN(n715) );
  NAND2_X1 U821 ( .A1(n520), .A2(n715), .ZN(n722) );
  NAND2_X1 U822 ( .A1(n722), .A2(G1341), .ZN(n717) );
  NAND2_X1 U823 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U824 ( .A(n720), .B(KEYINPUT64), .ZN(n726) );
  NAND2_X1 U825 ( .A1(n726), .A2(n977), .ZN(n721) );
  XNOR2_X1 U826 ( .A(n721), .B(KEYINPUT92), .ZN(n725) );
  BUF_X1 U827 ( .A(n722), .Z(n755) );
  NOR2_X1 U828 ( .A1(n732), .A2(G1348), .ZN(n723) );
  INV_X1 U829 ( .A(G2067), .ZN(n1007) );
  NOR2_X1 U830 ( .A1(n726), .A2(n977), .ZN(n728) );
  NOR2_X1 U831 ( .A1(n730), .A2(n729), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n732), .A2(G2072), .ZN(n731) );
  XOR2_X1 U833 ( .A(KEYINPUT27), .B(n731), .Z(n734) );
  NAND2_X1 U834 ( .A1(G1956), .A2(n755), .ZN(n733) );
  NAND2_X1 U835 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U836 ( .A1(G299), .A2(n738), .ZN(n735) );
  NOR2_X1 U837 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U838 ( .A1(G299), .A2(n738), .ZN(n739) );
  XOR2_X1 U839 ( .A(n739), .B(KEYINPUT28), .Z(n740) );
  XNOR2_X1 U840 ( .A(n744), .B(n743), .ZN(n773) );
  OR2_X1 U841 ( .A1(n732), .A2(G1961), .ZN(n746) );
  XNOR2_X1 U842 ( .A(KEYINPUT25), .B(G2078), .ZN(n1015) );
  NAND2_X1 U843 ( .A1(n732), .A2(n1015), .ZN(n745) );
  NAND2_X1 U844 ( .A1(n746), .A2(n745), .ZN(n761) );
  AND2_X1 U845 ( .A1(n761), .A2(G171), .ZN(n747) );
  XOR2_X1 U846 ( .A(KEYINPUT90), .B(n747), .Z(n772) );
  NOR2_X1 U847 ( .A1(G1971), .A2(n810), .ZN(n749) );
  NOR2_X1 U848 ( .A1(G2090), .A2(n755), .ZN(n748) );
  NOR2_X1 U849 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U850 ( .A1(n750), .A2(G303), .ZN(n766) );
  INV_X1 U851 ( .A(n766), .ZN(n751) );
  OR2_X1 U852 ( .A1(n751), .A2(G286), .ZN(n752) );
  AND2_X1 U853 ( .A1(n772), .A2(n754), .ZN(n753) );
  NAND2_X1 U854 ( .A1(n773), .A2(n753), .ZN(n770) );
  INV_X1 U855 ( .A(n754), .ZN(n768) );
  XNOR2_X1 U856 ( .A(n756), .B(KEYINPUT89), .ZN(n777) );
  NAND2_X1 U857 ( .A1(G8), .A2(n777), .ZN(n757) );
  NOR2_X1 U858 ( .A1(n776), .A2(n757), .ZN(n758) );
  XNOR2_X1 U859 ( .A(n758), .B(KEYINPUT30), .ZN(n760) );
  AND2_X1 U860 ( .A1(n760), .A2(n759), .ZN(n763) );
  NOR2_X1 U861 ( .A1(G171), .A2(n761), .ZN(n762) );
  NOR2_X1 U862 ( .A1(n763), .A2(n762), .ZN(n765) );
  XNOR2_X1 U863 ( .A(n765), .B(n764), .ZN(n775) );
  AND2_X1 U864 ( .A1(n775), .A2(n766), .ZN(n767) );
  NAND2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n781) );
  INV_X1 U867 ( .A(n776), .ZN(n780) );
  INV_X1 U868 ( .A(n777), .ZN(n778) );
  NAND2_X1 U869 ( .A1(G8), .A2(n778), .ZN(n779) );
  NOR2_X2 U870 ( .A1(n783), .A2(n782), .ZN(n799) );
  INV_X1 U871 ( .A(n799), .ZN(n788) );
  NOR2_X1 U872 ( .A1(G1971), .A2(G303), .ZN(n784) );
  XOR2_X1 U873 ( .A(n784), .B(KEYINPUT96), .Z(n786) );
  NOR2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n1000) );
  NAND2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NOR2_X1 U877 ( .A1(n792), .A2(KEYINPUT33), .ZN(n796) );
  NAND2_X1 U878 ( .A1(n1000), .A2(KEYINPUT33), .ZN(n793) );
  XOR2_X1 U879 ( .A(KEYINPUT97), .B(n793), .Z(n794) );
  NOR2_X1 U880 ( .A1(n810), .A2(n794), .ZN(n795) );
  XNOR2_X1 U881 ( .A(n797), .B(KEYINPUT98), .ZN(n798) );
  XOR2_X1 U882 ( .A(G1981), .B(G305), .Z(n982) );
  NAND2_X1 U883 ( .A1(n798), .A2(n982), .ZN(n806) );
  BUF_X1 U884 ( .A(n799), .Z(n802) );
  NAND2_X1 U885 ( .A1(G166), .A2(G8), .ZN(n800) );
  NOR2_X1 U886 ( .A1(G2090), .A2(n800), .ZN(n801) );
  NOR2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U888 ( .A(n803), .B(KEYINPUT99), .ZN(n804) );
  NAND2_X1 U889 ( .A1(n804), .A2(n810), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U891 ( .A(n807), .B(KEYINPUT100), .ZN(n812) );
  NOR2_X1 U892 ( .A1(G1981), .A2(G305), .ZN(n808) );
  XOR2_X1 U893 ( .A(n808), .B(KEYINPUT24), .Z(n809) );
  NOR2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U895 ( .A1(n812), .A2(n811), .ZN(n846) );
  NAND2_X1 U896 ( .A1(G160), .A2(G40), .ZN(n814) );
  NOR2_X1 U897 ( .A1(n813), .A2(n814), .ZN(n861) );
  XNOR2_X1 U898 ( .A(G2067), .B(KEYINPUT37), .ZN(n859) );
  NAND2_X1 U899 ( .A1(G140), .A2(n913), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G104), .A2(n576), .ZN(n815) );
  NAND2_X1 U901 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U902 ( .A(KEYINPUT34), .B(n817), .ZN(n823) );
  NAND2_X1 U903 ( .A1(G116), .A2(n590), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G128), .A2(n916), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U906 ( .A(KEYINPUT84), .B(n820), .Z(n821) );
  XNOR2_X1 U907 ( .A(KEYINPUT35), .B(n821), .ZN(n822) );
  NOR2_X1 U908 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U909 ( .A(KEYINPUT36), .B(n824), .ZN(n927) );
  NOR2_X1 U910 ( .A1(n859), .A2(n927), .ZN(n953) );
  NAND2_X1 U911 ( .A1(n861), .A2(n953), .ZN(n857) );
  NAND2_X1 U912 ( .A1(G107), .A2(n590), .ZN(n826) );
  NAND2_X1 U913 ( .A1(G119), .A2(n916), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n826), .A2(n825), .ZN(n831) );
  NAND2_X1 U915 ( .A1(G131), .A2(n913), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G95), .A2(n576), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U918 ( .A(KEYINPUT85), .B(n829), .Z(n830) );
  NOR2_X1 U919 ( .A1(n831), .A2(n830), .ZN(n832) );
  XOR2_X1 U920 ( .A(KEYINPUT86), .B(n832), .Z(n925) );
  AND2_X1 U921 ( .A1(G1991), .A2(n925), .ZN(n842) );
  NAND2_X1 U922 ( .A1(G105), .A2(n576), .ZN(n833) );
  XNOR2_X1 U923 ( .A(n833), .B(KEYINPUT38), .ZN(n840) );
  NAND2_X1 U924 ( .A1(G129), .A2(n916), .ZN(n835) );
  NAND2_X1 U925 ( .A1(G141), .A2(n913), .ZN(n834) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n838) );
  NAND2_X1 U927 ( .A1(G117), .A2(n590), .ZN(n836) );
  XNOR2_X1 U928 ( .A(KEYINPUT87), .B(n836), .ZN(n837) );
  NOR2_X1 U929 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U930 ( .A1(n840), .A2(n839), .ZN(n926) );
  AND2_X1 U931 ( .A1(n926), .A2(G1996), .ZN(n841) );
  NOR2_X1 U932 ( .A1(n842), .A2(n841), .ZN(n962) );
  XOR2_X1 U933 ( .A(n861), .B(KEYINPUT88), .Z(n843) );
  NOR2_X1 U934 ( .A1(n962), .A2(n843), .ZN(n854) );
  INV_X1 U935 ( .A(n854), .ZN(n844) );
  NAND2_X1 U936 ( .A1(n857), .A2(n844), .ZN(n845) );
  NOR2_X2 U937 ( .A1(n846), .A2(n845), .ZN(n848) );
  XNOR2_X1 U938 ( .A(n848), .B(n847), .ZN(n850) );
  XNOR2_X1 U939 ( .A(G1986), .B(G290), .ZN(n996) );
  NAND2_X1 U940 ( .A1(n996), .A2(n861), .ZN(n849) );
  NAND2_X1 U941 ( .A1(n850), .A2(n849), .ZN(n864) );
  NOR2_X1 U942 ( .A1(G1996), .A2(n926), .ZN(n957) );
  NOR2_X1 U943 ( .A1(n925), .A2(G1991), .ZN(n851) );
  XNOR2_X1 U944 ( .A(n851), .B(KEYINPUT102), .ZN(n964) );
  NOR2_X1 U945 ( .A1(G1986), .A2(G290), .ZN(n852) );
  NOR2_X1 U946 ( .A1(n964), .A2(n852), .ZN(n853) );
  NOR2_X1 U947 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U948 ( .A1(n957), .A2(n855), .ZN(n856) );
  XNOR2_X1 U949 ( .A(KEYINPUT39), .B(n856), .ZN(n858) );
  NAND2_X1 U950 ( .A1(n858), .A2(n857), .ZN(n860) );
  NAND2_X1 U951 ( .A1(n859), .A2(n927), .ZN(n966) );
  NAND2_X1 U952 ( .A1(n860), .A2(n966), .ZN(n862) );
  NAND2_X1 U953 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U954 ( .A1(n864), .A2(n863), .ZN(n866) );
  XOR2_X1 U955 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n865) );
  XNOR2_X1 U956 ( .A(n866), .B(n865), .ZN(G329) );
  NAND2_X1 U957 ( .A1(G2106), .A2(n867), .ZN(G217) );
  AND2_X1 U958 ( .A1(G15), .A2(G2), .ZN(n868) );
  NAND2_X1 U959 ( .A1(G661), .A2(n868), .ZN(G259) );
  NAND2_X1 U960 ( .A1(G3), .A2(G1), .ZN(n869) );
  NAND2_X1 U961 ( .A1(n870), .A2(n869), .ZN(G188) );
  INV_X1 U963 ( .A(G120), .ZN(G236) );
  INV_X1 U964 ( .A(G96), .ZN(G221) );
  INV_X1 U965 ( .A(G69), .ZN(G235) );
  NOR2_X1 U966 ( .A1(n872), .A2(n871), .ZN(G325) );
  INV_X1 U967 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U968 ( .A(KEYINPUT104), .B(n873), .ZN(G319) );
  XNOR2_X1 U969 ( .A(G1996), .B(KEYINPUT41), .ZN(n883) );
  XOR2_X1 U970 ( .A(G1971), .B(G1961), .Z(n875) );
  XNOR2_X1 U971 ( .A(G1991), .B(G1956), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n879) );
  XOR2_X1 U973 ( .A(G1966), .B(G1976), .Z(n877) );
  XNOR2_X1 U974 ( .A(G1986), .B(G1981), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U976 ( .A(n879), .B(n878), .Z(n881) );
  XNOR2_X1 U977 ( .A(KEYINPUT108), .B(G2474), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(G229) );
  XNOR2_X1 U980 ( .A(G2067), .B(G2078), .ZN(n884) );
  XNOR2_X1 U981 ( .A(n884), .B(KEYINPUT42), .ZN(n894) );
  XOR2_X1 U982 ( .A(KEYINPUT107), .B(G2678), .Z(n886) );
  XNOR2_X1 U983 ( .A(KEYINPUT106), .B(G2096), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U985 ( .A(G2100), .B(G2090), .Z(n888) );
  XNOR2_X1 U986 ( .A(G2072), .B(G2084), .ZN(n887) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U988 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U989 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(G227) );
  NAND2_X1 U992 ( .A1(G112), .A2(n590), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G100), .A2(n576), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n902) );
  NAND2_X1 U995 ( .A1(n916), .A2(G124), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n897), .B(KEYINPUT44), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G136), .A2(n913), .ZN(n898) );
  NAND2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U999 ( .A(KEYINPUT109), .B(n900), .Z(n901) );
  NOR2_X1 U1000 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(KEYINPUT110), .B(n903), .ZN(G162) );
  XNOR2_X1 U1002 ( .A(KEYINPUT111), .B(KEYINPUT112), .ZN(n908) );
  NAND2_X1 U1003 ( .A1(G142), .A2(n913), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(G106), .A2(n576), .ZN(n904) );
  NAND2_X1 U1005 ( .A1(n905), .A2(n904), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n906), .B(KEYINPUT45), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(G118), .A2(n590), .ZN(n910) );
  NAND2_X1 U1009 ( .A1(G130), .A2(n916), .ZN(n909) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(n912), .A2(n911), .ZN(n923) );
  NAND2_X1 U1012 ( .A1(G139), .A2(n913), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(G103), .A2(n576), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n921) );
  NAND2_X1 U1015 ( .A1(G115), .A2(n590), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(G127), .A2(n916), .ZN(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT47), .B(n919), .Z(n920) );
  NOR2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n968) );
  XNOR2_X1 U1020 ( .A(n968), .B(G164), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n923), .B(n922), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n925), .B(n924), .ZN(n929) );
  XOR2_X1 U1023 ( .A(n927), .B(n926), .Z(n928) );
  XNOR2_X1 U1024 ( .A(n929), .B(n928), .ZN(n936) );
  XOR2_X1 U1025 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n930) );
  XNOR2_X1 U1026 ( .A(n954), .B(n930), .ZN(n931) );
  XOR2_X1 U1027 ( .A(n931), .B(KEYINPUT114), .Z(n933) );
  XNOR2_X1 U1028 ( .A(G160), .B(KEYINPUT48), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n933), .B(n932), .ZN(n934) );
  XOR2_X1 U1030 ( .A(G162), .B(n934), .Z(n935) );
  XNOR2_X1 U1031 ( .A(n936), .B(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(G37), .A2(n937), .ZN(G395) );
  XOR2_X1 U1033 ( .A(n938), .B(G286), .Z(n940) );
  XNOR2_X1 U1034 ( .A(n977), .B(G171), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(n940), .B(n939), .ZN(n941) );
  XNOR2_X1 U1036 ( .A(n941), .B(n986), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(G37), .A2(n942), .ZN(G397) );
  INV_X1 U1038 ( .A(G319), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(G401), .A2(n943), .ZN(n944) );
  XOR2_X1 U1040 ( .A(KEYINPUT115), .B(n944), .Z(n948) );
  NOR2_X1 U1041 ( .A1(G229), .A2(G227), .ZN(n945) );
  XOR2_X1 U1042 ( .A(KEYINPUT116), .B(n945), .Z(n946) );
  XNOR2_X1 U1043 ( .A(KEYINPUT49), .B(n946), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(KEYINPUT117), .B(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(G395), .A2(G397), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(G225) );
  INV_X1 U1048 ( .A(G225), .ZN(G308) );
  INV_X1 U1049 ( .A(G108), .ZN(G238) );
  INV_X1 U1050 ( .A(KEYINPUT55), .ZN(n1025) );
  XOR2_X1 U1051 ( .A(G160), .B(G2084), .Z(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n960) );
  XOR2_X1 U1054 ( .A(G2090), .B(G162), .Z(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1056 ( .A(n958), .B(KEYINPUT51), .ZN(n959) );
  NOR2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT118), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n973) );
  XOR2_X1 U1062 ( .A(G2072), .B(n968), .Z(n970) );
  XOR2_X1 U1063 ( .A(G164), .B(G2078), .Z(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1065 ( .A(KEYINPUT50), .B(n971), .Z(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(KEYINPUT52), .B(n974), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n1025), .A2(n975), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n976), .A2(G29), .ZN(n1032) );
  XOR2_X1 U1070 ( .A(KEYINPUT56), .B(G16), .Z(n1002) );
  XNOR2_X1 U1071 ( .A(G1348), .B(n977), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(n978), .B(KEYINPUT124), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n992) );
  XNOR2_X1 U1075 ( .A(G1966), .B(G168), .ZN(n981) );
  XNOR2_X1 U1076 ( .A(n981), .B(KEYINPUT122), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n984) );
  XNOR2_X1 U1079 ( .A(n985), .B(n984), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(n986), .B(G1341), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(G299), .B(G1956), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G166), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1030) );
  XNOR2_X1 U1091 ( .A(KEYINPUT54), .B(G34), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT121), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G2084), .B(n1004), .ZN(n1023) );
  XNOR2_X1 U1094 ( .A(G2090), .B(G35), .ZN(n1021) );
  XNOR2_X1 U1095 ( .A(G1991), .B(G25), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(G33), .B(G2072), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(G26), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(G28), .ZN(n1012) );
  INV_X1 U1100 ( .A(G1996), .ZN(n1009) );
  XOR2_X1 U1101 ( .A(G32), .B(n1009), .Z(n1010) );
  XNOR2_X1 U1102 ( .A(KEYINPUT120), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G27), .B(n1015), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT119), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT53), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1111 ( .A(n1025), .B(n1024), .ZN(n1027) );
  INV_X1 U1112 ( .A(G29), .ZN(n1026) );
  NAND2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(G11), .A2(n1028), .ZN(n1029) );
  NOR2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1058) );
  XNOR2_X1 U1117 ( .A(G1348), .B(KEYINPUT59), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(n1033), .B(G4), .ZN(n1037) );
  XNOR2_X1 U1119 ( .A(G1981), .B(G6), .ZN(n1035) );
  XNOR2_X1 U1120 ( .A(G1341), .B(G19), .ZN(n1034) );
  NOR2_X1 U1121 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1122 ( .A1(n1037), .A2(n1036), .ZN(n1039) );
  XNOR2_X1 U1123 ( .A(G20), .B(G1956), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XOR2_X1 U1125 ( .A(KEYINPUT60), .B(n1040), .Z(n1042) );
  XNOR2_X1 U1126 ( .A(G1966), .B(G21), .ZN(n1041) );
  NOR2_X1 U1127 ( .A1(n1042), .A2(n1041), .ZN(n1043) );
  XOR2_X1 U1128 ( .A(KEYINPUT125), .B(n1043), .Z(n1051) );
  XNOR2_X1 U1129 ( .A(G1976), .B(G23), .ZN(n1045) );
  XNOR2_X1 U1130 ( .A(G22), .B(G1971), .ZN(n1044) );
  NOR2_X1 U1131 ( .A1(n1045), .A2(n1044), .ZN(n1046) );
  XOR2_X1 U1132 ( .A(KEYINPUT126), .B(n1046), .Z(n1048) );
  XNOR2_X1 U1133 ( .A(G1986), .B(G24), .ZN(n1047) );
  NOR2_X1 U1134 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  XNOR2_X1 U1135 ( .A(KEYINPUT58), .B(n1049), .ZN(n1050) );
  NAND2_X1 U1136 ( .A1(n1051), .A2(n1050), .ZN(n1053) );
  XNOR2_X1 U1137 ( .A(G5), .B(G1961), .ZN(n1052) );
  NOR2_X1 U1138 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  XOR2_X1 U1139 ( .A(KEYINPUT61), .B(n1054), .Z(n1055) );
  NOR2_X1 U1140 ( .A1(G16), .A2(n1055), .ZN(n1056) );
  XOR2_X1 U1141 ( .A(KEYINPUT127), .B(n1056), .Z(n1057) );
  NOR2_X1 U1142 ( .A1(n1058), .A2(n1057), .ZN(n1059) );
  XNOR2_X1 U1143 ( .A(n1059), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1144 ( .A(G311), .ZN(G150) );
endmodule

