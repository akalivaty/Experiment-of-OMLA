//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1224,
    new_n1225, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  INV_X1    g0011(.A(G58), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT65), .Z(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n217), .A2(KEYINPUT64), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT64), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n219), .A2(G1), .A3(G13), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n206), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n216), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n208), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n211), .B(new_n224), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  OAI211_X1 g0051(.A(G1), .B(G13), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G45), .ZN(new_n253));
  AOI21_X1  g0053(.A(G1), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n252), .A2(G274), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT72), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT72), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n252), .A2(new_n257), .A3(new_n254), .A4(G274), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G97), .ZN(new_n259));
  INV_X1    g0059(.A(G232), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G1698), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G226), .B2(G1698), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n259), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n250), .A2(new_n251), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n218), .B2(new_n220), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n256), .A2(new_n258), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT67), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n205), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n272), .A2(new_n252), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT73), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT73), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n272), .A2(new_n276), .A3(new_n252), .A4(new_n273), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G238), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n281), .B1(new_n269), .B2(new_n278), .ZN(new_n282));
  OAI21_X1  g0082(.A(G200), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(G20), .A2(G33), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G50), .B1(G20), .B2(new_n213), .ZN(new_n285));
  INV_X1    g0085(.A(G77), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n206), .A2(G33), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n218), .A2(new_n220), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n213), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT12), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n290), .A2(new_n294), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n206), .A2(G1), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(G68), .A3(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n292), .A2(new_n296), .A3(new_n297), .A4(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n283), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(G190), .B1(new_n279), .B2(KEYINPUT13), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT74), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n281), .B1(new_n279), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n269), .A2(new_n278), .A3(KEYINPUT74), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT79), .ZN(new_n311));
  AND2_X1   g0111(.A1(G226), .A2(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n263), .B2(new_n264), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT78), .ZN(new_n314));
  NAND2_X1  g0114(.A1(G33), .A2(G87), .ZN(new_n315));
  INV_X1    g0115(.A(G1698), .ZN(new_n316));
  OAI211_X1 g0116(.A(G223), .B(new_n316), .C1(new_n263), .C2(new_n264), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT78), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n318), .B(new_n312), .C1(new_n263), .C2(new_n264), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n314), .A2(new_n315), .A3(new_n317), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n268), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n272), .A2(G232), .A3(new_n252), .A4(new_n273), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  AND3_X1   g0123(.A1(new_n322), .A2(new_n323), .A3(new_n255), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n311), .B1(new_n321), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n255), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n321), .A2(new_n311), .A3(new_n324), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g0133(.A(KEYINPUT8), .B(G58), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n334), .A2(KEYINPUT77), .A3(new_n299), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT77), .B1(new_n334), .B2(new_n299), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n298), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n294), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n290), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n265), .B2(new_n206), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  NOR4_X1   g0142(.A1(new_n263), .A2(new_n264), .A3(new_n342), .A4(G20), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G58), .A2(G68), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT76), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n347), .A2(G58), .A3(G68), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n346), .A2(new_n348), .A3(new_n214), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(G20), .B1(G159), .B2(new_n284), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n340), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT75), .B1(new_n263), .B2(new_n264), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n250), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(new_n359), .A3(new_n206), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n343), .B1(new_n360), .B2(new_n342), .ZN(new_n361));
  OAI211_X1 g0161(.A(KEYINPUT16), .B(new_n350), .C1(new_n361), .C2(new_n213), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n339), .B1(new_n353), .B2(new_n362), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n333), .A2(KEYINPUT80), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT80), .B1(new_n333), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT17), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n339), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n356), .A2(new_n206), .A3(new_n358), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n342), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n213), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n349), .A2(G20), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n284), .A2(G159), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n352), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n290), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n350), .A2(KEYINPUT16), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n360), .A2(new_n342), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n370), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n379), .B2(G68), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n367), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n327), .B1(new_n268), .B2(new_n320), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  INV_X1    g0183(.A(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(new_n382), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(KEYINPUT18), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n381), .B2(new_n385), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT17), .B1(new_n333), .B2(new_n363), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n366), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(G169), .B1(new_n280), .B2(new_n282), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(KEYINPUT14), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n307), .A2(new_n308), .ZN(new_n396));
  INV_X1    g0196(.A(G179), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n280), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT14), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n400), .B(G169), .C1(new_n280), .C2(new_n282), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n310), .B(new_n393), .C1(new_n302), .C2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G50), .A2(G58), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n206), .B1(new_n404), .B2(new_n213), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT68), .ZN(new_n406));
  INV_X1    g0206(.A(new_n334), .ZN(new_n407));
  INV_X1    g0207(.A(new_n287), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n407), .A2(new_n408), .B1(G150), .B2(new_n284), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n340), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  OR2_X1    g0210(.A1(new_n410), .A2(KEYINPUT69), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n298), .A2(G50), .A3(new_n300), .ZN(new_n412));
  INV_X1    g0212(.A(G50), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n294), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n410), .B2(KEYINPUT69), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT9), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT70), .ZN(new_n420));
  XNOR2_X1  g0220(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n265), .A2(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G222), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n356), .A2(new_n358), .ZN(new_n424));
  INV_X1    g0224(.A(G223), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(G1698), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n423), .B1(new_n286), .B2(new_n424), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n268), .ZN(new_n428));
  INV_X1    g0228(.A(new_n255), .ZN(new_n429));
  INV_X1    g0229(.A(new_n274), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n429), .B1(new_n430), .B2(G226), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  INV_X1    g0233(.A(new_n417), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT9), .ZN(new_n435));
  INV_X1    g0235(.A(new_n432), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G190), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n421), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  OR2_X1    g0239(.A1(new_n433), .A2(KEYINPUT71), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT10), .B1(new_n433), .B2(KEYINPUT71), .ZN(new_n441));
  AND4_X1   g0241(.A1(new_n435), .A2(new_n440), .A3(new_n437), .A4(new_n441), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n439), .A2(KEYINPUT10), .B1(new_n442), .B2(new_n421), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n432), .A2(new_n384), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(G179), .B2(new_n432), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(new_n434), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n407), .A2(new_n284), .B1(G20), .B2(G77), .ZN(new_n448));
  XNOR2_X1  g0248(.A(KEYINPUT15), .B(G87), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n287), .B2(new_n449), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n290), .B1(new_n286), .B2(new_n294), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n298), .A2(G77), .A3(new_n300), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n422), .A2(G232), .B1(G107), .B2(new_n265), .ZN(new_n454));
  INV_X1    g0254(.A(G238), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n426), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n268), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n429), .B1(new_n430), .B2(G244), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n453), .B1(new_n460), .B2(G190), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(G200), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n397), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n459), .A2(new_n384), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(new_n453), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n403), .A2(new_n447), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n205), .A2(G45), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(G257), .A3(new_n252), .ZN(new_n474));
  OR2_X1    g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  NAND2_X1  g0275(.A1(KEYINPUT5), .A2(G41), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n477), .A2(G274), .A3(new_n252), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT81), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G244), .B(new_n316), .C1(new_n263), .C2(new_n264), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT4), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n424), .A2(KEYINPUT4), .A3(G244), .A4(new_n316), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n424), .A2(G250), .A3(G1698), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n268), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n474), .A2(KEYINPUT81), .A3(new_n478), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n481), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G190), .ZN(new_n493));
  INV_X1    g0293(.A(G107), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(KEYINPUT6), .A3(G97), .ZN(new_n495));
  INV_X1    g0295(.A(G97), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n496), .A2(new_n494), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n202), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n500));
  OAI21_X1  g0300(.A(G107), .B1(new_n341), .B2(new_n343), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n340), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n294), .A2(new_n496), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n205), .A2(G33), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n298), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n503), .B1(new_n505), .B2(new_n496), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n491), .A2(G200), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n493), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT82), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n491), .A2(G169), .ZN(new_n511));
  AND3_X1   g0311(.A1(new_n474), .A2(KEYINPUT81), .A3(new_n478), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT81), .B1(new_n474), .B2(new_n478), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(G179), .A3(new_n489), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n510), .B(new_n507), .C1(new_n511), .C2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n511), .A2(new_n515), .ZN(new_n517));
  INV_X1    g0317(.A(new_n507), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT82), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n509), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n477), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n252), .A2(G274), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(G270), .B1(new_n523), .B2(new_n477), .ZN(new_n524));
  OAI211_X1 g0324(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n525));
  OAI211_X1 g0325(.A(G257), .B(new_n316), .C1(new_n263), .C2(new_n264), .ZN(new_n526));
  INV_X1    g0326(.A(G303), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(new_n424), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n268), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n340), .A2(G116), .A3(new_n293), .A4(new_n504), .ZN(new_n531));
  INV_X1    g0331(.A(G116), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n294), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(G20), .B1(G33), .B2(G283), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n250), .A2(G97), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n535), .B1(G20), .B2(new_n532), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n536), .A2(new_n290), .A3(KEYINPUT20), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT20), .B1(new_n536), .B2(new_n290), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n531), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n530), .A2(new_n539), .A3(G169), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT21), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n530), .A2(G200), .ZN(new_n543));
  INV_X1    g0343(.A(new_n539), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n524), .A2(G190), .A3(new_n529), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n524), .A2(G179), .A3(new_n529), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n539), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n530), .A2(new_n539), .A3(KEYINPUT21), .A4(G169), .ZN(new_n549));
  AND4_X1   g0349(.A1(new_n542), .A2(new_n546), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n551));
  OAI211_X1 g0351(.A(G238), .B(new_n316), .C1(new_n263), .C2(new_n264), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n551), .B(new_n552), .C1(new_n250), .C2(new_n532), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n268), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n252), .A2(G274), .A3(new_n472), .ZN(new_n555));
  OAI211_X1 g0355(.A(G250), .B(new_n471), .C1(new_n267), .C2(new_n217), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n554), .A2(G190), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n206), .B1(new_n259), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(G87), .B2(new_n203), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n206), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n560), .B1(new_n287), .B2(new_n496), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(new_n290), .B1(new_n294), .B2(new_n449), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n298), .A2(G87), .A3(new_n504), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n557), .B1(new_n268), .B2(new_n553), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n330), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n559), .B1(new_n569), .B2(KEYINPUT83), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n554), .A2(new_n558), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT83), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n572), .A2(new_n573), .A3(new_n566), .A4(new_n567), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n449), .B2(new_n505), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n568), .A2(G169), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n554), .A2(new_n397), .A3(new_n558), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n570), .A2(new_n574), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT23), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n206), .B2(G107), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n494), .A2(KEYINPUT23), .A3(G20), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n408), .A2(G116), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n424), .A2(new_n206), .A3(G87), .ZN(new_n587));
  NOR2_X1   g0387(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n586), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n424), .A2(new_n206), .A3(G87), .A4(new_n588), .ZN(new_n591));
  AOI211_X1 g0391(.A(KEYINPUT24), .B(new_n584), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n587), .A2(new_n589), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n591), .A3(new_n585), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n593), .B1(new_n595), .B2(new_n583), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n290), .B1(new_n592), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n505), .A2(new_n494), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT25), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n293), .B2(G107), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n494), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n604));
  OAI211_X1 g0404(.A(G250), .B(new_n316), .C1(new_n263), .C2(new_n264), .ZN(new_n605));
  INV_X1    g0405(.A(G294), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n604), .B(new_n605), .C1(new_n250), .C2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT85), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n268), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n522), .A2(G264), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n609), .A2(new_n478), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n607), .B2(new_n268), .ZN(new_n612));
  OAI21_X1  g0412(.A(G169), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n607), .A2(new_n268), .B1(new_n522), .B2(G264), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n478), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n397), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n603), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n330), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n607), .A2(new_n268), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT85), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n620), .A2(new_n478), .A3(new_n609), .A4(new_n610), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n618), .B1(new_n621), .B2(G190), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n622), .A2(new_n597), .A3(new_n602), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n550), .A2(new_n579), .A3(new_n617), .A4(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n469), .A2(new_n520), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g0425(.A(new_n625), .B(KEYINPUT86), .Z(G372));
  NAND2_X1  g0426(.A1(new_n566), .A2(new_n567), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n566), .A2(KEYINPUT87), .A3(new_n567), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n559), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(new_n572), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n623), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n548), .A2(new_n549), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n542), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n637), .B2(new_n617), .ZN(new_n638));
  INV_X1    g0438(.A(new_n509), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n517), .A2(new_n518), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n510), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n517), .A2(KEYINPUT82), .A3(new_n518), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n638), .A2(new_n643), .B1(new_n575), .B2(new_n578), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(KEYINPUT26), .A3(new_n642), .A4(new_n579), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT88), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n517), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT88), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n647), .A2(new_n518), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n578), .A2(new_n575), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n633), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n645), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n644), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n468), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT89), .Z(new_n656));
  INV_X1    g0456(.A(new_n446), .ZN(new_n657));
  INV_X1    g0457(.A(new_n390), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n402), .A2(new_n302), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n466), .B2(new_n310), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n366), .A2(new_n392), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n657), .B1(new_n662), .B2(new_n443), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n544), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n636), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n550), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n673), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n617), .A2(new_n623), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n603), .A2(new_n671), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n617), .B2(new_n672), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n603), .A2(new_n616), .A3(new_n672), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n637), .A2(new_n671), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n679), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n683), .A2(new_n684), .A3(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n209), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G1), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n215), .B2(new_n690), .ZN(new_n693));
  XOR2_X1   g0493(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n694));
  XNOR2_X1  g0494(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n638), .A2(new_n643), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n650), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n516), .A2(new_n519), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT26), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(new_n699), .A3(new_n579), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n699), .B2(new_n652), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n672), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n520), .A2(new_n624), .A3(new_n671), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n568), .A2(new_n614), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n705), .A2(new_n547), .A3(new_n514), .A4(new_n489), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n492), .A2(KEYINPUT30), .A3(new_n547), .A4(new_n705), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n568), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n491), .A2(new_n530), .A3(new_n615), .A4(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n671), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT31), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(G330), .B1(new_n704), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n671), .B1(new_n644), .B2(new_n653), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT29), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n703), .A2(new_n718), .A3(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n695), .B1(new_n723), .B2(G1), .ZN(G364));
  NAND2_X1  g0524(.A1(new_n206), .A2(G13), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n253), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n689), .A2(new_n205), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n678), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G330), .B2(new_n676), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n222), .B1(G20), .B2(new_n384), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G13), .A2(G33), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n354), .A2(new_n359), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n688), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n253), .B2(new_n216), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n245), .B2(new_n253), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n209), .A2(new_n424), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT92), .Z(new_n743));
  AOI22_X1  g0543(.A1(new_n743), .A2(G355), .B1(new_n532), .B2(new_n688), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n736), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n731), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n206), .A2(new_n323), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(G179), .A3(new_n330), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n206), .A2(G190), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(G179), .A3(new_n330), .ZN(new_n750));
  OAI22_X1  g0550(.A1(new_n748), .A2(new_n212), .B1(new_n750), .B2(new_n286), .ZN(new_n751));
  NAND3_X1  g0551(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n752), .A2(new_n323), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n754), .A2(new_n213), .B1(new_n756), .B2(new_n413), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n206), .B1(new_n758), .B2(G190), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n751), .B(new_n757), .C1(G97), .C2(new_n760), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n206), .A2(KEYINPUT93), .A3(G190), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT93), .B1(new_n206), .B2(G190), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n762), .A2(new_n758), .A3(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G159), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT32), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n330), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n747), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G87), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n424), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT94), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n762), .A2(new_n763), .A3(new_n768), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n775), .A2(G107), .B1(new_n771), .B2(new_n772), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n761), .A2(new_n767), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n750), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n265), .B1(new_n769), .B2(new_n527), .ZN(new_n780));
  INV_X1    g0580(.A(new_n748), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n779), .B(new_n780), .C1(G322), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(KEYINPUT95), .B(G326), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n756), .A2(new_n783), .B1(new_n606), .B2(new_n759), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n784), .B1(new_n753), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n764), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G329), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n775), .A2(G283), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n782), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n746), .B1(new_n777), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n728), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n745), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n734), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n793), .B1(new_n676), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n730), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G396));
  NOR2_X1   g0597(.A1(new_n466), .A2(new_n671), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n453), .A2(new_n671), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n463), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n798), .B1(new_n466), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n719), .B(new_n801), .Z(new_n802));
  INV_X1    g0602(.A(new_n718), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n804), .A2(new_n792), .A3(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n532), .A2(new_n750), .B1(new_n769), .B2(new_n494), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n424), .B(new_n807), .C1(G294), .C2(new_n781), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n753), .A2(KEYINPUT96), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(G283), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n760), .A2(G97), .B1(G303), .B2(new_n755), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G87), .A2(new_n775), .B1(new_n787), .B2(G311), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n808), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n750), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G143), .A2(new_n781), .B1(new_n817), .B2(G159), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  INV_X1    g0619(.A(G150), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n819), .B2(new_n756), .C1(new_n820), .C2(new_n754), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT34), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n737), .B1(new_n212), .B2(new_n759), .C1(new_n764), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n822), .B2(new_n821), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n774), .A2(new_n213), .B1(new_n413), .B2(new_n769), .ZN(new_n828));
  XOR2_X1   g0628(.A(new_n828), .B(KEYINPUT97), .Z(new_n829));
  OAI21_X1  g0629(.A(new_n816), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n731), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n731), .A2(new_n732), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n792), .B1(new_n286), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n831), .B(new_n833), .C1(new_n801), .C2(new_n733), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n806), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(G384));
  OR2_X1    g0636(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n837), .A2(G116), .A3(new_n223), .A4(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT36), .Z(new_n840));
  INV_X1    g0640(.A(new_n215), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n841), .A2(G77), .A3(new_n348), .A4(new_n346), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n413), .A2(G68), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT98), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n205), .B(G13), .C1(new_n842), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n659), .A2(new_n671), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT80), .ZN(new_n849));
  INV_X1    g0649(.A(new_n332), .ZN(new_n850));
  AOI21_X1  g0650(.A(G200), .B1(new_n321), .B2(new_n328), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n850), .A2(new_n325), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n849), .B1(new_n852), .B2(new_n381), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n333), .A2(KEYINPUT80), .A3(new_n363), .ZN(new_n854));
  INV_X1    g0654(.A(new_n669), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n381), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT37), .B1(new_n381), .B2(new_n385), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n853), .A2(new_n854), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n362), .A2(new_n290), .A3(new_n375), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n332), .B1(G200), .B2(new_n382), .ZN(new_n860));
  OAI211_X1 g0660(.A(new_n859), .B(new_n367), .C1(new_n860), .C2(new_n325), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(new_n386), .A3(new_n856), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT99), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n858), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n864), .B1(new_n858), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n856), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n393), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(KEYINPUT38), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n374), .B1(new_n379), .B2(G68), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n290), .B(new_n362), .C1(new_n871), .C2(KEYINPUT16), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n669), .B1(new_n872), .B2(new_n367), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n393), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n367), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n385), .B2(new_n855), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n853), .A3(new_n854), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT37), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n858), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n874), .A2(KEYINPUT38), .A3(new_n879), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n870), .A2(new_n880), .A3(KEYINPUT39), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n874), .A2(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n874), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n882), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT100), .B1(new_n881), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n858), .A2(new_n863), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT99), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n858), .A2(new_n863), .A3(new_n864), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n869), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n884), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n882), .A3(new_n886), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n874), .B2(new_n879), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT39), .B1(new_n880), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT100), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n848), .B1(new_n888), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n798), .B1(new_n719), .B2(new_n801), .ZN(new_n900));
  INV_X1    g0700(.A(new_n310), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n302), .A2(new_n671), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n659), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n302), .B(new_n671), .C1(new_n402), .C2(new_n310), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n885), .A2(new_n886), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n906), .A2(new_n907), .B1(new_n658), .B2(new_n669), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n703), .A2(new_n721), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n468), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n664), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n910), .B(new_n913), .Z(new_n914));
  INV_X1    g0714(.A(G330), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n704), .A2(new_n717), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n469), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n801), .B1(new_n704), .B2(new_n717), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n918), .A2(new_n905), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n919), .B(new_n920), .C1(new_n880), .C2(new_n895), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n903), .A2(new_n904), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n922), .B(new_n801), .C1(new_n704), .C2(new_n717), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n893), .B2(new_n886), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n921), .B1(new_n924), .B2(new_n920), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n915), .B1(new_n917), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n917), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n914), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n726), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n928), .B1(new_n205), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n914), .A2(new_n927), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n846), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NOR2_X1   g0732(.A1(new_n649), .A2(new_n672), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n518), .A2(new_n671), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n933), .B1(new_n643), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n686), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT42), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n617), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n672), .B1(new_n938), .B2(new_n698), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n631), .A2(new_n672), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n575), .A3(new_n578), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n651), .B2(new_n941), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT101), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT102), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n683), .A2(new_n935), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT103), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n727), .A2(new_n205), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n686), .B1(new_n682), .B2(new_n685), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(new_n677), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n723), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT104), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n686), .A2(new_n684), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n935), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT44), .Z(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n935), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT45), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(new_n683), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n722), .B1(new_n960), .B2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n689), .B(KEYINPUT41), .Z(new_n969));
  OAI21_X1  g0769(.A(new_n955), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n950), .A2(KEYINPUT103), .A3(new_n951), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n954), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n449), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n736), .B1(new_n688), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n738), .A2(new_n240), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n792), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n748), .A2(new_n820), .B1(new_n750), .B2(new_n413), .ZN(new_n977));
  INV_X1    g0777(.A(new_n769), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n265), .B(new_n977), .C1(G58), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n812), .A2(G159), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n760), .A2(G68), .B1(G143), .B2(new_n755), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G77), .A2(new_n775), .B1(new_n787), .B2(G137), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT106), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT46), .B1(new_n978), .B2(G116), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT105), .ZN(new_n986));
  INV_X1    g0786(.A(G317), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n985), .A2(new_n986), .B1(new_n987), .B2(new_n764), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n986), .B2(new_n985), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n759), .A2(new_n494), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n978), .A2(KEYINPUT46), .A3(G116), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G311), .C2(new_n755), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n812), .A2(G294), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G303), .A2(new_n781), .B1(new_n817), .B2(G283), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n775), .A2(G97), .ZN(new_n995));
  INV_X1    g0795(.A(new_n737), .ZN(new_n996));
  AND3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n989), .A2(new_n992), .A3(new_n993), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n984), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n976), .B1(new_n794), .B2(new_n943), .C1(new_n1001), .C2(new_n746), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n972), .A2(new_n1002), .ZN(G387));
  INV_X1    g0803(.A(new_n955), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n682), .A2(new_n794), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n738), .B1(new_n237), .B2(new_n253), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n743), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n691), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n334), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1009));
  OAI21_X1  g0809(.A(KEYINPUT50), .B1(new_n334), .B2(G50), .ZN(new_n1010));
  AOI21_X1  g0810(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1009), .A2(new_n691), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1008), .A2(new_n1012), .B1(new_n494), .B2(new_n688), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n728), .B1(new_n1013), .B2(new_n736), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n787), .A2(G150), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n978), .A2(G77), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n995), .A2(new_n1015), .A3(new_n737), .A4(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT108), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n748), .A2(new_n413), .B1(new_n750), .B2(new_n213), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n407), .B2(new_n753), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n760), .A2(new_n973), .B1(G159), .B2(new_n755), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n737), .B1(new_n775), .B2(G116), .ZN(new_n1023));
  INV_X1    g0823(.A(G283), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n769), .A2(new_n606), .B1(new_n759), .B2(new_n1024), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT109), .Z(new_n1026));
  OAI22_X1  g0826(.A1(new_n748), .A2(new_n987), .B1(new_n750), .B2(new_n527), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(G322), .B2(new_n755), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n811), .B2(new_n778), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT48), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1026), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT49), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1023), .B1(new_n783), .B2(new_n764), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1022), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1014), .B1(new_n1036), .B2(new_n731), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n958), .A2(new_n1004), .B1(new_n1005), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n689), .B1(new_n723), .B2(new_n958), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n960), .B2(new_n1039), .ZN(G393));
  AOI21_X1  g0840(.A(new_n690), .B1(new_n960), .B2(new_n967), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n960), .B2(new_n967), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n334), .A2(new_n750), .B1(new_n769), .B2(new_n213), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n996), .B(new_n1043), .C1(G77), .C2(new_n760), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G87), .A2(new_n775), .B1(new_n787), .B2(G143), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(new_n413), .C2(new_n811), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n781), .A2(G159), .B1(G150), .B2(new_n755), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT51), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n769), .A2(new_n1024), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n265), .B1(new_n750), .B2(new_n606), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G116), .C2(new_n760), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(G107), .A2(new_n775), .B1(new_n787), .B2(G322), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n527), .C2(new_n811), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n781), .A2(G311), .B1(G317), .B2(new_n755), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n1046), .A2(new_n1048), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n731), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n735), .B1(new_n496), .B2(new_n209), .C1(new_n739), .C2(new_n248), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n728), .B1(new_n1058), .B2(KEYINPUT110), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(KEYINPUT110), .B2(new_n1058), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT111), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1057), .B(new_n1061), .C1(new_n935), .C2(new_n734), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n967), .B2(new_n1004), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1042), .A2(new_n1063), .ZN(G390));
  OAI21_X1  g0864(.A(new_n848), .B1(new_n900), .B2(new_n905), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n888), .A2(new_n898), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n918), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(G330), .A3(new_n922), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT112), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n893), .A2(new_n886), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n800), .A2(new_n466), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n672), .B(new_n1072), .C1(new_n697), .C2(new_n701), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n798), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n848), .B(new_n1071), .C1(new_n1075), .C2(new_n905), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1066), .A2(new_n1070), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1070), .B1(new_n1066), .B2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1004), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n888), .A2(new_n732), .A3(new_n898), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n792), .B1(new_n334), .B2(new_n832), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n769), .A2(new_n820), .ZN(new_n1082));
  XOR2_X1   g0882(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1083));
  XNOR2_X1  g0883(.A(new_n1082), .B(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G125), .B2(new_n787), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n413), .B2(new_n774), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n811), .A2(new_n819), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT54), .B(G143), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n424), .B1(new_n750), .B2(new_n1088), .C1(new_n824), .C2(new_n748), .ZN(new_n1089));
  INV_X1    g0889(.A(G128), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n756), .A2(new_n1090), .B1(new_n759), .B2(new_n765), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1086), .A2(new_n1087), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(KEYINPUT115), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(KEYINPUT115), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n748), .A2(new_n532), .B1(new_n750), .B2(new_n496), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n424), .B(new_n1095), .C1(G87), .C2(new_n978), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n812), .A2(G107), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n760), .A2(G77), .B1(G283), .B2(new_n755), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G68), .A2(new_n775), .B1(new_n787), .B2(G294), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1093), .A2(new_n1094), .A3(new_n1100), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1080), .B(new_n1081), .C1(new_n746), .C2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1079), .A2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n468), .A2(new_n803), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n912), .A2(new_n664), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1075), .A2(new_n1068), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n718), .A2(KEYINPUT113), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n718), .A2(KEYINPUT113), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n801), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n905), .B2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n905), .B1(new_n918), .B2(new_n915), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n900), .B1(new_n1068), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1106), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n690), .B1(new_n1104), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1070), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n894), .A2(new_n897), .A3(new_n896), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n897), .B1(new_n894), .B2(new_n896), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n654), .A2(new_n672), .A3(new_n801), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1074), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n847), .B1(new_n1120), .B2(new_n922), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1117), .A2(new_n1118), .A3(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1076), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1066), .A2(new_n1070), .A3(new_n1076), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1114), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1103), .B1(new_n1115), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G378));
  NOR2_X1   g0929(.A1(new_n434), .A2(new_n669), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n419), .B(KEYINPUT70), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n435), .A2(new_n433), .A3(new_n437), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT10), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n442), .A2(new_n421), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n657), .B(new_n1131), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1130), .B1(new_n443), .B2(new_n446), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT120), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n1138), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n925), .A2(G330), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n925), .B2(G330), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n1146), .B1(new_n899), .B2(new_n909), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n919), .B1(new_n870), .B2(new_n880), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT40), .B1(new_n885), .B2(new_n886), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1148), .A2(KEYINPUT40), .B1(new_n1149), .B2(new_n919), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n1150), .A2(new_n915), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n847), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n925), .A2(new_n1144), .A3(G330), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n908), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1147), .A2(KEYINPUT121), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT121), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n910), .A2(new_n1156), .A3(new_n1153), .A4(new_n1151), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1106), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1155), .B(new_n1157), .C1(new_n1126), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT57), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1106), .B1(new_n1104), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT122), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n899), .B2(new_n909), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1147), .A2(KEYINPUT122), .A3(new_n1154), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(KEYINPUT57), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1161), .A2(new_n1167), .A3(new_n689), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1155), .A2(new_n1157), .A3(new_n1004), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n832), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n728), .B1(new_n1170), .B2(G50), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n774), .A2(new_n212), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n781), .A2(G107), .B1(new_n760), .B2(G68), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n532), .B2(new_n756), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1172), .B(new_n1174), .C1(G283), .C2(new_n787), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n817), .A2(new_n973), .B1(G97), .B2(new_n753), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT117), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n996), .A2(new_n1016), .A3(new_n251), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT116), .Z(new_n1179));
  NAND3_X1  g0979(.A1(new_n1175), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n1181));
  NAND2_X1  g0981(.A1(new_n996), .A2(new_n251), .ZN(new_n1182));
  AOI21_X1  g0982(.A(G50), .B1(new_n250), .B2(new_n251), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1180), .A2(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n748), .A2(new_n1090), .B1(new_n769), .B2(new_n1088), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT119), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n817), .A2(G137), .B1(G125), .B2(new_n755), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n760), .A2(G150), .B1(G132), .B2(new_n753), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n775), .A2(G159), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1184), .B(new_n1194), .C1(new_n1181), .C2(new_n1180), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1171), .B1(new_n1195), .B2(new_n731), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1144), .B2(new_n733), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1169), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1168), .A2(new_n1199), .ZN(G375));
  OAI21_X1  g1000(.A(new_n728), .B1(new_n1170), .B2(G68), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n996), .B1(G50), .B2(new_n760), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1202), .B1(new_n824), .B2(new_n756), .C1(new_n811), .C2(new_n1088), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n820), .A2(new_n750), .B1(new_n769), .B2(new_n765), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n748), .A2(new_n819), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1172), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n1090), .B2(new_n764), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G77), .A2(new_n775), .B1(new_n787), .B2(G303), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n424), .B1(new_n817), .B2(G107), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n781), .A2(G283), .B1(new_n978), .B2(G97), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n760), .A2(new_n973), .B1(G294), .B2(new_n755), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n811), .A2(new_n532), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n1203), .A2(new_n1207), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1201), .B1(new_n1214), .B2(new_n731), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n922), .B2(new_n733), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1162), .B2(new_n955), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1114), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n1219), .A2(new_n969), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1162), .A2(new_n1158), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1218), .B1(new_n1220), .B2(new_n1222), .ZN(G381));
  OR2_X1    g1023(.A1(G393), .A2(G396), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1224), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G387), .A2(new_n1225), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1026(.A1(new_n670), .A2(G213), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1128), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G375), .C2(new_n1229), .ZN(G409));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1114), .A2(KEYINPUT60), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n689), .B1(new_n1232), .B2(new_n1221), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1232), .B2(new_n1221), .ZN(new_n1234));
  OR3_X1    g1034(.A1(new_n1234), .A2(new_n835), .A3(new_n1217), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n835), .B1(new_n1234), .B2(new_n1217), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1228), .A2(G2897), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1237), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1168), .A2(G378), .A3(new_n1199), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1159), .A2(new_n969), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1166), .A2(new_n1004), .A3(new_n1165), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1197), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1128), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1228), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1231), .B1(new_n1240), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(KEYINPUT125), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1249), .B(new_n1231), .C1(new_n1240), .C2(new_n1246), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n690), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1198), .B(new_n1128), .C1(new_n1253), .C2(new_n1167), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1245), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1252), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1241), .A2(KEYINPUT123), .A3(new_n1245), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1256), .A2(new_n1227), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT124), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1241), .A2(new_n1245), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1228), .B1(new_n1261), .B2(new_n1252), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1257), .A4(new_n1258), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT62), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1246), .A2(KEYINPUT62), .A3(new_n1257), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT126), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1251), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(KEYINPUT127), .ZN(new_n1269));
  XNOR2_X1  g1069(.A(G393), .B(G396), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(G390), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G387), .B(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1251), .B(new_n1274), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1269), .A2(new_n1273), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1240), .B1(new_n1262), .B2(new_n1258), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1257), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(new_n1277), .A2(new_n1273), .A3(new_n1278), .A4(KEYINPUT61), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1260), .A2(new_n1264), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1279), .B1(KEYINPUT63), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(new_n1128), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1241), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(new_n1284), .B(new_n1257), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(new_n1285), .B(new_n1273), .ZN(G402));
endmodule


