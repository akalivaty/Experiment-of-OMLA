//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:10 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT10), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(KEYINPUT65), .A2(G143), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(G146), .A3(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n192), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G146), .B1(new_n193), .B2(new_n194), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT1), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT78), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  AND2_X1   g019(.A1(KEYINPUT65), .A2(G143), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT65), .A2(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT78), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(G128), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n195), .A2(new_n197), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n201), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G101), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  AOI22_X1  g030(.A1(KEYINPUT77), .A2(new_n215), .B1(new_n216), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT77), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  AND4_X1   g033(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT3), .A4(G104), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n218), .A2(KEYINPUT3), .B1(new_n219), .B2(G104), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n214), .B(new_n217), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(G107), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(G104), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n214), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n190), .B1(new_n213), .B2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G101), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n230), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n205), .A2(G143), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n208), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n195), .A2(new_n235), .A3(new_n197), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n229), .A2(new_n240), .A3(G101), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n231), .A2(new_n238), .A3(new_n239), .A4(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n222), .A2(new_n226), .ZN(new_n243));
  OAI21_X1  g057(.A(G128), .B1(new_n196), .B2(new_n203), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n202), .B2(new_n232), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n200), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n246), .A3(KEYINPUT10), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G134), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT11), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n251), .B1(G134), .B2(new_n248), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n253), .A2(KEYINPUT11), .A3(G137), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT67), .A2(G131), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT11), .B1(new_n253), .B2(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n251), .A2(new_n248), .A3(G134), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n249), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(KEYINPUT79), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n265), .B1(new_n258), .B2(new_n262), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n228), .A2(new_n242), .A3(new_n247), .A4(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  XNOR2_X1  g083(.A(G110), .B(G140), .ZN(new_n270));
  INV_X1    g084(.A(G227), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(G953), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n270), .B(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n268), .A2(new_n269), .A3(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n228), .A2(new_n242), .A3(new_n247), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n263), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n268), .A2(new_n274), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT80), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n210), .A2(G128), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n209), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n212), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n227), .B1(new_n283), .B2(new_n200), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n206), .A2(new_n207), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n196), .B1(new_n285), .B2(G146), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n286), .A2(new_n199), .B1(new_n234), .B2(new_n244), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n227), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT12), .B(new_n263), .C1(new_n284), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n288), .B1(new_n213), .B2(new_n227), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT12), .B1(new_n292), .B2(new_n263), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n268), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  AOI22_X1  g108(.A1(new_n278), .A2(new_n280), .B1(new_n294), .B2(new_n273), .ZN(new_n295));
  OAI21_X1  g109(.A(G469), .B1(new_n295), .B2(G902), .ZN(new_n296));
  XOR2_X1   g110(.A(KEYINPUT71), .B(G902), .Z(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT81), .B(G469), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n268), .A2(new_n300), .A3(new_n274), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n291), .A2(new_n293), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n268), .B2(new_n274), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n274), .B1(new_n277), .B2(new_n268), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n297), .B(new_n299), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n189), .B1(new_n296), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G214), .B1(G237), .B2(G902), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n309), .B(KEYINPUT83), .Z(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT2), .A2(G113), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT70), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n313));
  INV_X1    g127(.A(G113), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(KEYINPUT70), .A2(KEYINPUT2), .A3(G113), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n311), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G119), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G116), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G119), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n317), .B(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n231), .A2(new_n323), .A3(new_n241), .ZN(new_n324));
  NOR3_X1   g138(.A1(new_n320), .A2(KEYINPUT5), .A3(G119), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n314), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT5), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n317), .A2(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n243), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n324), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(G110), .B(G122), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n329), .A3(new_n331), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT6), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n336), .A3(new_n332), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n287), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT65), .B(G143), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n232), .B1(new_n340), .B2(new_n205), .ZN(new_n341));
  INV_X1    g155(.A(new_n237), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n239), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G224), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n345), .B(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n335), .A2(new_n337), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT84), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT84), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n335), .A2(new_n351), .A3(new_n337), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n334), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n317), .A2(new_n322), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT85), .B1(new_n325), .B2(new_n314), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n327), .ZN(new_n358));
  NOR3_X1   g172(.A1(new_n325), .A2(KEYINPUT85), .A3(new_n314), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n243), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n331), .B(KEYINPUT8), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n227), .A2(new_n328), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT7), .B1(new_n346), .B2(G953), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n246), .A2(G125), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n338), .B1(new_n238), .B2(new_n239), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n339), .A2(new_n344), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n364), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n354), .B1(new_n355), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n353), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G210), .B1(G237), .B2(G902), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(KEYINPUT87), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n353), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n310), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G140), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n338), .A2(G140), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT16), .ZN(new_n385));
  OR3_X1    g199(.A1(new_n338), .A2(KEYINPUT16), .A3(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G146), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n384), .A3(KEYINPUT88), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT19), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n391), .B2(new_n205), .ZN(new_n392));
  INV_X1    g206(.A(G237), .ZN(new_n393));
  INV_X1    g207(.A(G953), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G143), .A4(G214), .ZN(new_n395));
  INV_X1    g209(.A(G214), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n396), .A2(G237), .A3(G953), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n395), .B1(new_n340), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G131), .ZN(new_n399));
  INV_X1    g213(.A(G131), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(new_n395), .C1(new_n340), .C2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n398), .B(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n383), .A2(new_n384), .A3(new_n205), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT74), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n383), .A2(new_n384), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G146), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n403), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  XOR2_X1   g228(.A(G113), .B(G122), .Z(new_n415));
  XOR2_X1   g229(.A(KEYINPUT89), .B(G104), .Z(new_n416));
  XOR2_X1   g230(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n392), .A2(new_n402), .B1(new_n405), .B2(new_n411), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT90), .B1(new_n420), .B2(new_n417), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT17), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n399), .A2(new_n401), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT91), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n385), .A2(new_n386), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n205), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(KEYINPUT72), .A3(new_n387), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT72), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(new_n205), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n398), .A2(KEYINPUT17), .A3(G131), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n399), .A2(new_n401), .A3(KEYINPUT91), .A4(new_n422), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n425), .A2(new_n431), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(new_n417), .A3(new_n412), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n419), .A2(new_n421), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(G475), .A2(G902), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT20), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n436), .A2(new_n440), .A3(new_n437), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n394), .A2(G952), .ZN(new_n443));
  INV_X1    g257(.A(G234), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n393), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI211_X1 g260(.A(new_n394), .B(new_n297), .C1(G234), .C2(G237), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(G898), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G478), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n451), .A2(KEYINPUT15), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G217), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n187), .A2(new_n454), .A3(G953), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G116), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n320), .A2(G122), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n219), .B1(new_n460), .B2(KEYINPUT14), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n219), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n459), .A2(new_n461), .B1(new_n462), .B2(KEYINPUT94), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n462), .A2(KEYINPUT94), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n192), .A2(G128), .ZN(new_n465));
  AOI211_X1 g279(.A(G134), .B(new_n465), .C1(new_n285), .C2(G128), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n285), .A2(G128), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n253), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n463), .B(new_n464), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n457), .B(new_n219), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n467), .A2(new_n253), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n467), .B1(new_n475), .B2(new_n465), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n285), .A2(KEYINPUT13), .A3(G128), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G134), .B1(new_n478), .B2(new_n477), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n474), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n456), .B1(new_n471), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT93), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n480), .B1(new_n485), .B2(new_n476), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n470), .B(new_n455), .C1(new_n486), .C2(new_n474), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n453), .B1(new_n488), .B2(new_n297), .ZN(new_n489));
  INV_X1    g303(.A(new_n297), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n490), .B(new_n452), .C1(new_n483), .C2(new_n487), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n435), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n417), .B1(new_n434), .B2(new_n412), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n354), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT92), .B(G475), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n442), .A2(new_n450), .A3(new_n492), .A4(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n308), .A2(new_n381), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(G472), .ZN(new_n501));
  INV_X1    g315(.A(new_n323), .ZN(new_n502));
  AOI211_X1 g316(.A(G131), .B(new_n249), .C1(new_n259), .C2(new_n260), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT68), .B1(new_n248), .B2(G134), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT68), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n253), .A3(G137), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n248), .A2(G134), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n400), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n246), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n255), .A2(new_n257), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n261), .A2(new_n256), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n238), .B(new_n239), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n502), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT28), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT28), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n502), .A2(new_n511), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n343), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n238), .A2(KEYINPUT66), .A3(new_n239), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n263), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n400), .B(new_n250), .C1(new_n252), .C2(new_n254), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n504), .A2(new_n506), .B1(G134), .B2(new_n248), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n400), .B2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n287), .A2(new_n525), .A3(KEYINPUT69), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT69), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n510), .B2(new_n246), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n522), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n516), .A2(new_n518), .B1(new_n529), .B2(new_n323), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n393), .A2(new_n394), .A3(G210), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT27), .Z(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT26), .B(G101), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  AOI21_X1  g348(.A(KEYINPUT29), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n515), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT30), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n537), .B1(new_n529), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n539), .B2(new_n323), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n535), .B1(new_n534), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n516), .A2(new_n518), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n511), .A2(new_n514), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n323), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n542), .A2(KEYINPUT29), .A3(new_n534), .A4(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n545), .A2(new_n297), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n501), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT32), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n530), .A2(new_n534), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT31), .B1(new_n540), .B2(new_n534), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n511), .A2(new_n514), .A3(KEYINPUT30), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT69), .B1(new_n287), .B2(new_n525), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n510), .A2(new_n527), .A3(new_n246), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n343), .A2(new_n519), .B1(new_n258), .B2(new_n262), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n554), .A2(new_n555), .B1(new_n556), .B2(new_n521), .ZN(new_n557));
  INV_X1    g371(.A(new_n538), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n323), .B(new_n553), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n559), .A2(KEYINPUT31), .A3(new_n515), .A4(new_n534), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n551), .B1(new_n552), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n549), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n559), .A2(new_n515), .A3(new_n534), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT31), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n550), .B1(new_n567), .B2(new_n560), .ZN(new_n568));
  INV_X1    g382(.A(new_n563), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n568), .A2(KEYINPUT32), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n548), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n394), .A2(G221), .A3(G234), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  NAND2_X1  g388(.A1(new_n318), .A2(G128), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n198), .A2(G119), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT24), .B(G110), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n318), .A2(G128), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n575), .B(new_n580), .C1(new_n581), .C2(KEYINPUT23), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n579), .B1(G110), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n428), .A2(new_n430), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n577), .A2(new_n578), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT73), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n582), .A2(G110), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n387), .B(new_n408), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n584), .A2(new_n591), .A3(KEYINPUT75), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT75), .B1(new_n584), .B2(new_n591), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n574), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n574), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n584), .A2(new_n591), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n454), .B1(new_n297), .B2(G234), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n599), .A2(G902), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n594), .A2(new_n297), .A3(new_n598), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT76), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT25), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n601), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n571), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n500), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n214), .ZN(G3));
  AND3_X1   g426(.A1(new_n353), .A2(new_n379), .A3(new_n374), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n379), .B1(new_n353), .B2(new_n374), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n450), .B(new_n309), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n436), .A2(new_n440), .A3(new_n437), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n440), .B1(new_n436), .B2(new_n437), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n497), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n490), .A2(new_n451), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n488), .A2(KEYINPUT33), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT33), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n483), .B2(new_n487), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n488), .A2(new_n297), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT95), .B(G478), .Z(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT96), .B1(new_n615), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n309), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n378), .B2(new_n380), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  INV_X1    g446(.A(new_n628), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n450), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(G472), .B1(new_n568), .B2(new_n490), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n562), .A2(new_n563), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n637), .A3(new_n609), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n308), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(new_n492), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n442), .A2(new_n644), .A3(new_n497), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n615), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  AND2_X1   g463(.A1(new_n636), .A2(new_n637), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n600), .A2(G902), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n596), .B(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n607), .A2(new_n608), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n498), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n308), .A2(new_n650), .A3(new_n381), .A4(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT37), .B(G110), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G12));
  NAND2_X1  g472(.A1(new_n607), .A2(new_n608), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n653), .A2(new_n651), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n446), .B1(new_n447), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n645), .A2(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n571), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n263), .B1(new_n284), .B2(new_n289), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT12), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n279), .A2(KEYINPUT82), .B1(new_n290), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n306), .B1(new_n669), .B2(new_n301), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n670), .A2(new_n490), .A3(new_n298), .ZN(new_n671));
  INV_X1    g485(.A(G469), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n280), .A2(new_n277), .A3(new_n275), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n294), .A2(new_n273), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n672), .B1(new_n675), .B2(new_n354), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n188), .B1(new_n671), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n309), .B1(new_n613), .B2(new_n614), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n665), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G128), .ZN(G30));
  NAND2_X1  g495(.A1(new_n378), .A2(new_n380), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT38), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n309), .B1(new_n489), .B2(new_n491), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n442), .B2(new_n497), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n683), .A2(new_n654), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n663), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n308), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  INV_X1    g504(.A(new_n534), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n540), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n536), .A2(new_n534), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n693), .B2(new_n544), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n696), .B1(new_n564), .B2(new_n570), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n686), .A2(new_n689), .A3(new_n690), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(new_n340), .ZN(G45));
  INV_X1    g513(.A(new_n663), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n618), .A2(new_n627), .A3(new_n700), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n654), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n571), .A2(new_n308), .A3(new_n631), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT97), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n562), .A2(new_n549), .A3(new_n563), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT32), .B1(new_n568), .B2(new_n569), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n547), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n618), .A2(new_n627), .A3(new_n700), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n661), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT97), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n710), .A2(new_n679), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n704), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  OAI21_X1  g528(.A(G469), .B1(new_n670), .B2(new_n490), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(new_n307), .A3(new_n188), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT98), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT98), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n307), .A3(new_n718), .A4(new_n188), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n717), .A2(new_n571), .A3(new_n609), .A4(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n635), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT99), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT41), .B(G113), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND2_X1  g539(.A1(new_n721), .A2(new_n646), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  AND3_X1   g541(.A1(new_n717), .A2(new_n631), .A3(new_n719), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n707), .A2(new_n498), .A3(new_n654), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n618), .A2(new_n644), .A3(new_n309), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n378), .B2(new_n380), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n562), .A2(new_n297), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n542), .A2(new_n544), .ZN(new_n736));
  OAI22_X1  g550(.A1(new_n552), .A2(new_n561), .B1(new_n534), .B2(new_n736), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n735), .A2(G472), .B1(new_n563), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n734), .A2(new_n738), .A3(new_n609), .A4(new_n450), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n717), .A2(new_n719), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n732), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n450), .B(new_n685), .C1(new_n613), .C2(new_n614), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n737), .A2(new_n563), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n636), .A3(new_n609), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(KEYINPUT100), .A3(new_n719), .A4(new_n717), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n741), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  NAND2_X1  g562(.A1(new_n743), .A2(new_n636), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n654), .A3(new_n701), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n728), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  NAND3_X1  g566(.A1(new_n378), .A2(new_n380), .A3(new_n309), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n189), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT101), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n673), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n278), .A2(KEYINPUT101), .A3(new_n280), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(G469), .A3(new_n674), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n672), .A2(new_n354), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(new_n307), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n609), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n707), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT103), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n701), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n766), .B1(KEYINPUT102), .B2(new_n767), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n763), .A2(new_n765), .A3(new_n768), .A4(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n765), .A2(new_n762), .A3(new_n754), .A4(new_n768), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n769), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n771), .A2(new_n773), .A3(KEYINPUT104), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT104), .B1(new_n771), .B2(new_n773), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G131), .ZN(G33));
  NAND4_X1  g591(.A1(new_n765), .A2(new_n664), .A3(new_n754), .A4(new_n762), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  NAND3_X1  g593(.A1(new_n758), .A2(KEYINPUT45), .A3(new_n674), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n672), .B1(new_n675), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(KEYINPUT105), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT105), .B1(new_n780), .B2(new_n782), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n761), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT46), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n671), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n780), .A2(new_n782), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT105), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n760), .B1(new_n791), .B2(new_n783), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n189), .B1(new_n788), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n627), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n795), .A2(new_n618), .A3(KEYINPUT43), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n795), .B1(KEYINPUT106), .B2(new_n618), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(KEYINPUT106), .B2(new_n618), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n796), .B1(new_n798), .B2(KEYINPUT43), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n650), .A2(new_n654), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(KEYINPUT44), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT44), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n753), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n794), .A2(new_n687), .A3(new_n801), .A4(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(KEYINPUT107), .B(G137), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(G39));
  OAI21_X1  g620(.A(new_n307), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n786), .A2(new_n787), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n188), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(KEYINPUT47), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n188), .B(new_n814), .C1(new_n807), .C2(new_n808), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n571), .A2(new_n753), .A3(new_n609), .A4(new_n701), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  INV_X1    g632(.A(KEYINPUT51), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n799), .A2(new_n446), .ZN(new_n820));
  INV_X1    g634(.A(new_n744), .ZN(new_n821));
  INV_X1    g635(.A(new_n753), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT113), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n812), .A2(new_n815), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n715), .A2(new_n307), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n189), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n825), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT50), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n820), .A2(new_n821), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n683), .A2(new_n309), .ZN(new_n833));
  INV_X1    g647(.A(new_n740), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n831), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n799), .A2(new_n446), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n744), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n838), .A2(KEYINPUT50), .A3(new_n834), .A4(new_n833), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n834), .A2(new_n822), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n837), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n842), .A2(new_n661), .A3(new_n738), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n697), .A2(new_n764), .A3(new_n445), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n439), .A2(new_n441), .B1(new_n495), .B2(new_n496), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n795), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n840), .B(new_n843), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n819), .B1(new_n830), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT114), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n819), .C1(new_n830), .C2(new_n848), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OR3_X1    g667(.A1(new_n830), .A2(new_n848), .A3(new_n819), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n845), .A2(new_n628), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n838), .A2(new_n728), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n443), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n858), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n842), .A2(new_n765), .ZN(new_n861));
  XOR2_X1   g675(.A(new_n861), .B(KEYINPUT48), .Z(new_n862));
  NOR3_X1   g676(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n853), .A2(new_n854), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n734), .A2(new_n188), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT111), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n661), .B2(new_n663), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n654), .A2(KEYINPUT111), .A3(new_n700), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n866), .A2(new_n697), .A3(new_n762), .A4(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n713), .A2(new_n680), .A3(new_n751), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n704), .A2(new_n712), .B1(new_n679), .B2(new_n665), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n751), .A4(new_n871), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n721), .A2(new_n646), .B1(new_n728), .B2(new_n729), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n449), .B1(new_n628), .B2(new_n645), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n638), .A2(new_n381), .A3(new_n308), .A4(new_n879), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n880), .B(new_n656), .C1(new_n610), .C2(new_n500), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n878), .A2(new_n882), .A3(new_n747), .A4(new_n722), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n846), .A2(KEYINPUT110), .A3(new_n492), .A4(new_n700), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT110), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n492), .B(new_n497), .C1(new_n616), .C2(new_n617), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n663), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n753), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n571), .A3(new_n308), .A4(new_n661), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n750), .A2(new_n754), .A3(new_n762), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n778), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n883), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n877), .A2(new_n894), .A3(new_n776), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT53), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n720), .B1(new_n634), .B2(new_n629), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n881), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n747), .A3(new_n878), .A4(new_n892), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n901), .B1(new_n874), .B2(new_n876), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n771), .A2(KEYINPUT53), .A3(new_n773), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT112), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n895), .A2(new_n906), .A3(new_n896), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n906), .B1(new_n895), .B2(new_n896), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n895), .A2(new_n896), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n905), .B1(new_n910), .B2(new_n898), .ZN(new_n911));
  OAI22_X1  g725(.A1(new_n864), .A2(new_n911), .B1(G952), .B2(G953), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n764), .A2(new_n189), .A3(new_n310), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT109), .Z(new_n914));
  OR2_X1    g728(.A1(new_n827), .A2(KEYINPUT49), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n683), .A2(new_n798), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n697), .B1(new_n827), .B2(KEYINPUT49), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n918), .ZN(G75));
  INV_X1    g733(.A(KEYINPUT116), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n877), .A2(new_n894), .A3(new_n903), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n896), .B2(new_n895), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(new_n297), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n897), .A2(new_n904), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(KEYINPUT116), .A3(new_n490), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n377), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n335), .A2(new_n337), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(new_n348), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT55), .Z(new_n930));
  OAI21_X1  g744(.A(new_n927), .B1(new_n930), .B2(KEYINPUT118), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(KEYINPUT118), .B2(new_n930), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n394), .A2(G952), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT119), .Z(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n924), .A2(new_n490), .A3(new_n377), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT56), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n936), .B1(new_n939), .B2(new_n930), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n933), .A2(new_n940), .ZN(G51));
  AND3_X1   g755(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n898), .B1(new_n897), .B2(new_n904), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n760), .B(KEYINPUT57), .Z(new_n945));
  OAI22_X1  g759(.A1(new_n944), .A2(new_n945), .B1(new_n306), .B2(new_n305), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n923), .A2(new_n791), .A3(new_n783), .A4(new_n925), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n934), .B1(new_n946), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n923), .A2(new_n925), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n436), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(new_n934), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n923), .A2(new_n436), .A3(new_n925), .A4(new_n949), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(G60));
  OR2_X1    g769(.A1(new_n620), .A2(new_n622), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT120), .Z(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT59), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT53), .B1(new_n902), .B2(new_n776), .ZN(new_n961));
  OAI21_X1  g775(.A(KEYINPUT54), .B1(new_n961), .B2(new_n921), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n962), .B2(new_n905), .ZN(new_n963));
  OAI21_X1  g777(.A(KEYINPUT121), .B1(new_n963), .B2(new_n936), .ZN(new_n964));
  INV_X1    g778(.A(new_n960), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n942), .B2(new_n943), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n967), .A3(new_n935), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n964), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n957), .B1(new_n911), .B2(new_n959), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G63));
  NAND2_X1  g785(.A1(G217), .A2(G902), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n924), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n599), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n924), .A2(new_n653), .A3(new_n974), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n935), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(KEYINPUT61), .B1(new_n977), .B2(KEYINPUT123), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G66));
  OAI21_X1  g794(.A(G953), .B1(new_n448), .B2(new_n346), .ZN(new_n981));
  INV_X1    g795(.A(new_n883), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n928), .B1(G898), .B2(new_n394), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  NAND3_X1  g800(.A1(new_n713), .A2(new_n680), .A3(new_n751), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n778), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n794), .A2(new_n765), .A3(new_n687), .A4(new_n734), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n989), .A2(new_n776), .A3(new_n804), .A4(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n817), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n991), .A2(new_n992), .A3(KEYINPUT126), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT126), .B1(new_n991), .B2(new_n992), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n394), .A3(new_n994), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n539), .B(new_n391), .Z(new_n996));
  AOI21_X1  g810(.A(new_n996), .B1(G900), .B2(G953), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(G953), .B1(new_n271), .B2(new_n662), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n999), .A2(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n988), .A2(new_n698), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n628), .A2(new_n645), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT125), .Z(new_n1005));
  OR4_X1    g819(.A1(new_n610), .A2(new_n1005), .A3(new_n688), .A4(new_n753), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n804), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1003), .A2(new_n817), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n394), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1000), .B1(new_n1009), .B2(new_n996), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n999), .A2(KEYINPUT127), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n998), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1011), .B1(new_n998), .B2(new_n1010), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1012), .A2(new_n1013), .ZN(G72));
  NAND2_X1  g828(.A1(new_n559), .A2(new_n693), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n993), .A2(new_n982), .A3(new_n994), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  AOI21_X1  g832(.A(new_n1015), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n1008), .B2(new_n883), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n1020), .A2(new_n692), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n540), .B(new_n534), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n1018), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n910), .A2(new_n1023), .ZN(new_n1024));
  NOR4_X1   g838(.A1(new_n1019), .A2(new_n1021), .A3(new_n1024), .A4(new_n934), .ZN(G57));
endmodule


