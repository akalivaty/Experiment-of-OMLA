//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:31 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT64), .Z(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT65), .B(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G107), .A2(G264), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT67), .B(G50), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  NAND3_X1  g0047(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(new_n217), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n252), .B(G50), .C1(G1), .C2(new_n208), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G50), .B2(new_n248), .ZN(new_n254));
  INV_X1    g0054(.A(new_n251), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n208), .B1(new_n201), .B2(new_n202), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n208), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n260), .A2(new_n262), .B1(G150), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n255), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G169), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G1698), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n270), .B1(new_n203), .B2(new_n268), .C1(new_n271), .C2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  INV_X1    g0080(.A(G45), .ZN(new_n281));
  AOI21_X1  g0081(.A(G1), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(new_n284), .A3(G274), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n286), .B1(G226), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n279), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n266), .B1(new_n267), .B2(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G179), .B2(new_n291), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g0094(.A1(KEYINPUT9), .A2(new_n266), .B1(new_n291), .B2(G200), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n295), .B1(KEYINPUT9), .B2(new_n266), .C1(new_n296), .C2(new_n291), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n248), .A2(KEYINPUT70), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT70), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n302), .A2(new_n207), .A3(G13), .A4(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n251), .B1(new_n301), .B2(new_n303), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n305), .A2(new_n203), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n263), .ZN(new_n309));
  OAI22_X1  g0109(.A1(new_n259), .A2(new_n309), .B1(new_n208), .B2(new_n203), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT15), .B(G87), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT69), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n312), .B2(new_n262), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n308), .B1(new_n313), .B2(new_n255), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n286), .B1(G244), .B2(new_n289), .ZN(new_n315));
  INV_X1    g0115(.A(G107), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n276), .A2(new_n220), .B1(new_n268), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n273), .A2(new_n275), .ZN(new_n318));
  INV_X1    g0118(.A(G232), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n278), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G179), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n315), .A2(new_n321), .A3(KEYINPUT71), .A4(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(G169), .B1(new_n315), .B2(new_n321), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n315), .A2(new_n321), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n325), .A2(new_n326), .B1(new_n327), .B2(G179), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n324), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n314), .B1(G200), .B2(new_n327), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n296), .B2(new_n327), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n300), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n268), .A2(G226), .A3(new_n269), .ZN(new_n334));
  NAND2_X1  g0134(.A1(G33), .A2(G97), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n278), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n286), .B1(G238), .B2(new_n289), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n337), .B2(new_n338), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT14), .B1(new_n342), .B2(new_n267), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(G169), .C1(new_n340), .C2(new_n341), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT74), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n342), .B2(G179), .ZN(new_n347));
  NOR4_X1   g0147(.A1(new_n340), .A2(new_n341), .A3(KEYINPUT74), .A4(new_n322), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n343), .B(new_n345), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n221), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n203), .B2(new_n261), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n351), .A2(KEYINPUT72), .A3(new_n251), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT72), .B1(new_n351), .B2(new_n251), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n352), .A2(new_n353), .A3(KEYINPUT11), .ZN(new_n354));
  INV_X1    g0154(.A(G13), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G1), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT12), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(G20), .A4(new_n221), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT73), .Z(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT12), .B1(new_n304), .B2(G68), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n221), .B1(new_n207), .B2(G20), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n359), .A2(new_n360), .B1(new_n306), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT11), .B1(new_n352), .B2(new_n353), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n354), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n349), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n342), .A2(G190), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n337), .A2(new_n338), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT13), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G200), .ZN(new_n371));
  INV_X1    g0171(.A(new_n364), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n366), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n268), .A2(new_n376), .A3(G20), .ZN(new_n377));
  AOI21_X1  g0177(.A(KEYINPUT7), .B1(new_n318), .B2(new_n208), .ZN(new_n378));
  OAI21_X1  g0178(.A(G68), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n263), .A2(G159), .ZN(new_n380));
  INV_X1    g0180(.A(G58), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n221), .ZN(new_n382));
  OAI21_X1  g0182(.A(G20), .B1(new_n382), .B2(new_n201), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n379), .A2(KEYINPUT16), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n376), .B1(new_n268), .B2(G20), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n318), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n221), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n383), .A2(new_n380), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n384), .A2(new_n390), .A3(new_n251), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n259), .B1(new_n207), .B2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n252), .B1(new_n249), .B2(new_n259), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n285), .B1(new_n319), .B2(new_n288), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n273), .A2(new_n275), .A3(G223), .A4(new_n269), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G87), .ZN(new_n397));
  INV_X1    g0197(.A(G226), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n397), .C1(new_n276), .C2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n395), .B1(new_n278), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(new_n322), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(G169), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n375), .B1(new_n394), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n399), .A2(new_n278), .ZN(new_n406));
  INV_X1    g0206(.A(new_n395), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n407), .A3(new_n296), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(G200), .B2(new_n400), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n391), .A2(new_n409), .A3(new_n393), .ZN(new_n410));
  XNOR2_X1  g0210(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(KEYINPUT75), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n391), .A2(new_n409), .A3(new_n393), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n394), .A2(new_n403), .A3(new_n375), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n405), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n332), .A2(new_n374), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(G97), .B(G107), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT6), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G97), .ZN(new_n425));
  NOR3_X1   g0225(.A1(new_n423), .A2(new_n425), .A3(G107), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n429));
  OAI21_X1  g0229(.A(G107), .B1(new_n377), .B2(new_n378), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n255), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT76), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n248), .A2(G97), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n207), .A2(G33), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n252), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n436), .B2(new_n425), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n431), .A2(new_n432), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n426), .B1(new_n423), .B2(new_n422), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n439), .A2(new_n208), .B1(new_n203), .B2(new_n309), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n316), .B1(new_n386), .B2(new_n387), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n251), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n437), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT76), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(new_n269), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT4), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n448));
  NAND2_X1  g0248(.A1(G33), .A2(G283), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n447), .A2(new_n448), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n278), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n207), .A2(G45), .ZN(new_n453));
  NOR2_X1   g0253(.A1(KEYINPUT5), .A2(G41), .ZN(new_n454));
  INV_X1    g0254(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n453), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G274), .ZN(new_n458));
  INV_X1    g0258(.A(new_n217), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n283), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n281), .A2(G1), .ZN(new_n462));
  INV_X1    g0262(.A(new_n456), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(new_n454), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G257), .A3(new_n284), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n267), .B1(new_n452), .B2(new_n467), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n322), .B(new_n466), .C1(new_n278), .C2(new_n451), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n438), .A2(new_n444), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n452), .A2(new_n467), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n466), .B1(new_n451), .B2(new_n278), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G190), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n472), .A2(new_n474), .A3(new_n442), .A4(new_n443), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n284), .A2(G274), .A3(new_n462), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n284), .A2(G250), .A3(new_n453), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(G1698), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n273), .A2(new_n275), .A3(G238), .A4(new_n269), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G116), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n479), .B1(new_n278), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n322), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(KEYINPUT77), .C1(G169), .C2(new_n484), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT77), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n278), .ZN(new_n488));
  INV_X1    g0288(.A(new_n479), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n488), .A2(new_n322), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(G169), .B1(new_n488), .B2(new_n489), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n493), .A2(KEYINPUT78), .A3(new_n208), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT78), .B1(new_n493), .B2(new_n208), .ZN(new_n495));
  NOR3_X1   g0295(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n273), .A2(new_n275), .A3(new_n208), .A4(G68), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT19), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(new_n261), .B2(new_n425), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n251), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  XOR2_X1   g0302(.A(KEYINPUT15), .B(G87), .Z(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT69), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT69), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n311), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n305), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n504), .A2(new_n252), .A3(new_n506), .A4(new_n435), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n502), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n486), .A2(new_n492), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(new_n502), .A2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n488), .A2(new_n489), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  INV_X1    g0314(.A(new_n436), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n484), .A2(G190), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n512), .A2(new_n514), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G116), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n305), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n306), .A2(G116), .A3(new_n435), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n250), .A2(new_n217), .B1(G20), .B2(new_n520), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n449), .B(new_n208), .C1(G33), .C2(new_n425), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT20), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n523), .A2(KEYINPUT20), .A3(new_n524), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n521), .B(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g0328(.A(KEYINPUT5), .B(G41), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n462), .B1(new_n459), .B2(new_n283), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(G270), .B1(new_n460), .B2(new_n457), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n274), .A2(G33), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n272), .A2(KEYINPUT3), .ZN(new_n533));
  OAI21_X1  g0333(.A(G303), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n273), .A2(new_n275), .A3(G264), .A4(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(new_n269), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n278), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n531), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G200), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n528), .B(new_n540), .C1(new_n296), .C2(new_n539), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n527), .A2(new_n539), .A3(G169), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT21), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n531), .A2(new_n538), .A3(G179), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n527), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n527), .A2(new_n539), .A3(KEYINPUT21), .A4(G169), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n541), .A2(new_n544), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n476), .A2(new_n519), .A3(new_n548), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n273), .A2(new_n275), .A3(G250), .A4(new_n269), .ZN(new_n551));
  NAND2_X1  g0351(.A1(G33), .A2(G294), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g0353(.A1(new_n553), .A2(new_n278), .B1(new_n530), .B2(G264), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n461), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n267), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G179), .B2(new_n555), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n482), .A2(G20), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT23), .B1(new_n316), .B2(G20), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n316), .A2(KEYINPUT23), .A3(G20), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n273), .A2(new_n275), .A3(new_n208), .A4(G87), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT79), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n208), .A3(G87), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n318), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(G87), .ZN(new_n569));
  NOR3_X1   g0369(.A1(new_n569), .A2(KEYINPUT22), .A3(G20), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n268), .A2(KEYINPUT79), .A3(new_n570), .ZN(new_n571));
  AOI221_X4 g0371(.A(KEYINPUT80), .B1(new_n564), .B2(KEYINPUT22), .C1(new_n568), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT80), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n571), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n563), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT24), .ZN(new_n578));
  NOR3_X1   g0378(.A1(new_n318), .A2(new_n565), .A3(new_n567), .ZN(new_n579));
  AOI21_X1  g0379(.A(KEYINPUT79), .B1(new_n268), .B2(new_n570), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n575), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT80), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n573), .A3(new_n575), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT24), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n563), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n255), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n249), .A2(new_n316), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n588), .B(KEYINPUT25), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(G107), .B2(new_n515), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n558), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n585), .B1(new_n584), .B2(new_n563), .ZN(new_n594));
  INV_X1    g0394(.A(new_n563), .ZN(new_n595));
  AOI211_X1 g0395(.A(KEYINPUT24), .B(new_n595), .C1(new_n582), .C2(new_n583), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n251), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(G200), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n555), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(G190), .B2(new_n555), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n597), .A2(new_n590), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n592), .A2(new_n593), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n592), .B2(new_n601), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n421), .A2(new_n549), .A3(new_n604), .ZN(G372));
  AOI21_X1  g0405(.A(new_n344), .B1(new_n370), .B2(G169), .ZN(new_n606));
  INV_X1    g0406(.A(new_n345), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT74), .B1(new_n370), .B2(new_n322), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n342), .A2(new_n346), .A3(G179), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n372), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n329), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n373), .B(new_n418), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n419), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(new_n404), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n298), .A2(new_n299), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n294), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g0419(.A(new_n619), .B(KEYINPUT83), .Z(new_n620));
  OAI21_X1  g0420(.A(new_n432), .B1(new_n431), .B2(new_n437), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n442), .A2(KEYINPUT76), .A3(new_n443), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n471), .A2(G169), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n473), .A2(G179), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n621), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n442), .B(new_n443), .C1(new_n473), .C2(new_n598), .ZN(new_n626));
  INV_X1    g0426(.A(new_n474), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n518), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n625), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n557), .B1(new_n597), .B2(new_n590), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n630), .B(new_n601), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n513), .A2(KEYINPUT82), .A3(new_n267), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT82), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n484), .B2(G169), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n634), .A2(new_n636), .A3(new_n485), .A4(new_n510), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n518), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n442), .A2(new_n443), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n469), .B2(new_n468), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n638), .A2(new_n640), .A3(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n625), .A2(new_n518), .A3(new_n511), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(KEYINPUT26), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n633), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n421), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n620), .A2(new_n645), .ZN(G369));
  NAND2_X1  g0446(.A1(new_n356), .A2(new_n208), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n528), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n632), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n548), .B2(new_n654), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G330), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n652), .B1(new_n587), .B2(new_n591), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n604), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n592), .A2(new_n653), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n597), .A2(new_n590), .A3(new_n600), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT81), .B1(new_n663), .B2(new_n631), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n592), .A2(new_n601), .A3(new_n593), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n632), .A2(new_n653), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n631), .A2(new_n653), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n662), .A2(new_n669), .ZN(G399));
  INV_X1    g0470(.A(new_n211), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n496), .A2(new_n520), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G1), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n215), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n633), .A2(new_n637), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n638), .A2(new_n640), .ZN(new_n680));
  MUX2_X1   g0480(.A(new_n642), .B(new_n680), .S(KEYINPUT26), .Z(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n678), .B1(new_n682), .B2(new_n653), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n644), .A2(new_n653), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  NOR4_X1   g0486(.A1(new_n476), .A2(new_n519), .A3(new_n548), .A4(new_n652), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n664), .A2(new_n687), .A3(new_n665), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n484), .A2(new_n554), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n545), .A3(KEYINPUT30), .A4(new_n473), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n484), .A2(G179), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n471), .A2(new_n691), .A3(new_n539), .A4(new_n555), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n484), .A2(new_n554), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n531), .A2(new_n538), .A3(G179), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n471), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n690), .B(new_n692), .C1(new_n695), .C2(KEYINPUT30), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT31), .B1(new_n696), .B2(new_n652), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(KEYINPUT31), .A3(new_n652), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n686), .B1(new_n688), .B2(new_n700), .ZN(new_n701));
  NOR3_X1   g0501(.A1(new_n683), .A2(new_n685), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n677), .B1(new_n702), .B2(G1), .ZN(G364));
  INV_X1    g0503(.A(new_n657), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n355), .A2(G20), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n207), .B1(new_n705), .B2(G45), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n672), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(G330), .B2(new_n656), .ZN(new_n710));
  OAI21_X1  g0510(.A(G20), .B1(KEYINPUT85), .B2(G169), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(KEYINPUT85), .A2(G169), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n217), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n208), .A2(new_n322), .ZN(new_n716));
  NOR2_X1   g0516(.A1(G190), .A2(G200), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G311), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n318), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(G20), .A3(new_n322), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(G329), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n716), .A2(new_n296), .A3(G200), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT33), .B(G317), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n296), .A2(G200), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n322), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n725), .A2(new_n726), .B1(new_n729), .B2(G294), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n716), .A2(KEYINPUT86), .A3(new_n727), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT86), .B1(new_n716), .B2(new_n727), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n731), .B1(G322), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n716), .A2(G190), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR4_X1   g0538(.A1(new_n208), .A2(new_n598), .A3(G179), .A4(G190), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n738), .A2(G326), .B1(G283), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G303), .ZN(new_n741));
  NOR4_X1   g0541(.A1(new_n208), .A2(new_n296), .A3(new_n598), .A4(G179), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n736), .B(new_n740), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n569), .B1(new_n221), .B2(new_n724), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n722), .A2(G159), .ZN(new_n746));
  OAI22_X1  g0546(.A1(new_n746), .A2(KEYINPUT32), .B1(new_n202), .B2(new_n737), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n735), .A2(G58), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n268), .B1(new_n718), .B2(new_n203), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(KEYINPUT32), .B2(new_n746), .ZN(new_n751));
  AOI22_X1  g0551(.A1(new_n729), .A2(G97), .B1(new_n739), .B2(G107), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n748), .A2(new_n749), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n715), .B1(new_n744), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G13), .A2(G33), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n714), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n671), .A2(new_n318), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT84), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n761), .A2(G355), .B1(new_n520), .B2(new_n671), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n216), .A2(new_n281), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n671), .A2(new_n268), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n763), .B(new_n764), .C1(new_n243), .C2(new_n281), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n759), .B1(new_n762), .B2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n708), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n754), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n757), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n768), .B1(new_n656), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n710), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(G396));
  NAND3_X1  g0572(.A1(new_n324), .A2(new_n328), .A3(new_n652), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT91), .ZN(new_n774));
  INV_X1    g0574(.A(KEYINPUT91), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n324), .A2(new_n775), .A3(new_n328), .A4(new_n652), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n314), .A2(new_n652), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n331), .A2(new_n329), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT92), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n777), .A2(KEYINPUT92), .A3(new_n779), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n756), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n714), .A2(new_n755), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n739), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n788), .A2(new_n569), .B1(new_n719), .B2(new_n721), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT89), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT87), .B(G283), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n724), .A2(new_n791), .B1(new_n718), .B2(new_n520), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n792), .B(KEYINPUT88), .Z(new_n793));
  INV_X1    g0593(.A(G294), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n734), .A2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n738), .A2(G303), .B1(new_n742), .B2(G107), .ZN(new_n796));
  INV_X1    g0596(.A(new_n729), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n318), .C1(new_n425), .C2(new_n797), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n790), .A2(new_n793), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G137), .ZN(new_n800));
  INV_X1    g0600(.A(G150), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n800), .A2(new_n737), .B1(new_n724), .B2(new_n801), .ZN(new_n802));
  XOR2_X1   g0602(.A(new_n802), .B(KEYINPUT90), .Z(new_n803));
  INV_X1    g0603(.A(G143), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n803), .B1(new_n804), .B2(new_n734), .C1(new_n805), .C2(new_n718), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT34), .ZN(new_n807));
  INV_X1    g0607(.A(G132), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n268), .B1(new_n721), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n739), .A2(G68), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n810), .B1(new_n743), .B2(new_n202), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(G58), .C2(new_n729), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n799), .B1(new_n807), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n708), .B1(G77), .B2(new_n787), .C1(new_n813), .C2(new_n715), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n785), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n783), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT92), .B1(new_n777), .B2(new_n779), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n684), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n784), .A2(new_n644), .A3(new_n653), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n701), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n819), .A2(new_n820), .A3(new_n701), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n767), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n823), .B2(KEYINPUT93), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT93), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n822), .A2(new_n825), .A3(new_n767), .ZN(new_n826));
  AOI211_X1 g0626(.A(KEYINPUT94), .B(new_n815), .C1(new_n824), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT94), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n823), .A2(KEYINPUT93), .ZN(new_n829));
  INV_X1    g0629(.A(new_n821), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n829), .A2(new_n826), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n815), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n827), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G384));
  NOR2_X1   g0635(.A1(new_n705), .A2(new_n207), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT40), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT95), .B1(new_n372), .B2(new_n653), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT95), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n364), .A2(new_n839), .A3(new_n652), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n373), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n612), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n365), .A2(new_n373), .A3(new_n838), .A4(new_n840), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n843), .B(new_n844), .C1(new_n816), .C2(new_n817), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n625), .A2(new_n628), .ZN(new_n846));
  INV_X1    g0646(.A(new_n548), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n511), .A2(new_n518), .ZN(new_n848));
  NAND4_X1  g0648(.A1(new_n846), .A2(new_n847), .A3(new_n848), .A4(new_n653), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n602), .A2(new_n603), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT98), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n699), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n698), .ZN(new_n853));
  AOI211_X1 g0653(.A(KEYINPUT98), .B(KEYINPUT31), .C1(new_n696), .C2(new_n652), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT99), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n697), .B1(new_n851), .B2(new_n699), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n858), .A2(new_n854), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT99), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n688), .A3(new_n860), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n837), .B(new_n845), .C1(new_n857), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n650), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n394), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n394), .B1(new_n403), .B2(new_n866), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT97), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n869), .A2(new_n410), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n420), .A2(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n870), .A2(KEYINPUT37), .A3(new_n410), .A4(new_n869), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n865), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n867), .B1(new_n616), .B2(new_n418), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n869), .A2(KEYINPUT37), .A3(new_n410), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n876), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n863), .B1(new_n875), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n420), .A2(new_n868), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n871), .A2(new_n872), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n874), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n864), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n878), .A4(new_n879), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(KEYINPUT100), .A3(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n881), .B1(new_n876), .B2(new_n880), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n888), .ZN(new_n892));
  INV_X1    g0692(.A(new_n845), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n859), .A2(new_n688), .A3(new_n860), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n860), .B1(new_n859), .B2(new_n688), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI22_X1  g0696(.A1(new_n862), .A2(new_n890), .B1(new_n896), .B2(new_n837), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n857), .A2(new_n861), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n421), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n897), .A2(new_n899), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n900), .A2(new_n901), .A3(new_n686), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n421), .B1(new_n683), .B2(new_n685), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n620), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT39), .B1(new_n887), .B2(new_n888), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n891), .A2(new_n888), .A3(KEYINPUT39), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n612), .A2(new_n653), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n329), .A2(new_n652), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n820), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n844), .A2(new_n843), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(new_n892), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n650), .B1(new_n615), .B2(new_n404), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n911), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n905), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n836), .B1(new_n903), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n903), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n428), .A2(KEYINPUT35), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n922), .A2(G116), .A3(new_n218), .A4(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n924), .B(KEYINPUT36), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n215), .A2(new_n203), .A3(new_n382), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n221), .A2(G50), .ZN(new_n927));
  OAI211_X1 g0727(.A(G1), .B(new_n355), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n921), .A2(new_n925), .A3(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n512), .A2(new_n516), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n652), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n637), .A3(new_n518), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n637), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT42), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n639), .A2(new_n652), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n846), .A2(new_n937), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n640), .A2(new_n653), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OR3_X1    g0741(.A1(new_n667), .A2(KEYINPUT102), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT102), .B1(new_n667), .B2(new_n941), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n940), .B(KEYINPUT101), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n631), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n652), .B1(new_n946), .B2(new_n470), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n942), .A2(new_n936), .A3(new_n943), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n949), .A2(KEYINPUT103), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(KEYINPUT103), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n662), .A2(new_n945), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n954), .A2(KEYINPUT104), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(KEYINPUT104), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AND3_X1   g0757(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n957), .B1(new_n952), .B2(new_n953), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n935), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n952), .A2(new_n953), .ZN(new_n961));
  INV_X1    g0761(.A(new_n957), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n934), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n672), .B(KEYINPUT41), .Z(new_n966));
  INV_X1    g0766(.A(new_n702), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n659), .A2(new_n661), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n667), .B1(new_n968), .B2(new_n666), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n704), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n704), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n667), .A2(KEYINPUT45), .A3(new_n668), .A4(new_n940), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n669), .B2(new_n941), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n973), .A2(new_n975), .B1(new_n662), .B2(KEYINPUT105), .ZN(new_n976));
  INV_X1    g0776(.A(new_n662), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT105), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n940), .B1(new_n667), .B2(new_n668), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT44), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n976), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n979), .B1(new_n976), .B2(new_n981), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n972), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n966), .B1(new_n985), .B2(new_n702), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n960), .B(new_n965), .C1(new_n986), .C2(new_n707), .ZN(new_n987));
  INV_X1    g0787(.A(new_n764), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n758), .B1(new_n211), .B2(new_n507), .C1(new_n988), .C2(new_n238), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n989), .A2(new_n708), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n318), .B1(new_n991), .B2(new_n721), .C1(new_n788), .C2(new_n425), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT106), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n724), .A2(new_n794), .B1(new_n718), .B2(new_n791), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n797), .A2(new_n316), .B1(new_n737), .B2(new_n719), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n993), .B2(new_n992), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT46), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n743), .B2(new_n520), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n742), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(new_n741), .C2(new_n734), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n797), .A2(new_n221), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G143), .B2(new_n738), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n381), .B2(new_n743), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n788), .A2(new_n203), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n268), .B1(new_n721), .B2(new_n800), .C1(new_n718), .C2(new_n202), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G159), .C2(new_n725), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n801), .B2(new_n734), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n998), .A2(new_n1002), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n990), .B1(new_n769), .B2(new_n933), .C1(new_n1012), .C2(new_n715), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n987), .A2(new_n1013), .ZN(G387));
  NAND2_X1  g0814(.A1(new_n970), .A2(new_n971), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n764), .B1(new_n235), .B2(new_n281), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n761), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n674), .B2(new_n1017), .ZN(new_n1018));
  OR3_X1    g0818(.A1(new_n259), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT50), .B1(new_n259), .B2(G50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1019), .A2(new_n674), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1018), .A2(new_n1022), .B1(new_n316), .B2(new_n671), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n708), .B1(new_n1023), .B2(new_n759), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT108), .B(G150), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n268), .B1(new_n1025), .B2(new_n721), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n743), .A2(new_n203), .B1(new_n805), .B2(new_n737), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(G97), .C2(new_n739), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n724), .A2(new_n259), .B1(new_n718), .B2(new_n221), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT109), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n735), .A2(G50), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n312), .A2(new_n729), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1028), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n268), .B1(new_n722), .B2(G326), .ZN(new_n1034));
  INV_X1    g0834(.A(G322), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n737), .A2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n724), .A2(new_n719), .B1(new_n718), .B2(new_n741), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n735), .C2(G317), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT110), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(KEYINPUT48), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n797), .A2(new_n791), .B1(new_n743), .B2(new_n794), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1034), .B1(new_n520), .B2(new_n788), .C1(new_n1044), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1044), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1047), .A2(KEYINPUT49), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1033), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1024), .B1(new_n1049), .B2(new_n714), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n659), .A2(new_n661), .A3(new_n757), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1015), .A2(new_n707), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n972), .A2(new_n673), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n1015), .A2(new_n702), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(G393));
  NOR2_X1   g0855(.A1(new_n945), .A2(new_n769), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n734), .A2(new_n719), .B1(new_n991), .B2(new_n737), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n318), .B1(new_n721), .B2(new_n1035), .C1(new_n718), .C2(new_n794), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n788), .A2(new_n316), .B1(new_n741), .B2(new_n724), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n797), .A2(new_n520), .B1(new_n743), .B2(new_n791), .ZN(new_n1061));
  NOR4_X1   g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n734), .A2(new_n805), .B1(new_n801), .B2(new_n737), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  OAI221_X1 g0864(.A(new_n268), .B1(new_n721), .B2(new_n804), .C1(new_n718), .C2(new_n259), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n797), .A2(new_n203), .B1(new_n569), .B2(new_n788), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n743), .A2(new_n221), .B1(new_n202), .B2(new_n724), .ZN(new_n1067));
  NOR4_X1   g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n714), .B1(new_n1062), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n988), .A2(new_n246), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n758), .B1(new_n425), .B2(new_n211), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n708), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1056), .A2(new_n1072), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n983), .A2(new_n984), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1073), .B1(new_n1074), .B2(new_n707), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n972), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n985), .A2(new_n672), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1075), .B1(new_n1076), .B2(new_n1077), .ZN(G390));
  OAI21_X1  g0878(.A(new_n708), .B1(new_n787), .B2(new_n260), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT112), .Z(new_n1080));
  AOI21_X1  g0880(.A(new_n268), .B1(new_n742), .B2(G87), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT115), .Z(new_n1082));
  OAI221_X1 g0882(.A(new_n810), .B1(new_n425), .B2(new_n718), .C1(new_n794), .C2(new_n721), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G116), .B2(new_n735), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n797), .A2(new_n203), .B1(new_n724), .B2(new_n316), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G283), .B2(new_n738), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT54), .B(G143), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n797), .A2(new_n805), .B1(new_n718), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G137), .B2(new_n725), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT113), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n318), .B1(new_n722), .B2(G125), .ZN(new_n1092));
  INV_X1    g0892(.A(G128), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n737), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(G50), .B2(new_n739), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n735), .A2(G132), .ZN(new_n1096));
  XOR2_X1   g0896(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OR3_X1    g0898(.A1(new_n743), .A2(new_n1098), .A3(new_n1025), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1098), .B1(new_n743), .B2(new_n1025), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1095), .A2(new_n1096), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1087), .B1(new_n1091), .B2(new_n1101), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1102), .A2(KEYINPUT116), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n715), .B1(new_n1102), .B2(KEYINPUT116), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1080), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n908), .B2(new_n756), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n910), .B1(new_n914), .B2(new_n915), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n915), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n682), .A2(new_n784), .A3(new_n653), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1108), .B1(new_n1109), .B2(new_n913), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n883), .A2(new_n889), .A3(new_n909), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1107), .A2(new_n908), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(KEYINPUT111), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT111), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n898), .A2(new_n1115), .A3(G330), .A4(new_n893), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n701), .A2(new_n784), .A3(new_n915), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n1110), .B2(new_n1111), .C1(new_n1107), .C2(new_n908), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1106), .B1(new_n1121), .B2(new_n706), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT117), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n701), .A2(new_n784), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1108), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1114), .A2(new_n1116), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n914), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1119), .A2(new_n913), .A3(new_n1109), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n898), .A2(G330), .A3(new_n784), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1129), .B2(new_n1108), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n686), .B1(new_n857), .B2(new_n861), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n421), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n620), .A2(new_n904), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(new_n1121), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1121), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n672), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1123), .B1(new_n1138), .B2(new_n1140), .ZN(G378));
  NOR2_X1   g0941(.A1(new_n266), .A2(new_n650), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n300), .A2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n300), .B1(new_n266), .B2(new_n650), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1144), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n897), .B2(G330), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n845), .B1(new_n857), .B2(new_n861), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1153), .A2(KEYINPUT40), .A3(new_n883), .A4(new_n889), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n896), .A2(new_n837), .ZN(new_n1155));
  AND4_X1   g0955(.A1(G330), .A2(new_n1154), .A3(new_n1151), .A4(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n918), .B1(new_n1152), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(G330), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1151), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n897), .A2(G330), .A3(new_n1151), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n918), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1157), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1159), .A2(new_n755), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n708), .B1(new_n787), .B2(G50), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT118), .Z(new_n1167));
  NOR2_X1   g0967(.A1(new_n268), .A2(G41), .ZN(new_n1168));
  AOI211_X1 g0968(.A(G50), .B(new_n1168), .C1(new_n272), .C2(new_n280), .ZN(new_n1169));
  INV_X1    g0969(.A(G283), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1168), .B1(new_n1170), .B2(new_n721), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n1003), .C1(G107), .C2(new_n735), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n743), .A2(new_n203), .B1(new_n788), .B2(new_n381), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n425), .A2(new_n724), .B1(new_n737), .B2(new_n520), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(new_n507), .C2(new_n718), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1169), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n724), .A2(new_n808), .B1(new_n718), .B2(new_n800), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n735), .B2(G128), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G125), .A2(new_n738), .B1(new_n729), .B2(G150), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n743), .C2(new_n1088), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n739), .A2(G159), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n722), .C2(G124), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1178), .B1(new_n1177), .B2(new_n1176), .C1(new_n1183), .C2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1167), .B1(new_n1188), .B2(new_n714), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n1164), .A2(new_n707), .B1(new_n1165), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1130), .B1(new_n1126), .B2(new_n914), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1136), .B1(new_n1121), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1164), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1194), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n673), .B1(new_n1196), .B2(new_n1192), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT119), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(KEYINPUT119), .B(new_n673), .C1(new_n1196), .C2(new_n1192), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1190), .B1(new_n1199), .B2(new_n1200), .ZN(G375));
  INV_X1    g1001(.A(new_n966), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1127), .A2(new_n1135), .A3(new_n1131), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1137), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n915), .A2(new_n756), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT120), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n787), .A2(G68), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n520), .A2(new_n724), .B1(new_n737), .B2(new_n794), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(new_n1006), .C1(G97), .C2(new_n742), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n318), .B1(new_n721), .B2(new_n741), .C1(new_n718), .C2(new_n316), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n312), .B2(new_n729), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(new_n1170), .C2(new_n734), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT121), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n808), .A2(new_n737), .B1(new_n724), .B2(new_n1088), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G159), .B2(new_n742), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n735), .A2(G137), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n268), .B1(new_n718), .B2(new_n801), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G128), .B2(new_n722), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n729), .A2(G50), .B1(new_n739), .B2(G58), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1214), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n767), .B(new_n1207), .C1(new_n1223), .C2(new_n714), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1206), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1191), .B2(new_n706), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1204), .A2(new_n1227), .ZN(G381));
  OR2_X1    g1028(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1230));
  OR4_X1    g1030(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1231), .A2(G378), .A3(G387), .A4(G381), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .ZN(G407));
  NOR2_X1   g1033(.A1(new_n1140), .A2(new_n1138), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT117), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1122), .B(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n651), .A2(G213), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(new_n1238), .B(KEYINPUT123), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1229), .A2(new_n1237), .A3(new_n1230), .A4(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(G213), .A3(G407), .ZN(G409));
  AND3_X1   g1041(.A1(new_n987), .A2(new_n1013), .A3(G390), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n987), .B2(new_n1013), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT127), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(G393), .B(new_n771), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1245), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1247), .B(KEYINPUT127), .C1(new_n1242), .C2(new_n1243), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G378), .B(new_n1190), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1165), .A2(new_n1189), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n1193), .B2(new_n966), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT124), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1164), .A2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT124), .B1(new_n1157), .B2(new_n1163), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1254), .A2(new_n706), .A3(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1237), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1250), .A2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT125), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n827), .B2(new_n833), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n673), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1191), .A2(KEYINPUT60), .A3(new_n1135), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT60), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1203), .A2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n833), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n831), .A2(new_n828), .A3(new_n832), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1227), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1266), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1226), .B1(new_n834), .B2(KEYINPUT125), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1262), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1272), .A2(new_n1273), .A3(new_n1260), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1258), .A2(new_n1238), .A3(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1239), .B1(new_n1250), .B2(new_n1257), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1275), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(new_n1277), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n1276), .A2(new_n1277), .B1(new_n1278), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n651), .A2(G213), .A3(G2897), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1272), .A2(new_n1273), .A3(new_n1260), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1260), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1284), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1239), .A2(G2897), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1271), .A2(new_n1274), .A3(new_n1288), .ZN(new_n1289));
  AND3_X1   g1089(.A1(new_n1287), .A2(new_n1289), .A3(KEYINPUT126), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT126), .B1(new_n1287), .B2(new_n1289), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1282), .B1(new_n1292), .B2(new_n1278), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1249), .B1(new_n1281), .B2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1246), .A2(new_n1282), .A3(new_n1248), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT63), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1279), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1295), .B1(new_n1278), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT126), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1287), .A2(new_n1289), .A3(KEYINPUT126), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1258), .A2(new_n1238), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1296), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1276), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1298), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1294), .A2(new_n1307), .ZN(G405));
  NAND2_X1  g1108(.A1(new_n1249), .A2(new_n1279), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1246), .A2(new_n1248), .A3(new_n1275), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(G375), .B(G378), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1311), .B(new_n1312), .ZN(G402));
endmodule


