//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n811, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G228gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208));
  OR2_X1    g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(KEYINPUT81), .B(G155gat), .Z(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G162gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n211), .B1(new_n213), .B2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n208), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT80), .A3(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n209), .A2(new_n210), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n216), .A2(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT82), .B1(new_n214), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT81), .B(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n221), .A3(new_n208), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n222), .A2(new_n209), .A3(new_n210), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT80), .B1(new_n218), .B2(new_n219), .ZN(new_n230));
  INV_X1    g029(.A(new_n219), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n231), .A2(new_n217), .A3(new_n215), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n229), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n224), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  INV_X1    g036(.A(G204gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G197gat), .ZN(new_n239));
  INV_X1    g038(.A(G197gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G204gat), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(G211gat), .ZN(new_n243));
  OR2_X1    g042(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n242), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT76), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n239), .A2(new_n241), .ZN(new_n250));
  AND2_X1   g049(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n252));
  OAI21_X1  g051(.A(G211gat), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n254));
  NOR2_X1   g053(.A1(KEYINPUT74), .A2(KEYINPUT22), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n250), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT76), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT77), .ZN(new_n260));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n249), .A2(new_n259), .A3(new_n260), .A4(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n261), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n248), .B2(KEYINPUT76), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n260), .B1(new_n266), .B2(new_n259), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n237), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT3), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n236), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n267), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(new_n264), .A3(new_n263), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n228), .A2(new_n233), .A3(new_n269), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n274));
  AND2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n207), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n274), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n248), .A2(new_n262), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n264), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n280), .A2(KEYINPUT88), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n269), .B1(new_n280), .B2(KEYINPUT88), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n214), .A2(new_n223), .ZN(new_n284));
  OAI221_X1 g083(.A(new_n206), .B1(new_n272), .B2(new_n275), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n277), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n277), .B2(new_n285), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n205), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n277), .A2(new_n285), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n286), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n285), .A3(new_n287), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n204), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G15gat), .B(G43gat), .Z(new_n296));
  XNOR2_X1  g095(.A(G71gat), .B(G99gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(G227gat), .ZN(new_n299));
  INV_X1    g098(.A(G233gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(G169gat), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT23), .ZN(new_n304));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(KEYINPUT64), .ZN(new_n314));
  OR3_X1    g113(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n309), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n303), .A2(KEYINPUT65), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(G169gat), .B2(G176gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(KEYINPUT23), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n305), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n324), .A2(new_n327), .A3(new_n305), .ZN(new_n328));
  NAND2_X1  g127(.A1(G183gat), .A2(G190gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT24), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT67), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n313), .A3(new_n316), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n333));
  OR2_X1    g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n319), .B1(new_n308), .B2(new_n307), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n326), .A2(new_n328), .A3(new_n334), .A4(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n339), .A3(new_n312), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT28), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT27), .B(G183gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(new_n343), .A3(new_n312), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT26), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n321), .A2(new_n346), .A3(new_n323), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n348), .A2(new_n305), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n347), .A2(new_n349), .B1(G183gat), .B2(G190gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT68), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n345), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n347), .A2(new_n349), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n329), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT68), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n320), .A2(new_n336), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n357));
  INV_X1    g156(.A(G134gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G127gat), .ZN(new_n359));
  INV_X1    g158(.A(G127gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G134gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT1), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  INV_X1    g163(.A(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G113gat), .A2(G120gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n357), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(G113gat), .A2(G120gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(G113gat), .A2(G120gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G127gat), .B(G134gat), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT70), .A4(new_n362), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT69), .B1(new_n370), .B2(new_n371), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT69), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n366), .A2(new_n377), .A3(new_n367), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n376), .A2(new_n378), .A3(new_n362), .ZN(new_n379));
  INV_X1    g178(.A(new_n373), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n375), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n356), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n324), .A2(new_n327), .A3(new_n305), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n327), .B1(new_n324), .B2(new_n305), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n335), .B1(new_n332), .B2(new_n333), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT25), .B1(new_n309), .B2(new_n317), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n353), .A2(new_n351), .A3(new_n329), .ZN(new_n392));
  AND2_X1   g191(.A1(new_n341), .A2(new_n344), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n350), .A2(new_n351), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n390), .A2(new_n391), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n383), .A2(new_n385), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n302), .B1(new_n386), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n400));
  OAI21_X1  g199(.A(new_n298), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT32), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n398), .ZN(new_n405));
  AOI221_X4 g204(.A(new_n402), .B1(new_n400), .B2(new_n298), .C1(new_n405), .C2(new_n301), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n302), .A3(new_n398), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(KEYINPUT34), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n404), .A2(KEYINPUT73), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(KEYINPUT73), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n401), .A2(new_n403), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n411), .B1(new_n412), .B2(new_n406), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n295), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n265), .A2(new_n267), .ZN(new_n416));
  NAND2_X1  g215(.A1(G226gat), .A2(G233gat), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n396), .B2(new_n274), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n320), .A2(new_n336), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n352), .A2(new_n355), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n416), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n418), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT29), .B1(new_n420), .B2(new_n421), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n424), .B(new_n272), .C1(new_n425), .C2(new_n418), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n430), .A2(KEYINPUT30), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(KEYINPUT30), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n423), .A2(new_n426), .ZN(new_n434));
  INV_X1    g233(.A(new_n429), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI211_X1 g235(.A(KEYINPUT79), .B(new_n429), .C1(new_n423), .C2(new_n426), .ZN(new_n437));
  OAI22_X1  g236(.A1(new_n431), .A2(new_n432), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n440));
  NAND3_X1  g239(.A1(new_n224), .A2(new_n382), .A3(new_n235), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n375), .A2(new_n228), .A3(new_n381), .A4(new_n233), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G225gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n440), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n383), .A2(new_n284), .A3(new_n385), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT4), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n224), .A2(KEYINPUT3), .A3(new_n235), .ZN(new_n450));
  AND2_X1   g249(.A1(new_n273), .A2(new_n382), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT83), .B1(new_n442), .B2(KEYINPUT4), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n454), .B1(new_n447), .B2(KEYINPUT4), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n446), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n383), .A2(new_n457), .A3(new_n284), .A4(new_n385), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n442), .A2(KEYINPUT4), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n461));
  INV_X1    g260(.A(new_n440), .ZN(new_n462));
  AOI211_X1 g261(.A(new_n445), .B(new_n462), .C1(new_n450), .C2(new_n451), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT85), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n464), .A3(new_n459), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n456), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G1gat), .B(G29gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT0), .ZN(new_n469));
  XNOR2_X1  g268(.A(G57gat), .B(G85gat), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n469), .B(new_n470), .Z(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n474));
  NAND3_X1  g273(.A1(new_n456), .A2(new_n466), .A3(new_n471), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n474), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n467), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n439), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT35), .B1(new_n415), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n404), .A2(new_n407), .A3(new_n409), .ZN(new_n482));
  INV_X1    g281(.A(new_n409), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n412), .B2(new_n406), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n471), .B1(new_n456), .B2(new_n466), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n487), .A2(KEYINPUT89), .A3(new_n477), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT89), .B1(new_n487), .B2(new_n477), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n476), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n438), .A2(KEYINPUT35), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n486), .A2(new_n295), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n481), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT36), .B1(new_n482), .B2(new_n484), .ZN(new_n496));
  INV_X1    g295(.A(new_n414), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n496), .B1(new_n497), .B2(KEYINPUT36), .ZN(new_n498));
  INV_X1    g297(.A(new_n295), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n480), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n430), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n418), .B1(new_n396), .B2(new_n237), .ZN(new_n503));
  NOR3_X1   g302(.A1(new_n503), .A2(new_n422), .A3(new_n416), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n417), .B1(new_n356), .B2(new_n278), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n272), .B1(new_n505), .B2(new_n424), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n435), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n435), .A2(KEYINPUT37), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n396), .A2(new_n237), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n422), .B1(new_n511), .B2(new_n417), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n510), .B1(new_n512), .B2(new_n416), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n272), .B1(new_n419), .B2(new_n422), .ZN(new_n514));
  AOI21_X1  g313(.A(KEYINPUT38), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n502), .B1(new_n509), .B2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n478), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n487), .A2(KEYINPUT89), .A3(new_n477), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n516), .A2(new_n476), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n490), .A2(KEYINPUT90), .A3(new_n476), .A4(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n434), .A2(KEYINPUT37), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT38), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n450), .A2(new_n451), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n461), .A2(new_n529), .A3(new_n465), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT39), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n445), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(new_n471), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT39), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n535), .B1(new_n530), .B2(new_n445), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n528), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n445), .ZN(new_n538));
  INV_X1    g337(.A(new_n535), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT40), .A3(new_n471), .A4(new_n532), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n438), .A2(new_n537), .A3(new_n473), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n295), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT91), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n501), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n526), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n548), .B1(new_n520), .B2(new_n521), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n543), .B1(new_n549), .B2(new_n523), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n495), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  OR2_X1    g352(.A1(G43gat), .A2(G50gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(G43gat), .A2(G50gat), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT93), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n557), .A2(new_n553), .B1(G43gat), .B2(G50gat), .ZN(new_n558));
  XOR2_X1   g357(.A(KEYINPUT94), .B(G50gat), .Z(new_n559));
  OAI221_X1 g358(.A(new_n558), .B1(new_n557), .B2(new_n553), .C1(new_n559), .C2(G43gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(G29gat), .A2(G36gat), .ZN(new_n561));
  XOR2_X1   g360(.A(new_n561), .B(KEYINPUT92), .Z(new_n562));
  NOR2_X1   g361(.A1(G29gat), .A2(G36gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT14), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n556), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n565), .A2(new_n556), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT17), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G15gat), .B(G22gat), .ZN(new_n571));
  INV_X1    g370(.A(G1gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(KEYINPUT16), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n573), .B(new_n574), .C1(new_n572), .C2(new_n571), .ZN(new_n575));
  NAND2_X1  g374(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n575), .B(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT17), .B1(new_n566), .B2(new_n567), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n570), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n575), .B(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n568), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT18), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n580), .A2(new_n581), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n578), .B1(new_n566), .B2(new_n567), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n588), .A2(new_n583), .A3(KEYINPUT98), .ZN(new_n589));
  OR3_X1    g388(.A1(new_n568), .A2(new_n582), .A3(KEYINPUT98), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n581), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G197gat), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT11), .B(G169gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT12), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n584), .A3(new_n585), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n594), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n599), .B1(new_n594), .B2(new_n601), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n552), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT106), .ZN(new_n606));
  XOR2_X1   g405(.A(G99gat), .B(G106gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(G85gat), .A2(G92gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT7), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT102), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  INV_X1    g411(.A(G85gat), .ZN(new_n613));
  INV_X1    g412(.A(G92gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(KEYINPUT8), .A2(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n611), .B1(new_n610), .B2(new_n615), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n608), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n607), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n570), .A2(new_n579), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n568), .ZN(new_n625));
  NAND3_X1  g424(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G190gat), .B(G218gat), .Z(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n627), .A2(new_n628), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n632), .B1(new_n629), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  XOR2_X1   g436(.A(G57gat), .B(G64gat), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT9), .ZN(new_n639));
  XOR2_X1   g438(.A(G71gat), .B(G78gat), .Z(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n640), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n638), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n644), .A2(new_n645), .A3(new_n637), .A4(new_n638), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT101), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n651), .B1(new_n647), .B2(new_n648), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n582), .B1(new_n653), .B2(KEYINPUT21), .ZN(new_n654));
  OAI211_X1 g453(.A(G231gat), .B(G233gat), .C1(new_n653), .C2(KEYINPUT21), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT21), .ZN(new_n656));
  NAND2_X1  g455(.A1(G231gat), .A2(G233gat), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n656), .B(new_n657), .C1(new_n650), .C2(new_n652), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n360), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n360), .B1(new_n655), .B2(new_n658), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n654), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n661), .ZN(new_n663));
  INV_X1    g462(.A(new_n654), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(new_n664), .A3(new_n659), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G155gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G183gat), .B(G211gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n662), .A2(new_n665), .A3(new_n670), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n636), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n622), .B1(new_n650), .B2(new_n652), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n647), .A2(new_n648), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n622), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n649), .A2(KEYINPUT103), .A3(new_n619), .A4(new_n621), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n676), .A2(new_n677), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n653), .A2(KEYINPUT10), .A3(new_n624), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n682), .A2(KEYINPUT104), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT104), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n676), .A2(new_n680), .A3(new_n681), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n687), .ZN(new_n690));
  XNOR2_X1  g489(.A(G120gat), .B(G148gat), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n691), .B(new_n692), .Z(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n687), .B1(new_n682), .B2(new_n683), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n695), .B1(new_n689), .B2(new_n687), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n693), .B(KEYINPUT105), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI22_X1  g497(.A1(new_n688), .A2(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n606), .B1(new_n675), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n699), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n674), .A2(KEYINPUT106), .A3(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n605), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n479), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(new_n572), .ZN(G1324gat));
  NAND3_X1  g505(.A1(new_n605), .A2(new_n438), .A3(new_n703), .ZN(new_n707));
  AND2_X1   g506(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n707), .A2(G8gat), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT42), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(KEYINPUT42), .B2(new_n710), .ZN(G1325gat));
  OAI21_X1  g512(.A(G15gat), .B1(new_n704), .B2(new_n498), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n485), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n704), .B2(new_n715), .ZN(G1326gat));
  OAI21_X1  g515(.A(KEYINPUT107), .B1(new_n704), .B2(new_n295), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n605), .A2(new_n718), .A3(new_n499), .A4(new_n703), .ZN(new_n719));
  XNOR2_X1  g518(.A(KEYINPUT43), .B(G22gat), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n717), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n717), .B2(new_n719), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(G1327gat));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  INV_X1    g523(.A(new_n636), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n552), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n479), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n295), .B1(new_n479), .B2(new_n439), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n410), .A2(new_n413), .A3(KEYINPUT36), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n485), .B2(KEYINPUT36), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n550), .B2(KEYINPUT91), .ZN(new_n732));
  AOI211_X1 g531(.A(new_n546), .B(new_n543), .C1(new_n523), .C2(new_n549), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n494), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(KEYINPUT44), .A3(new_n636), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n672), .A2(new_n673), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(KEYINPUT110), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n699), .B(KEYINPUT111), .Z(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(new_n604), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n726), .A2(new_n727), .A3(new_n735), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G29gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n736), .A2(new_n725), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n701), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n604), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n479), .A2(G29gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n747), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n743), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT112), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n743), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1328gat));
  AND2_X1   g556(.A1(new_n726), .A2(new_n735), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n438), .A3(new_n741), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G36gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n734), .A2(new_n748), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n745), .B(KEYINPUT108), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n439), .A2(G36gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT113), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n768), .A3(new_n764), .ZN(new_n769));
  AND3_X1   g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n760), .B1(new_n770), .B2(new_n771), .ZN(G1329gat));
  NAND4_X1  g571(.A1(new_n726), .A2(new_n730), .A3(new_n735), .A4(new_n741), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n485), .A2(G43gat), .ZN(new_n774));
  AOI22_X1  g573(.A1(new_n773), .A2(G43gat), .B1(new_n763), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g575(.A1(new_n726), .A2(new_n499), .A3(new_n735), .A4(new_n741), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n777), .A2(new_n778), .A3(new_n559), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n295), .A2(new_n559), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n734), .A2(new_n747), .A3(new_n748), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT48), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n777), .A2(new_n559), .B1(new_n778), .B2(new_n784), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n781), .A2(new_n787), .ZN(new_n789));
  OAI21_X1  g588(.A(KEYINPUT48), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n791), .ZN(G1331gat));
  NOR4_X1   g591(.A1(new_n552), .A2(new_n748), .A3(new_n675), .A4(new_n739), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n727), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g594(.A(new_n438), .B(KEYINPUT117), .Z(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT49), .B(G64gat), .Z(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(G1333gat));
  NAND2_X1  g600(.A1(new_n793), .A2(new_n730), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G71gat), .ZN(new_n803));
  INV_X1    g602(.A(G71gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n793), .A2(new_n804), .A3(new_n486), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n803), .A2(KEYINPUT50), .A3(new_n805), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(G1334gat));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n499), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g611(.A1(new_n736), .A2(new_n748), .A3(new_n701), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n758), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G85gat), .B1(new_n814), .B2(new_n479), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n734), .A2(new_n604), .A3(new_n744), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n734), .A2(KEYINPUT51), .A3(new_n604), .A4(new_n744), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n820), .A2(new_n613), .A3(new_n727), .A4(new_n699), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n821), .ZN(G1336gat));
  NAND4_X1  g621(.A1(new_n726), .A2(new_n735), .A3(new_n797), .A4(new_n813), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G92gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n740), .A2(new_n797), .A3(new_n614), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n726), .A2(new_n438), .A3(new_n735), .A4(new_n813), .ZN(new_n830));
  AOI22_X1  g629(.A1(G92gat), .A2(new_n830), .B1(new_n820), .B2(new_n826), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n829), .B1(new_n831), .B2(new_n828), .ZN(G1337gat));
  OAI21_X1  g631(.A(G99gat), .B1(new_n814), .B2(new_n498), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n485), .A2(G99gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n820), .A2(new_n699), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1338gat));
  NAND4_X1  g635(.A1(new_n726), .A2(new_n499), .A3(new_n735), .A4(new_n813), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(G106gat), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n739), .A2(G106gat), .A3(new_n295), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n545), .A2(new_n546), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n551), .A3(new_n731), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n748), .B1(new_n841), .B2(new_n494), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n842), .B2(new_n744), .ZN(new_n843));
  INV_X1    g642(.A(new_n819), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n846));
  NOR2_X1   g645(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n847));
  XNOR2_X1  g646(.A(new_n847), .B(KEYINPUT119), .ZN(new_n848));
  AND4_X1   g647(.A1(new_n838), .A2(new_n845), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(new_n846), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n820), .B2(new_n839), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n848), .B1(new_n851), .B2(new_n838), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n849), .A2(new_n852), .ZN(G1339gat));
  NAND3_X1  g652(.A1(new_n674), .A2(new_n604), .A3(new_n701), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT120), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT120), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n674), .A2(new_n856), .A3(new_n604), .A4(new_n701), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n684), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n682), .A2(new_n683), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT104), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n687), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n694), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n693), .B1(new_n695), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT54), .B1(new_n860), .B2(new_n686), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n688), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n604), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n860), .A2(new_n866), .A3(new_n686), .ZN(new_n873));
  INV_X1    g672(.A(new_n693), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n868), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n863), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n872), .B1(new_n877), .B2(KEYINPUT55), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n868), .B1(new_n859), .B2(new_n862), .ZN(new_n879));
  NOR4_X1   g678(.A1(new_n879), .A2(KEYINPUT121), .A3(new_n870), .A4(new_n875), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n865), .B(new_n871), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n592), .B1(new_n589), .B2(new_n590), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n580), .A2(new_n583), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(G229gat), .A3(G233gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n601), .A2(new_n593), .A3(new_n587), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n888), .A2(new_n598), .B1(new_n889), .B2(new_n599), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n699), .A2(new_n890), .A3(KEYINPUT123), .ZN(new_n891));
  AOI21_X1  g690(.A(KEYINPUT123), .B1(new_n699), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n881), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n725), .ZN(new_n895));
  OAI211_X1 g694(.A(KEYINPUT55), .B(new_n867), .C1(new_n688), .C2(new_n868), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT121), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n863), .A2(new_n876), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n898), .A2(new_n872), .A3(KEYINPUT55), .A4(new_n867), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n897), .A2(new_n899), .B1(new_n863), .B2(new_n864), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n869), .A2(new_n870), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n636), .A3(new_n901), .A4(new_n890), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n858), .B1(new_n903), .B2(new_n737), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n904), .A2(new_n479), .A3(new_n415), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(new_n796), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n748), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n796), .A2(new_n727), .ZN(new_n908));
  NOR4_X1   g707(.A1(new_n904), .A2(new_n499), .A3(new_n485), .A4(new_n908), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n604), .A2(new_n364), .ZN(new_n910));
  AOI22_X1  g709(.A1(new_n907), .A2(new_n364), .B1(new_n909), .B2(new_n910), .ZN(G1340gat));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n699), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n739), .A2(new_n365), .ZN(new_n913));
  AOI22_X1  g712(.A1(new_n912), .A2(new_n365), .B1(new_n909), .B2(new_n913), .ZN(G1341gat));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n360), .A3(new_n736), .ZN(new_n915));
  INV_X1    g714(.A(new_n909), .ZN(new_n916));
  OAI21_X1  g715(.A(G127gat), .B1(new_n916), .B2(new_n737), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1342gat));
  NAND4_X1  g717(.A1(new_n905), .A2(new_n358), .A3(new_n439), .A4(new_n636), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT56), .ZN(new_n920));
  OAI21_X1  g719(.A(G134gat), .B1(new_n916), .B2(new_n725), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(KEYINPUT56), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(G1343gat));
  AND2_X1   g722(.A1(new_n699), .A2(new_n890), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(new_n900), .B2(new_n871), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n902), .B1(new_n925), .B2(new_n636), .ZN(new_n926));
  INV_X1    g725(.A(new_n736), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n858), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(KEYINPUT57), .B1(new_n928), .B2(new_n295), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT57), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n738), .B1(new_n895), .B2(new_n902), .ZN(new_n931));
  OAI211_X1 g730(.A(new_n930), .B(new_n499), .C1(new_n931), .C2(new_n858), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n908), .A2(new_n730), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n929), .A2(new_n932), .A3(new_n748), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(G141gat), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n904), .A2(new_n479), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n730), .A2(new_n295), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n604), .A2(G141gat), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n936), .A2(new_n796), .A3(new_n937), .A4(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT58), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n935), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1344gat));
  NAND2_X1  g743(.A1(new_n936), .A2(new_n937), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n945), .A2(new_n797), .ZN(new_n946));
  INV_X1    g745(.A(G148gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n699), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n701), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G148gat), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT57), .B1(new_n904), .B2(new_n295), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n926), .A2(new_n927), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n700), .A2(new_n604), .A3(new_n702), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n930), .B(new_n499), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n954), .A2(new_n957), .A3(new_n699), .A4(new_n933), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n951), .B1(new_n958), .B2(G148gat), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n948), .B1(new_n953), .B2(new_n959), .ZN(G1345gat));
  NAND3_X1  g759(.A1(new_n946), .A2(new_n225), .A3(new_n736), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n212), .B1(new_n949), .B2(new_n737), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1346gat));
  OAI21_X1  g762(.A(G162gat), .B1(new_n949), .B2(new_n725), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n439), .A2(new_n226), .A3(new_n636), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n945), .B2(new_n965), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n904), .A2(new_n727), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n796), .A2(new_n415), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT124), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(G169gat), .B1(new_n970), .B2(new_n748), .ZN(new_n971));
  INV_X1    g770(.A(new_n902), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n636), .B1(new_n881), .B2(new_n893), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n737), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n974), .A2(new_n857), .A3(new_n855), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n727), .A2(new_n439), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n977), .A2(new_n485), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n295), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n748), .A2(G169gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n971), .B1(new_n980), .B2(new_n981), .ZN(G1348gat));
  INV_X1    g781(.A(G176gat), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n970), .A2(new_n983), .A3(new_n699), .ZN(new_n984));
  OAI21_X1  g783(.A(G176gat), .B1(new_n979), .B2(new_n739), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1349gat));
  OAI21_X1  g785(.A(G183gat), .B1(new_n979), .B2(new_n737), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n967), .A2(new_n342), .A3(new_n736), .A4(new_n969), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(KEYINPUT60), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT60), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n987), .A2(new_n988), .A3(KEYINPUT125), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n990), .A2(new_n992), .ZN(G1350gat));
  NAND3_X1  g792(.A1(new_n970), .A2(new_n312), .A3(new_n636), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n636), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n995), .B1(new_n996), .B2(G190gat), .ZN(new_n997));
  AOI211_X1 g796(.A(KEYINPUT61), .B(new_n312), .C1(new_n980), .C2(new_n636), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G1351gat));
  NOR3_X1   g798(.A1(new_n796), .A2(new_n730), .A3(new_n295), .ZN(new_n1000));
  AND2_X1   g799(.A1(new_n967), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n748), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n954), .A2(new_n957), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n977), .A2(new_n730), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n604), .A2(new_n240), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1002), .B1(new_n1006), .B2(new_n1007), .ZN(G1352gat));
  NAND4_X1  g807(.A1(new_n967), .A2(new_n238), .A3(new_n699), .A4(new_n1000), .ZN(new_n1009));
  OR2_X1    g808(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1011));
  NOR3_X1   g810(.A1(new_n1003), .A2(new_n739), .A3(new_n1005), .ZN(new_n1012));
  OAI211_X1 g811(.A(new_n1010), .B(new_n1011), .C1(new_n1012), .C2(new_n238), .ZN(G1353gat));
  NAND3_X1  g812(.A1(new_n1001), .A2(new_n243), .A3(new_n736), .ZN(new_n1014));
  NAND4_X1  g813(.A1(new_n954), .A2(new_n957), .A3(new_n736), .A4(new_n1004), .ZN(new_n1015));
  AND3_X1   g814(.A1(new_n1015), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1016));
  AOI21_X1  g815(.A(KEYINPUT63), .B1(new_n1015), .B2(G211gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(G1354gat));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1019));
  NAND4_X1  g818(.A1(new_n954), .A2(new_n957), .A3(new_n1019), .A4(new_n1004), .ZN(new_n1020));
  AOI21_X1  g819(.A(new_n725), .B1(new_n244), .B2(new_n245), .ZN(new_n1021));
  AND2_X1   g820(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g821(.A(KEYINPUT127), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1023));
  NAND4_X1  g822(.A1(new_n975), .A2(new_n479), .A3(new_n636), .A4(new_n1000), .ZN(new_n1024));
  INV_X1    g823(.A(G218gat), .ZN(new_n1025));
  NAND3_X1  g824(.A1(new_n1024), .A2(KEYINPUT126), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1027));
  INV_X1    g826(.A(KEYINPUT126), .ZN(new_n1028));
  NAND2_X1  g827(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g828(.A1(new_n1022), .A2(new_n1023), .B1(new_n1026), .B2(new_n1029), .ZN(G1355gat));
endmodule


