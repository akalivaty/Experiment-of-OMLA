//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT64), .B(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G107), .A2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n208), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT2), .B(G226), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G264), .B(G270), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G58), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(KEYINPUT72), .ZN(new_n243));
  INV_X1    g0043(.A(KEYINPUT3), .ZN(new_n244));
  INV_X1    g0044(.A(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  OAI221_X1 g0053(.A(new_n250), .B1(new_n251), .B2(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n245), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n260));
  NOR3_X1   g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n256), .A2(new_n260), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT65), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT65), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n256), .A2(new_n264), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n261), .B1(new_n266), .B2(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n258), .A2(new_n267), .A3(KEYINPUT66), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G200), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n273), .A2(new_n214), .ZN(new_n274));
  NOR2_X1   g0074(.A1(G58), .A2(G68), .ZN(new_n275));
  INV_X1    g0075(.A(G50), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n206), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XOR2_X1   g0077(.A(new_n277), .B(KEYINPUT67), .Z(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT8), .B(G58), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n245), .A2(G20), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G20), .A2(G33), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n280), .A2(new_n281), .B1(G150), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n274), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n205), .A2(G20), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n273), .A2(new_n214), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n287), .A2(G50), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G50), .B2(new_n288), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n272), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n270), .A2(new_n271), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G190), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  OR4_X1    g0102(.A1(new_n243), .A2(new_n298), .A3(new_n299), .A4(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G179), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n300), .A2(KEYINPUT69), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT69), .B1(new_n300), .B2(new_n304), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n295), .B1(G169), .B2(new_n300), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n243), .A2(new_n299), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n243), .A2(new_n299), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n309), .B(new_n310), .C1(new_n298), .C2(new_n302), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT74), .ZN(new_n313));
  INV_X1    g0113(.A(new_n265), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n264), .B1(new_n256), .B2(new_n260), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n263), .A2(KEYINPUT74), .A3(new_n265), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(G238), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n261), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n248), .A2(G232), .A3(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n248), .A2(G226), .A3(new_n249), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT73), .A4(new_n323), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n256), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n320), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G238), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n266), .B2(new_n313), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n261), .B1(new_n331), .B2(new_n317), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n326), .A2(new_n327), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n257), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n332), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n329), .A2(new_n336), .A3(G190), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n289), .A2(new_n218), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n282), .A2(G50), .B1(G20), .B2(new_n218), .ZN(new_n340));
  INV_X1    g0140(.A(new_n281), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n251), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n287), .A2(G68), .A3(new_n291), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n339), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT11), .B1(new_n342), .B2(new_n290), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n329), .B2(new_n336), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT75), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n350), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT75), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n352), .A2(new_n353), .A3(new_n337), .A4(new_n347), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n347), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n329), .A2(new_n336), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n358), .A3(G169), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n329), .A2(new_n336), .A3(G179), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n358), .B1(new_n357), .B2(G169), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n356), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G87), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n245), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(KEYINPUT76), .A2(G33), .ZN(new_n367));
  NOR2_X1   g0167(.A1(KEYINPUT76), .A2(G33), .ZN(new_n368));
  OAI21_X1  g0168(.A(KEYINPUT3), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n249), .B1(new_n369), .B2(new_n246), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n366), .B1(new_n370), .B2(G226), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT76), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n245), .ZN(new_n373));
  NAND2_X1  g0173(.A1(KEYINPUT76), .A2(G33), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n244), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  OAI211_X1 g0176(.A(G223), .B(new_n249), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT78), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G1698), .B1(new_n369), .B2(new_n246), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n380), .A2(KEYINPUT78), .A3(G223), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n371), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n257), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n256), .A2(G232), .A3(new_n260), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT79), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n256), .A2(KEYINPUT79), .A3(G232), .A4(new_n260), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n319), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n383), .A2(new_n384), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n390), .B1(new_n382), .B2(new_n257), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n392), .B1(G200), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT80), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n287), .A2(new_n280), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n274), .A2(new_n288), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n397), .B1(new_n288), .B2(new_n280), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n373), .A2(new_n374), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n376), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n399), .B1(new_n401), .B2(new_n206), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n369), .A2(new_n399), .A3(new_n206), .A4(new_n246), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G68), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT77), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n369), .A2(new_n246), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT7), .B1(new_n406), .B2(G20), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G68), .A4(new_n403), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(G58), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n218), .ZN(new_n412));
  OAI21_X1  g0212(.A(G20), .B1(new_n412), .B2(new_n275), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n282), .A2(G159), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n410), .A2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n415), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n367), .A2(new_n368), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n244), .ZN(new_n421));
  AOI21_X1  g0221(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n422), .A2(KEYINPUT7), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n246), .A2(new_n422), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n421), .A2(new_n423), .B1(new_n399), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n419), .B1(new_n425), .B2(new_n218), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n274), .B1(new_n426), .B2(new_n416), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n398), .B1(new_n418), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n394), .A2(new_n395), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n395), .B1(new_n394), .B2(new_n428), .ZN(new_n430));
  OAI21_X1  g0230(.A(KEYINPUT17), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT18), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n393), .A2(G179), .ZN(new_n433));
  INV_X1    g0233(.A(G169), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n393), .ZN(new_n435));
  INV_X1    g0235(.A(new_n398), .ZN(new_n436));
  INV_X1    g0236(.A(new_n417), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n405), .B2(new_n409), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n423), .B1(KEYINPUT3), .B2(new_n400), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n424), .A2(new_n399), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n415), .B1(new_n441), .B2(G68), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n290), .B1(new_n442), .B2(KEYINPUT16), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n436), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n432), .B1(new_n435), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n393), .A2(new_n434), .ZN(new_n446));
  AOI211_X1 g0246(.A(new_n304), .B(new_n390), .C1(new_n382), .C2(new_n257), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n444), .B(new_n432), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(KEYINPUT17), .B1(new_n394), .B2(new_n428), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n431), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n261), .B1(new_n266), .B2(G244), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n455));
  INV_X1    g0255(.A(G107), .ZN(new_n456));
  OAI221_X1 g0256(.A(new_n455), .B1(new_n456), .B2(new_n248), .C1(new_n252), .C2(new_n217), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n454), .B1(new_n458), .B2(new_n256), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT70), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(KEYINPUT70), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n434), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n287), .A2(G77), .A3(new_n291), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(G77), .B2(new_n288), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n280), .A2(new_n282), .B1(G20), .B2(G77), .ZN(new_n465));
  XOR2_X1   g0265(.A(KEYINPUT15), .B(G87), .Z(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n281), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n274), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(new_n469), .B(KEYINPUT71), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT70), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n459), .B(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n462), .B(new_n470), .C1(new_n472), .C2(G179), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n460), .A2(new_n461), .A3(G200), .ZN(new_n474));
  INV_X1    g0274(.A(new_n470), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n474), .B(new_n475), .C1(new_n384), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NOR4_X1   g0277(.A1(new_n312), .A2(new_n364), .A3(new_n453), .A4(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT91), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n288), .A2(G116), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n397), .B1(new_n205), .B2(G33), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n481), .B1(new_n482), .B2(G116), .ZN(new_n483));
  INV_X1    g0283(.A(G116), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n273), .A2(new_n214), .B1(G20), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT86), .ZN(new_n486));
  OR2_X1    g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  INV_X1    g0288(.A(G97), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n488), .B(new_n206), .C1(G33), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT87), .ZN(new_n491));
  AOI21_X1  g0291(.A(G20), .B1(new_n245), .B2(G97), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT87), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n493), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n485), .A2(new_n486), .ZN(new_n496));
  AND4_X1   g0296(.A1(KEYINPUT20), .A2(new_n487), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n491), .A2(new_n494), .B1(new_n486), .B2(new_n485), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT20), .B1(new_n498), .B2(new_n487), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n483), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n249), .A2(G257), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n401), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n248), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G303), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n406), .A2(G264), .A3(G1698), .ZN(new_n507));
  INV_X1    g0307(.A(new_n503), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n406), .A2(KEYINPUT85), .A3(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n257), .ZN(new_n511));
  XNOR2_X1  g0311(.A(KEYINPUT5), .B(G41), .ZN(new_n512));
  INV_X1    g0312(.A(G45), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G1), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n512), .A2(new_n256), .A3(G274), .A4(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n514), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(new_n256), .ZN(new_n517));
  INV_X1    g0317(.A(G270), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n511), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(KEYINPUT21), .A3(G169), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n519), .B1(new_n510), .B2(new_n257), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G179), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n501), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT85), .B1(new_n406), .B2(new_n508), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n502), .B(new_n503), .C1(new_n369), .C2(new_n246), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI22_X1  g0328(.A1(new_n370), .A2(G264), .B1(G303), .B2(new_n505), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n256), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n500), .B(G169), .C1(new_n530), .C2(new_n519), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT88), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT88), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n521), .A2(new_n534), .A3(G169), .A4(new_n500), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT21), .B1(new_n531), .B2(KEYINPUT88), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(KEYINPUT89), .A3(new_n535), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n525), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n521), .A2(G200), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n523), .A2(G190), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(new_n501), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT90), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n542), .A2(KEYINPUT90), .A3(new_n501), .A4(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n480), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n525), .ZN(new_n550));
  AND4_X1   g0350(.A1(KEYINPUT89), .A2(new_n532), .A3(new_n533), .A4(new_n535), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT89), .B1(new_n539), .B2(new_n535), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n548), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n370), .A2(G257), .B1(G294), .B2(new_n400), .ZN(new_n556));
  INV_X1    g0356(.A(G250), .ZN(new_n557));
  INV_X1    g0357(.A(new_n380), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n257), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n257), .B1(new_n514), .B2(new_n512), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G264), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n560), .A2(new_n304), .A3(new_n515), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n515), .ZN(new_n564));
  INV_X1    g0364(.A(new_n562), .ZN(new_n565));
  AOI211_X1 g0365(.A(new_n564), .B(new_n565), .C1(new_n559), .C2(new_n257), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n434), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  OR4_X1    g0369(.A1(KEYINPUT22), .A2(new_n505), .A3(G20), .A4(new_n365), .ZN(new_n570));
  AOI21_X1  g0370(.A(G20), .B1(new_n369), .B2(new_n246), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(KEYINPUT92), .A3(G87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT22), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT92), .B1(new_n571), .B2(G87), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n420), .A2(new_n484), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n206), .B2(G107), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n456), .A2(KEYINPUT23), .A3(G20), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n576), .A2(new_n206), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n569), .B1(new_n575), .B2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n575), .A2(new_n569), .A3(new_n580), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n274), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT25), .B1(new_n289), .B2(new_n456), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n289), .A2(KEYINPUT25), .A3(new_n456), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n482), .A2(G107), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n563), .B(new_n568), .C1(new_n584), .C2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n580), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n406), .A2(new_n206), .A3(G87), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT92), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(KEYINPUT22), .A3(new_n572), .ZN(new_n595));
  AOI211_X1 g0395(.A(KEYINPUT24), .B(new_n591), .C1(new_n595), .C2(new_n570), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n290), .B1(new_n596), .B2(new_n581), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n560), .A2(new_n384), .A3(new_n515), .A4(new_n562), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n598), .B1(new_n566), .B2(G200), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n597), .A2(new_n599), .A3(new_n588), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n590), .A2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n489), .A2(new_n456), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(new_n202), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n456), .A2(KEYINPUT6), .A3(G97), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(G20), .B1(G77), .B2(new_n282), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n607), .B1(new_n425), .B2(new_n456), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n290), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n288), .A2(G97), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n291), .B1(G1), .B2(new_n245), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n489), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n564), .B1(G257), .B2(new_n561), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n488), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT4), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n406), .A2(G244), .A3(new_n249), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n304), .B(new_n616), .C1(new_n622), .C2(new_n256), .ZN(new_n623));
  INV_X1    g0423(.A(new_n616), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n620), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n625), .A2(new_n488), .A3(new_n617), .A4(new_n618), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n257), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n615), .B(new_n623), .C1(new_n627), .C2(G169), .ZN(new_n628));
  OAI211_X1 g0428(.A(G190), .B(new_n616), .C1(new_n622), .C2(new_n256), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n613), .B1(new_n608), .B2(new_n290), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n629), .B(new_n630), .C1(new_n627), .C2(new_n349), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT81), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n628), .A2(new_n631), .A3(KEYINPUT81), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n256), .B(G250), .C1(G1), .C2(new_n513), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n256), .A2(G274), .A3(new_n514), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT82), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT82), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n637), .A2(new_n641), .A3(new_n638), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n576), .B1(new_n380), .B2(G238), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n406), .A2(G244), .A3(G1698), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n256), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(G200), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n466), .A2(new_n288), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n612), .A2(new_n365), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n406), .A2(new_n206), .A3(G68), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT19), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n652), .B1(new_n341), .B2(new_n489), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n206), .B1(new_n323), .B2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n202), .A2(new_n365), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT83), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n654), .A2(KEYINPUT83), .A3(new_n655), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n651), .B(new_n653), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  AOI211_X1 g0458(.A(new_n649), .B(new_n650), .C1(new_n658), .C2(new_n290), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n645), .A2(new_n646), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n257), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n661), .A2(new_n643), .A3(G190), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n648), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n434), .B1(new_n644), .B2(new_n647), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n643), .A3(new_n304), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n290), .ZN(new_n666));
  INV_X1    g0466(.A(new_n649), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n482), .A2(new_n466), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n664), .A2(new_n665), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT84), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n663), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n663), .B2(new_n670), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n636), .A2(new_n674), .ZN(new_n675));
  NOR4_X1   g0475(.A1(new_n479), .A2(new_n555), .A3(new_n601), .A4(new_n675), .ZN(G372));
  INV_X1    g0476(.A(new_n450), .ZN(new_n677));
  INV_X1    g0477(.A(new_n355), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n363), .B1(new_n678), .B2(new_n473), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n431), .A2(new_n452), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n677), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n303), .A2(new_n311), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n307), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n660), .A2(new_n257), .B1(new_n640), .B2(new_n642), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n649), .B1(new_n658), .B2(new_n290), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n304), .A2(new_n685), .B1(new_n686), .B2(new_n668), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n661), .A2(new_n643), .ZN(new_n688));
  AOI21_X1  g0488(.A(KEYINPUT93), .B1(new_n688), .B2(new_n434), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n685), .A2(new_n690), .A3(G169), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n687), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n664), .A2(new_n690), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n688), .A2(KEYINPUT93), .A3(new_n434), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n694), .B1(new_n697), .B2(new_n687), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n685), .A2(new_n349), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n666), .B(new_n667), .C1(new_n365), .C2(new_n612), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT94), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT94), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n648), .A2(new_n659), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n662), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n628), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(new_n707), .A4(new_n692), .ZN(new_n708));
  NOR3_X1   g0508(.A1(new_n672), .A2(new_n673), .A3(new_n628), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n699), .B(new_n708), .C1(new_n709), .C2(new_n707), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n590), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n628), .A2(new_n631), .ZN(new_n713));
  AND4_X1   g0513(.A1(new_n600), .A2(new_n713), .A3(new_n705), .A4(new_n692), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n684), .B1(new_n479), .B2(new_n717), .ZN(G369));
  NAND3_X1  g0518(.A1(new_n541), .A2(new_n480), .A3(new_n548), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n553), .A2(KEYINPUT91), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT27), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT27), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n722), .A2(G213), .A3(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(G343), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n719), .A2(new_n720), .B1(new_n500), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n726), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n541), .A2(new_n501), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n728), .B1(new_n597), .B2(new_n588), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n601), .A2(new_n733), .B1(new_n590), .B2(new_n728), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n541), .A2(new_n726), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n597), .A2(new_n599), .A3(new_n588), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n563), .B1(new_n566), .B2(G169), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n738), .B1(new_n597), .B2(new_n588), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n736), .A2(new_n740), .B1(new_n739), .B2(new_n728), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n735), .A2(new_n741), .ZN(G399));
  INV_X1    g0542(.A(new_n209), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G41), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n655), .A2(G116), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n745), .A2(G1), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n212), .B2(new_n745), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT28), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n726), .B1(new_n711), .B2(new_n715), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT29), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n705), .A2(new_n706), .A3(new_n692), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT26), .ZN(new_n754));
  INV_X1    g0554(.A(new_n673), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n663), .A2(new_n670), .A3(new_n671), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n756), .A3(new_n707), .A4(new_n706), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n754), .A2(new_n757), .A3(new_n699), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n715), .B2(KEYINPUT96), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT96), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n712), .A2(new_n714), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n726), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n752), .B1(new_n762), .B2(new_n751), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n740), .A2(new_n674), .A3(new_n636), .A4(new_n728), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(new_n549), .B2(new_n554), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n627), .A2(new_n562), .A3(new_n560), .A4(new_n685), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n767), .B1(new_n768), .B2(new_n524), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n627), .A2(new_n685), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n523), .A2(G179), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n770), .A2(new_n567), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NOR3_X1   g0573(.A1(new_n768), .A2(new_n767), .A3(new_n524), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n726), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT31), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n766), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n763), .B1(G330), .B2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n749), .B1(new_n778), .B2(G1), .ZN(G364));
  INV_X1    g0579(.A(G13), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n205), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n744), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n732), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n730), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(G330), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n214), .B1(G20), .B2(new_n434), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n206), .A2(new_n304), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n384), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n206), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(new_n384), .A3(G200), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(G50), .B1(new_n794), .B2(G107), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n384), .A2(G179), .A3(G200), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n206), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G97), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n790), .A2(G190), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n795), .B(new_n799), .C1(new_n218), .C2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(G190), .A2(G200), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n792), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G159), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n804), .A2(KEYINPUT32), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G87), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT32), .B1(new_n804), .B2(new_n805), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n789), .A2(new_n803), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n789), .A2(G190), .A3(new_n349), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n248), .B1(new_n812), .B2(new_n251), .C1(new_n411), .C2(new_n813), .ZN(new_n814));
  NOR4_X1   g0614(.A1(new_n802), .A2(new_n806), .A3(new_n811), .A4(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n813), .ZN(new_n816));
  INV_X1    g0616(.A(new_n804), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n816), .A2(G322), .B1(new_n817), .B2(G329), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n505), .C1(new_n819), .C2(new_n812), .ZN(new_n820));
  INV_X1    g0620(.A(G317), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(KEYINPUT33), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(KEYINPUT33), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n800), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n791), .A2(G326), .ZN(new_n825));
  INV_X1    g0625(.A(G303), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n807), .ZN(new_n827));
  INV_X1    g0627(.A(G294), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n797), .A2(new_n828), .B1(new_n793), .B2(new_n829), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n820), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n788), .B1(new_n815), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n209), .A2(new_n248), .ZN(new_n833));
  INV_X1    g0633(.A(G355), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n833), .A2(new_n834), .B1(G116), .B2(new_n209), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n743), .A2(new_n406), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n513), .B2(new_n213), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n238), .A2(new_n513), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n835), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(G13), .A2(G33), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(G20), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n844), .A2(new_n788), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT97), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n784), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n844), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n832), .B(new_n849), .C1(new_n786), .C2(new_n850), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n787), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(G396));
  NAND2_X1  g0653(.A1(new_n777), .A2(G330), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n470), .A2(new_n726), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n473), .A2(new_n476), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT99), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n473), .A2(new_n476), .A3(new_n858), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n712), .A2(new_n714), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n728), .B(new_n860), .C1(new_n861), .C2(new_n710), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n857), .B(new_n859), .C1(new_n473), .C2(new_n728), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n862), .B1(new_n750), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n784), .B1(new_n854), .B2(new_n864), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n788), .A2(new_n842), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n784), .B1(G77), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n791), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n829), .A2(new_n801), .B1(new_n871), .B2(new_n826), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G107), .B2(new_n808), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n813), .A2(new_n828), .B1(new_n804), .B2(new_n819), .ZN(new_n874));
  INV_X1    g0674(.A(new_n812), .ZN(new_n875));
  AOI211_X1 g0675(.A(new_n248), .B(new_n874), .C1(G116), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n794), .A2(G87), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n873), .A2(new_n799), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n816), .A2(G143), .B1(new_n875), .B2(G159), .ZN(new_n879));
  INV_X1    g0679(.A(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n879), .B1(new_n871), .B2(new_n880), .C1(new_n881), .C2(new_n801), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT34), .Z(new_n883));
  NAND2_X1  g0683(.A1(new_n794), .A2(G68), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n276), .B2(new_n807), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n885), .A2(KEYINPUT98), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(KEYINPUT98), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n798), .A2(G58), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n401), .B1(G132), .B2(new_n817), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n886), .A2(new_n887), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n878), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n870), .B1(new_n891), .B2(new_n788), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n863), .B2(new_n843), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT100), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n867), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(G384));
  NOR2_X1   g0696(.A1(new_n781), .A2(new_n205), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n429), .A2(new_n430), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT16), .B1(new_n410), .B2(new_n419), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n899), .A2(new_n274), .A3(new_n438), .ZN(new_n900));
  INV_X1    g0700(.A(new_n724), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n900), .A2(new_n398), .B1(new_n435), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n898), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n435), .A2(new_n444), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n444), .A2(new_n901), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n904), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n903), .A2(KEYINPUT37), .B1(new_n898), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n900), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n724), .B1(new_n910), .B2(new_n436), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n453), .A2(KEYINPUT103), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT103), .B1(new_n453), .B2(new_n911), .ZN(new_n913));
  OAI211_X1 g0713(.A(KEYINPUT38), .B(new_n909), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n453), .A2(new_n911), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n453), .A2(KEYINPUT103), .A3(new_n911), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT104), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n920), .A2(new_n921), .A3(KEYINPUT38), .A4(new_n909), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n453), .A2(new_n444), .A3(new_n901), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n394), .A2(new_n428), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n904), .A2(new_n924), .A3(new_n906), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n923), .A2(KEYINPUT37), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT38), .B1(new_n898), .B2(new_n907), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n915), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n347), .A2(new_n728), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n364), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n355), .B(new_n363), .C1(new_n347), .C2(new_n728), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n764), .B1(new_n719), .B2(new_n720), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT31), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n775), .B(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n933), .B(new_n863), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n929), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n937), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n920), .B2(new_n909), .ZN(new_n942));
  INV_X1    g0742(.A(new_n914), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n940), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n777), .A2(new_n478), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT105), .Z(new_n947));
  AOI21_X1  g0747(.A(new_n731), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n931), .A2(new_n932), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n473), .A2(new_n726), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n862), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n942), .B2(new_n943), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n677), .A2(new_n724), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n363), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n728), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT39), .B1(new_n942), .B2(new_n943), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT39), .B1(new_n926), .B2(new_n927), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n915), .A2(new_n922), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n956), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n683), .B1(new_n763), .B2(new_n478), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n897), .B1(new_n949), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n949), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n276), .A2(G68), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT102), .Z(new_n970));
  NOR3_X1   g0770(.A1(new_n412), .A2(new_n212), .A3(new_n251), .ZN(new_n971));
  OAI211_X1 g0771(.A(G1), .B(new_n780), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n606), .A2(KEYINPUT35), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n973), .A2(G116), .A3(new_n215), .A4(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(KEYINPUT101), .B(KEYINPUT36), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n975), .B(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n968), .A2(new_n972), .A3(new_n977), .ZN(G367));
  AOI21_X1  g0778(.A(new_n632), .B1(new_n615), .B2(new_n726), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT107), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n628), .B2(new_n728), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n741), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT45), .Z(new_n983));
  NOR2_X1   g0783(.A1(new_n981), .A2(new_n741), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT44), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(new_n735), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n736), .A2(new_n740), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n734), .B2(new_n736), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n732), .B(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n778), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n991), .A2(new_n778), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n744), .B(KEYINPUT41), .Z(new_n993));
  OAI21_X1  g0793(.A(new_n782), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n705), .A2(new_n692), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n659), .A2(new_n728), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT106), .ZN(new_n997));
  MUX2_X1   g0797(.A(new_n995), .B(new_n699), .S(new_n997), .Z(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n980), .A2(new_n590), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n726), .B1(new_n1001), .B2(new_n628), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n981), .A2(new_n740), .A3(new_n736), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1002), .B1(new_n1003), .B2(KEYINPUT42), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n998), .A2(new_n999), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n732), .A2(new_n734), .A3(new_n981), .ZN(new_n1009));
  OR3_X1    g0809(.A1(new_n1008), .A2(KEYINPUT108), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(KEYINPUT108), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n994), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n466), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n845), .B1(new_n209), .B2(new_n1015), .C1(new_n837), .C2(new_n234), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT109), .Z(new_n1017));
  OAI22_X1  g0817(.A1(new_n828), .A2(new_n801), .B1(new_n871), .B2(new_n819), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G97), .B2(new_n794), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n808), .A2(G116), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT46), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n813), .A2(new_n826), .B1(new_n812), .B2(new_n829), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G317), .B2(new_n817), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n406), .B1(new_n798), .B2(G107), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n797), .A2(new_n218), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n505), .B(new_n1026), .C1(G150), .C2(new_n816), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n808), .A2(G58), .B1(new_n817), .B2(G137), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT111), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(KEYINPUT111), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n791), .A2(G143), .B1(new_n794), .B2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n800), .A2(G159), .B1(new_n875), .B2(G50), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT110), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1025), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT47), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n848), .B(new_n1017), .C1(new_n1036), .C2(new_n788), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT112), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n998), .A2(new_n844), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT113), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1014), .A2(new_n1042), .ZN(G387));
  AOI21_X1  g0843(.A(new_n745), .B1(new_n990), .B2(new_n778), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n778), .B2(new_n990), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n734), .A2(new_n850), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n833), .A2(new_n746), .B1(G107), .B2(new_n209), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n231), .A2(new_n513), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n746), .ZN(new_n1049));
  AOI211_X1 g0849(.A(G45), .B(new_n1049), .C1(G68), .C2(G77), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n279), .A2(G50), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT50), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n837), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1047), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n784), .B1(new_n1054), .B2(new_n846), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n798), .A2(new_n466), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n276), .B2(new_n813), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT114), .Z(new_n1058));
  OAI221_X1 g0858(.A(new_n406), .B1(new_n218), .B2(new_n812), .C1(new_n881), .C2(new_n804), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n791), .A2(G159), .B1(new_n808), .B2(G77), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n489), .B2(new_n793), .C1(new_n279), .C2(new_n801), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n406), .B1(G326), .B2(new_n817), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n797), .A2(new_n829), .B1(new_n807), .B2(new_n828), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n816), .A2(G317), .B1(new_n875), .B2(G303), .ZN(new_n1065));
  INV_X1    g0865(.A(G322), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1065), .B1(new_n871), .B2(new_n1066), .C1(new_n819), .C2(new_n801), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1063), .B1(new_n484), .B2(new_n793), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1062), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1055), .B1(new_n1074), .B2(new_n788), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n990), .A2(new_n783), .B1(new_n1046), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1045), .A2(new_n1076), .ZN(G393));
  OR2_X1    g0877(.A1(new_n981), .A2(new_n850), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n845), .B1(new_n489), .B2(new_n209), .C1(new_n837), .C2(new_n241), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n784), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n797), .A2(new_n251), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n877), .B1(new_n218), .B2(new_n807), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G50), .C2(new_n800), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n280), .A2(new_n875), .B1(new_n817), .B2(G143), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G150), .A2(new_n791), .B1(new_n816), .B2(G159), .ZN(new_n1085));
  XOR2_X1   g0885(.A(KEYINPUT115), .B(KEYINPUT51), .Z(new_n1086));
  XNOR2_X1  g0886(.A(new_n1085), .B(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n406), .A3(new_n1084), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G317), .A2(new_n791), .B1(new_n816), .B2(G311), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n801), .A2(new_n826), .B1(new_n484), .B2(new_n797), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n505), .B1(new_n804), .B2(new_n1066), .C1(new_n828), .C2(new_n812), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n456), .A2(new_n793), .B1(new_n807), .B2(new_n829), .ZN(new_n1093));
  OR3_X1    g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1088), .B1(new_n1090), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1080), .B1(new_n1095), .B2(new_n788), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n987), .A2(new_n783), .B1(new_n1078), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n991), .A2(new_n744), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n987), .B1(new_n778), .B2(new_n990), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G390));
  INV_X1    g0900(.A(new_n860), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n726), .B(new_n1101), .C1(new_n759), .C2(new_n761), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n933), .B1(new_n1102), .B2(new_n951), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n958), .A3(new_n929), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n951), .B1(new_n750), .B2(new_n860), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n958), .B1(new_n1105), .B2(new_n950), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n960), .A2(new_n1106), .A3(new_n962), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n863), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n766), .B2(new_n776), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(KEYINPUT116), .A3(G330), .A4(new_n933), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT116), .ZN(new_n1111));
  OAI211_X1 g0911(.A(G330), .B(new_n863), .C1(new_n934), .C2(new_n936), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1112), .B2(new_n950), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1104), .A2(new_n1107), .A3(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n777), .A2(G330), .A3(new_n863), .A4(new_n933), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1104), .B2(new_n1107), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n960), .A2(new_n962), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n842), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n784), .B1(new_n280), .B2(new_n869), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1122), .A2(new_n871), .B1(new_n801), .B2(new_n880), .ZN(new_n1123));
  INV_X1    g0923(.A(G132), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n797), .A2(new_n805), .B1(new_n813), .B2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT121), .B(KEYINPUT53), .Z(new_n1127));
  NAND3_X1  g0927(.A1(new_n808), .A2(G150), .A3(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT119), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n875), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1127), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n881), .B2(new_n807), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G125), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n248), .B1(new_n804), .B2(new_n1135), .C1(new_n276), .C2(new_n793), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT120), .Z(new_n1137));
  OAI22_X1  g0937(.A1(new_n813), .A2(new_n484), .B1(new_n804), .B2(new_n828), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n248), .B(new_n1138), .C1(G97), .C2(new_n875), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(new_n809), .A3(new_n884), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1081), .B1(G283), .B2(new_n791), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n456), .B2(new_n801), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1134), .A2(new_n1137), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1121), .B1(new_n1143), .B2(new_n788), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1118), .A2(new_n783), .B1(new_n1120), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT118), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1116), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1104), .A2(new_n1107), .A3(new_n1114), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n951), .B1(new_n762), .B2(new_n860), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1112), .A2(new_n950), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1110), .A2(new_n1113), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1116), .A2(new_n1153), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1105), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT117), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT117), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1158), .B(new_n1105), .C1(new_n1116), .C2(new_n1153), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1154), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n777), .A2(new_n478), .A3(G330), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n965), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n745), .B1(new_n1151), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1149), .A2(new_n1160), .A3(new_n1150), .A4(new_n1163), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1146), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND4_X1   g0967(.A1(new_n1152), .A2(new_n1110), .A3(new_n1113), .A4(new_n1153), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1158), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1155), .A2(KEYINPUT117), .A3(new_n1156), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1172), .A2(new_n1162), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1173));
  AND4_X1   g0973(.A1(new_n1146), .A2(new_n1173), .A3(new_n744), .A4(new_n1166), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1145), .B1(new_n1167), .B2(new_n1174), .ZN(G378));
  OAI211_X1 g0975(.A(new_n954), .B(new_n955), .C1(new_n1119), .C2(new_n958), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT38), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n937), .B1(new_n1179), .B2(new_n914), .ZN(new_n1180));
  OAI21_X1  g0980(.A(G330), .B1(new_n1180), .B2(KEYINPUT40), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n294), .A2(new_n724), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT125), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n312), .B(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(new_n940), .A2(new_n1181), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n731), .B1(new_n944), .B2(new_n938), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n929), .A2(new_n939), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1176), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1186), .B1(new_n940), .B2(new_n1181), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1189), .A2(new_n1190), .A3(new_n1188), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n964), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1186), .A2(new_n842), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n869), .A2(G50), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n406), .A2(G41), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G50), .B(new_n1199), .C1(new_n245), .C2(new_n255), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n816), .A2(G107), .B1(new_n817), .B2(G283), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n1015), .B2(new_n812), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1026), .B(new_n1202), .C1(G77), .C2(new_n808), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n871), .A2(new_n484), .B1(new_n793), .B2(new_n411), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(G97), .B2(new_n800), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1205), .A3(new_n1199), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT122), .Z(new_n1207));
  XNOR2_X1  g1007(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1200), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n791), .A2(G125), .B1(new_n875), .B2(G137), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(G150), .A2(new_n798), .B1(new_n800), .B2(G132), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1130), .A2(new_n808), .B1(G128), .B2(new_n816), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1212), .A2(KEYINPUT124), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(KEYINPUT124), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1210), .B(new_n1211), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n794), .A2(G159), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n817), .C2(G124), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1209), .B1(new_n1216), .B2(new_n1220), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n848), .B(new_n1198), .C1(new_n1221), .C2(new_n788), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1196), .A2(new_n783), .B1(new_n1197), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1193), .A2(new_n964), .A3(new_n1194), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n964), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1162), .B1(new_n1118), .B2(new_n1160), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n744), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1166), .A2(new_n1163), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1229), .B2(new_n1196), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1223), .B1(new_n1228), .B2(new_n1230), .ZN(G375));
  OAI211_X1 g1031(.A(new_n1162), .B(new_n1154), .C1(new_n1157), .C2(new_n1159), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT126), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n993), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1164), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT127), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n484), .A2(new_n801), .B1(new_n871), .B2(new_n828), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(G97), .B2(new_n808), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n794), .A2(G77), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n813), .A2(new_n829), .B1(new_n812), .B2(new_n456), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n248), .B(new_n1240), .C1(G303), .C2(new_n817), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1239), .A3(new_n1056), .A4(new_n1241), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n871), .A2(new_n1124), .B1(new_n807), .B2(new_n805), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G50), .B2(new_n798), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n812), .A2(new_n881), .B1(new_n804), .B2(new_n1122), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G137), .B2(new_n816), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1130), .A2(new_n800), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n401), .B1(G58), .B2(new_n794), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1244), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n788), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n848), .B1(new_n218), .B2(new_n868), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n933), .C2(new_n843), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n1172), .B2(new_n782), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1236), .A2(new_n1255), .ZN(G381));
  NAND2_X1  g1056(.A1(new_n1197), .A2(new_n1222), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n782), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT57), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1260), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n745), .B1(new_n1261), .B2(new_n1229), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1260), .B1(new_n1258), .B2(new_n1227), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1259), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1173), .A2(new_n744), .A3(new_n1166), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(new_n1145), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1264), .A2(new_n1267), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1045), .A2(new_n852), .A3(new_n1076), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1269), .A2(new_n895), .A3(new_n1097), .A4(new_n1271), .ZN(new_n1272));
  OR4_X1    g1072(.A1(G387), .A2(G381), .A3(new_n1268), .A4(new_n1272), .ZN(G407));
  OAI211_X1 g1073(.A(G407), .B(G213), .C1(G343), .C2(new_n1268), .ZN(G409));
  NAND3_X1  g1074(.A1(new_n1229), .A2(new_n1196), .A3(new_n1234), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1223), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1267), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1120), .A2(new_n1144), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1151), .B2(new_n782), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1265), .A2(KEYINPUT118), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1165), .A2(new_n1146), .A3(new_n1166), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1277), .B1(G375), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(G213), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1284), .A2(G343), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1232), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1164), .A2(KEYINPUT60), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT126), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1232), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT60), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n744), .B1(new_n1232), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1292), .A2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(G384), .B1(new_n1296), .B2(new_n1255), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n895), .B(new_n1254), .C1(new_n1292), .C2(new_n1295), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1283), .A2(new_n1286), .A3(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(KEYINPUT62), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT61), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1283), .A2(new_n1303), .A3(new_n1299), .A4(new_n1286), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1294), .B1(new_n1233), .B2(new_n1289), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n895), .B1(new_n1305), .B2(new_n1254), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1296), .A2(G384), .A3(new_n1255), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1285), .A2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1308), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1266), .B1(new_n1223), .B2(new_n1275), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1264), .B2(G378), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1309), .B(new_n1311), .C1(new_n1313), .C2(new_n1285), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1301), .A2(new_n1302), .A3(new_n1304), .A4(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n852), .B1(new_n1045), .B2(new_n1076), .ZN(new_n1316));
  OAI211_X1 g1116(.A(new_n1269), .B(new_n1097), .C1(new_n1271), .C2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1316), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(G390), .A2(new_n1270), .A3(new_n1318), .ZN(new_n1319));
  AND4_X1   g1119(.A1(new_n1042), .A2(new_n1317), .A3(new_n1014), .A4(new_n1319), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1317), .A2(new_n1319), .B1(new_n1014), .B2(new_n1042), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1315), .A2(new_n1323), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1311), .A2(new_n1309), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1300), .A2(new_n1328), .ZN(new_n1329));
  NAND4_X1  g1129(.A1(new_n1283), .A2(KEYINPUT63), .A3(new_n1299), .A4(new_n1286), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1327), .A2(new_n1322), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1324), .A2(new_n1331), .ZN(G405));
  NAND2_X1  g1132(.A1(new_n1264), .A2(G378), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(G375), .A2(new_n1267), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1299), .ZN(new_n1336));
  OAI211_X1 g1136(.A(new_n1333), .B(new_n1334), .C1(new_n1297), .C2(new_n1298), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1337), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1323), .B(new_n1338), .ZN(G402));
endmodule


