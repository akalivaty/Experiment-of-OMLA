//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202));
  XNOR2_X1  g001(.A(G141gat), .B(G148gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  AOI21_X1  g003(.A(new_n203), .B1(KEYINPUT2), .B2(new_n204), .ZN(new_n205));
  OR2_X1    g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n204), .B(new_n206), .C1(new_n203), .C2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n205), .A2(new_n208), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT73), .ZN(new_n212));
  INV_X1    g011(.A(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G127gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT67), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT68), .B(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(new_n213), .ZN(new_n217));
  XNOR2_X1  g016(.A(G113gat), .B(G120gat), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n215), .A2(new_n217), .B1(KEYINPUT1), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT1), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n220), .B1(new_n213), .B2(G127gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT69), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n221), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G113gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n224), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n214), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n219), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n212), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G225gat), .A2(G233gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n228), .B1(KEYINPUT3), .B2(new_n211), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n211), .A2(new_n227), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n229), .B(new_n230), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n230), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n209), .A2(new_n210), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(new_n228), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n239), .B2(new_n235), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT74), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT74), .B(new_n237), .C1(new_n239), .C2(new_n235), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n244), .A3(KEYINPUT5), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n235), .A2(KEYINPUT4), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n237), .A2(KEYINPUT5), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT73), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n211), .B(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n249), .A2(new_n227), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n246), .B(new_n247), .C1(new_n250), .C2(new_n234), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT0), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G57gat), .ZN(new_n255));
  INV_X1    g054(.A(G85gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n202), .B1(new_n260), .B2(KEYINPUT6), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT6), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n245), .A2(new_n257), .A3(new_n251), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n262), .B2(new_n259), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n261), .B1(new_n265), .B2(new_n202), .ZN(new_n266));
  INV_X1    g065(.A(G169gat), .ZN(new_n267));
  INV_X1    g066(.A(G176gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(G169gat), .A2(G176gat), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n269), .B1(KEYINPUT23), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  OR2_X1    g072(.A1(new_n270), .A2(KEYINPUT23), .ZN(new_n274));
  NAND2_X1  g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n275), .B(KEYINPUT24), .Z(new_n276));
  NOR2_X1   g075(.A1(G183gat), .A2(G190gat), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n274), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(new_n277), .B(KEYINPUT64), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n271), .B(new_n274), .C1(new_n276), .C2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  INV_X1    g084(.A(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n287), .B(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT26), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n291), .B(new_n292), .C1(new_n267), .C2(new_n268), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n289), .A2(new_n275), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n284), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n289), .A2(new_n300), .A3(new_n275), .A4(new_n293), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n284), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n298), .B1(new_n303), .B2(new_n297), .ZN(new_n304));
  XNOR2_X1  g103(.A(G197gat), .B(G204gat), .ZN(new_n305));
  INV_X1    g104(.A(G211gat), .ZN(new_n306));
  INV_X1    g105(.A(G218gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(KEYINPUT22), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G211gat), .B(G218gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n299), .A2(new_n301), .B1(new_n283), .B2(new_n279), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n297), .B1(new_n313), .B2(KEYINPUT29), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n295), .A2(G226gat), .A3(G233gat), .ZN(new_n317));
  OAI211_X1 g116(.A(KEYINPUT70), .B(new_n297), .C1(new_n313), .C2(KEYINPUT29), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n311), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n312), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G8gat), .B(G36gat), .ZN(new_n322));
  INV_X1    g121(.A(G64gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(G92gat), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n321), .A2(KEYINPUT71), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT71), .B1(new_n321), .B2(new_n325), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT37), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n319), .B2(new_n320), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n304), .A2(new_n311), .ZN(new_n331));
  AND3_X1   g130(.A1(new_n330), .A2(KEYINPUT78), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT78), .B1(new_n330), .B2(new_n331), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n325), .B1(new_n321), .B2(new_n329), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT38), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n321), .A2(new_n329), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n337), .A2(KEYINPUT38), .A3(new_n335), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n266), .B(new_n328), .C1(new_n336), .C2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n311), .B1(new_n340), .B2(KEYINPUT29), .ZN(new_n341));
  NAND2_X1  g140(.A1(G228gat), .A2(G233gat), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT3), .B1(new_n320), .B2(new_n296), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n341), .B(new_n342), .C1(new_n212), .C2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n320), .B1(new_n233), .B2(new_n296), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n343), .A2(new_n238), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n344), .B1(new_n347), .B2(new_n342), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n348), .A2(G22gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(G22gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(KEYINPUT75), .A3(new_n350), .ZN(new_n354));
  XNOR2_X1  g153(.A(G78gat), .B(G106gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT31), .B(G50gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n351), .A2(new_n352), .A3(new_n357), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n246), .B1(new_n250), .B2(new_n234), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n237), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(KEYINPUT39), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n365), .A2(new_n258), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n239), .A2(new_n235), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n364), .B(KEYINPUT39), .C1(new_n237), .C2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT40), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n259), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g170(.A(KEYINPUT77), .B(KEYINPUT40), .C1(new_n366), .C2(new_n368), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT30), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n326), .B2(new_n327), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n321), .A2(KEYINPUT30), .A3(new_n325), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n321), .A2(new_n325), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n366), .A2(KEYINPUT40), .A3(new_n368), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n339), .A2(new_n362), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n303), .A2(new_n228), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n313), .A2(new_n227), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n385), .B1(G227gat), .B2(G233gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(G227gat), .A3(G233gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT34), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n387), .A2(KEYINPUT32), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n387), .B2(KEYINPUT32), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(KEYINPUT32), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT34), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(KEYINPUT32), .A3(new_n388), .ZN(new_n394));
  INV_X1    g193(.A(new_n386), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n399), .B(G71gat), .ZN(new_n400));
  INV_X1    g199(.A(G99gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n391), .A2(new_n396), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n404), .B1(new_n391), .B2(new_n396), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT36), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT36), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n405), .B2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n361), .B(KEYINPUT76), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n265), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n381), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n406), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n391), .A2(new_n396), .A3(new_n404), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n362), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT35), .B1(new_n414), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n266), .A2(new_n378), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT35), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n407), .A4(new_n362), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G1gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT16), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n427), .B(KEYINPUT85), .ZN(new_n428));
  XOR2_X1   g227(.A(G15gat), .B(G22gat), .Z(new_n429));
  OR2_X1    g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(G8gat), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n426), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n433), .B(KEYINPUT87), .Z(new_n434));
  NAND3_X1  g233(.A1(new_n430), .A2(KEYINPUT86), .A3(new_n432), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(G8gat), .C1(KEYINPUT86), .C2(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(G43gat), .B(G50gat), .Z(new_n439));
  INV_X1    g238(.A(KEYINPUT15), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n441), .B1(G29gat), .B2(G36gat), .ZN(new_n442));
  OR3_X1    g241(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n439), .A2(new_n440), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n444), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n443), .B2(KEYINPUT83), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(KEYINPUT83), .B2(new_n443), .ZN(new_n450));
  NAND2_X1  g249(.A1(G29gat), .A2(G36gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT84), .ZN(new_n453));
  AND3_X1   g252(.A1(new_n452), .A2(new_n453), .A3(new_n441), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n452), .B2(new_n441), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n447), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n438), .B(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(G229gat), .A2(G233gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT13), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT17), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n456), .A2(new_n461), .ZN(new_n462));
  OAI211_X1 g261(.A(KEYINPUT17), .B(new_n447), .C1(new_n454), .C2(new_n455), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n438), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n437), .A2(new_n456), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n458), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT18), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n467), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n460), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(KEYINPUT81), .ZN(new_n472));
  XNOR2_X1  g271(.A(G113gat), .B(G141gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(G169gat), .B(G197gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n474), .B(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n460), .A2(new_n468), .A3(new_n478), .A4(new_n469), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n425), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT7), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT7), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n488), .A2(KEYINPUT95), .A3(G85gat), .A4(G92gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491));
  INV_X1    g290(.A(G92gat), .ZN(new_n492));
  AOI22_X1  g291(.A1(KEYINPUT8), .A2(new_n491), .B1(new_n256), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G99gat), .B(G106gat), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n490), .A2(new_n495), .A3(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n462), .A2(new_n499), .A3(new_n463), .ZN(new_n500));
  INV_X1    g299(.A(new_n499), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n456), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(KEYINPUT93), .Z(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT41), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G190gat), .B(G218gat), .Z(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT97), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n505), .A2(KEYINPUT41), .ZN(new_n513));
  XNOR2_X1  g312(.A(G134gat), .B(G162gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n507), .A2(KEYINPUT97), .A3(new_n509), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n500), .A2(new_n508), .A3(new_n502), .A4(new_n506), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n512), .A2(new_n515), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n517), .A2(KEYINPUT96), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(KEYINPUT96), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n512), .A2(new_n520), .A3(new_n516), .A4(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n515), .B(KEYINPUT94), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT98), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n526), .A3(new_n523), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n519), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G231gat), .ZN(new_n529));
  INV_X1    g328(.A(G233gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(KEYINPUT89), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(G71gat), .A3(G78gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n323), .A2(G57gat), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G64gat), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT90), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT90), .B1(new_n538), .B2(new_n540), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(KEYINPUT89), .A2(KEYINPUT9), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n537), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n533), .A2(KEYINPUT9), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n546), .A2(new_n532), .B1(new_n538), .B2(new_n540), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n434), .A2(new_n549), .A3(new_n436), .ZN(new_n550));
  OR2_X1    g349(.A1(new_n550), .A2(KEYINPUT92), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(KEYINPUT92), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n531), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n531), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n554), .B(new_n555), .C1(KEYINPUT21), .C2(new_n548), .ZN(new_n556));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT91), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT19), .ZN(new_n559));
  XNOR2_X1  g358(.A(G127gat), .B(G155gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT20), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n563));
  INV_X1    g362(.A(new_n555), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n553), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n556), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n562), .B1(new_n556), .B2(new_n565), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n528), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n499), .B1(new_n545), .B2(new_n547), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n538), .A2(new_n540), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT90), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n544), .A3(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n537), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n547), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n498), .A4(new_n497), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n571), .A2(new_n572), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT99), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n548), .A2(KEYINPUT10), .A3(new_n501), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n571), .A2(new_n581), .A3(new_n585), .A4(new_n572), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G230gat), .A2(G233gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n571), .A2(new_n581), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G120gat), .B(G148gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT100), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G176gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G204gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n591), .B(new_n595), .Z(new_n596));
  NAND3_X1  g395(.A1(new_n425), .A2(KEYINPUT88), .A3(new_n482), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n485), .A2(new_n570), .A3(new_n596), .A4(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(KEYINPUT101), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT88), .B1(new_n425), .B2(new_n482), .ZN(new_n600));
  INV_X1    g399(.A(new_n482), .ZN(new_n601));
  AOI211_X1 g400(.A(new_n484), .B(new_n601), .C1(new_n416), .C2(new_n424), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n603), .A2(new_n604), .A3(new_n570), .A4(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n265), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g408(.A1(new_n606), .A2(new_n378), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G8gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT16), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n431), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n431), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n606), .A2(new_n378), .A3(new_n613), .A4(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT42), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT103), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI211_X1 g417(.A(new_n413), .B(new_n614), .C1(new_n599), .C2(new_n605), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT103), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT42), .A4(new_n613), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n617), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n623), .A2(KEYINPUT102), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(KEYINPUT102), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n611), .B(new_n622), .C1(new_n624), .C2(new_n625), .ZN(G1325gat));
  AOI21_X1  g425(.A(G15gat), .B1(new_n606), .B2(new_n407), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n411), .B1(new_n599), .B2(new_n605), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(G15gat), .B2(new_n628), .ZN(G1326gat));
  NAND2_X1  g428(.A1(new_n606), .A2(new_n412), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT43), .B(G22gat), .Z(new_n631));
  OR2_X1    g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n635), .A3(new_n633), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(G1327gat));
  NOR3_X1   g438(.A1(new_n600), .A2(new_n602), .A3(new_n528), .ZN(new_n640));
  INV_X1    g439(.A(new_n596), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n568), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n643), .A2(G29gat), .A3(new_n265), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT106), .B(KEYINPUT45), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n528), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n425), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g447(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(KEYINPUT44), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n482), .B(new_n642), .C1(new_n649), .C2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G29gat), .B1(new_n651), .B2(new_n265), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n646), .A2(new_n652), .ZN(G1328gat));
  NOR3_X1   g452(.A1(new_n643), .A2(G36gat), .A3(new_n413), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT46), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n656), .A2(KEYINPUT107), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(KEYINPUT107), .ZN(new_n659));
  OAI21_X1  g458(.A(G36gat), .B1(new_n651), .B2(new_n413), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n657), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(G1329gat));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662));
  OAI21_X1  g461(.A(G43gat), .B1(new_n651), .B2(new_n411), .ZN(new_n663));
  INV_X1    g462(.A(G43gat), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n640), .A2(new_n664), .A3(new_n407), .A4(new_n642), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n663), .A2(new_n662), .A3(new_n665), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n667), .A2(KEYINPUT47), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT47), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(G1330gat));
  INV_X1    g470(.A(new_n412), .ZN(new_n672));
  OR3_X1    g471(.A1(new_n643), .A2(G50gat), .A3(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(G50gat), .B1(new_n651), .B2(new_n362), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(KEYINPUT48), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G50gat), .B1(new_n651), .B2(new_n672), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n675), .B1(new_n677), .B2(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g477(.A1(new_n570), .A2(new_n425), .A3(new_n641), .A4(new_n601), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n607), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(G57gat), .ZN(G1332gat));
  INV_X1    g480(.A(KEYINPUT49), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n679), .B(new_n378), .C1(new_n682), .C2(new_n323), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n323), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1333gat));
  AOI21_X1  g484(.A(G71gat), .B1(new_n679), .B2(new_n407), .ZN(new_n686));
  INV_X1    g485(.A(new_n411), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(G71gat), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(new_n679), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g489(.A1(new_n679), .A2(new_n412), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G78gat), .ZN(G1335gat));
  INV_X1    g491(.A(new_n568), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n601), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT109), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n425), .A2(new_n647), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT51), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(KEYINPUT110), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n698), .A2(KEYINPUT110), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n699), .A2(new_n700), .A3(new_n596), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n256), .A3(new_n607), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n641), .B(new_n695), .C1(new_n649), .C2(new_n650), .ZN(new_n703));
  OAI21_X1  g502(.A(G85gat), .B1(new_n703), .B2(new_n265), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1336gat));
  OAI21_X1  g504(.A(G92gat), .B1(new_n703), .B2(new_n413), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n378), .A2(new_n492), .A3(new_n641), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n706), .B1(new_n697), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT52), .ZN(G1337gat));
  NAND3_X1  g508(.A1(new_n701), .A2(new_n401), .A3(new_n407), .ZN(new_n710));
  OAI21_X1  g509(.A(G99gat), .B1(new_n703), .B2(new_n411), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1338gat));
  NOR3_X1   g511(.A1(new_n362), .A2(G106gat), .A3(new_n596), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT112), .ZN(new_n715));
  OAI21_X1  g514(.A(G106gat), .B1(new_n703), .B2(new_n362), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT53), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n714), .A2(KEYINPUT112), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n703), .A2(new_n672), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n713), .B(KEYINPUT111), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n720), .A2(G106gat), .B1(new_n698), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n722), .B2(new_n717), .ZN(G1339gat));
  NAND4_X1  g522(.A1(new_n601), .A2(new_n528), .A3(new_n568), .A4(new_n596), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT113), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n587), .A2(new_n588), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT54), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n729), .A2(new_n595), .ZN(new_n730));
  INV_X1    g529(.A(new_n588), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n583), .A2(new_n731), .A3(new_n584), .A4(new_n586), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n728), .B1(new_n732), .B2(new_n733), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT115), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n583), .A2(new_n586), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n738), .A2(KEYINPUT114), .A3(new_n731), .A4(new_n584), .ZN(new_n739));
  AND4_X1   g538(.A1(KEYINPUT115), .A2(new_n739), .A3(new_n736), .A4(new_n589), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n730), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT55), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n591), .A2(new_n595), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g544(.A(KEYINPUT55), .B(new_n730), .C1(new_n737), .C2(new_n740), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n482), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n457), .A2(new_n459), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n476), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n481), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n641), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n647), .B1(new_n749), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n748), .A2(new_n753), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(new_n528), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n693), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n726), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n759), .A2(new_n407), .A3(new_n672), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n378), .A2(new_n265), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G113gat), .B1(new_n762), .B2(new_n601), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n759), .A2(new_n761), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n419), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n482), .A2(new_n224), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT116), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n763), .B1(new_n766), .B2(new_n768), .ZN(G1340gat));
  OAI21_X1  g568(.A(G120gat), .B1(new_n762), .B2(new_n596), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n764), .A2(new_n596), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n419), .A2(G120gat), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(G1341gat));
  INV_X1    g573(.A(new_n216), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n762), .A2(new_n775), .A3(new_n693), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n216), .B1(new_n765), .B2(new_n568), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(G1342gat));
  NAND3_X1  g577(.A1(new_n765), .A2(new_n213), .A3(new_n647), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT56), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(KEYINPUT117), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n779), .A2(KEYINPUT56), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(KEYINPUT117), .ZN(new_n783));
  OAI21_X1  g582(.A(G134gat), .B1(new_n762), .B2(new_n528), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(G1343gat));
  INV_X1    g584(.A(G141gat), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n362), .B1(new_n726), .B2(new_n758), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n787), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT118), .B1(new_n787), .B2(KEYINPUT57), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT57), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n747), .A2(KEYINPUT119), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n743), .A2(new_n793), .A3(new_n745), .A4(new_n746), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n482), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n647), .B1(new_n795), .B2(new_n754), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n693), .B1(new_n796), .B2(new_n757), .ZN(new_n797));
  AOI211_X1 g596(.A(new_n791), .B(new_n672), .C1(new_n726), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n790), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n411), .A2(new_n761), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n786), .B1(new_n801), .B2(new_n482), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n764), .A2(new_n362), .A3(new_n687), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n803), .A2(new_n786), .A3(new_n482), .ZN(new_n804));
  OR3_X1    g603(.A1(new_n802), .A2(KEYINPUT58), .A3(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT58), .B1(new_n802), .B2(new_n804), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1344gat));
  INV_X1    g606(.A(G148gat), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n687), .A2(new_n362), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n771), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n754), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n528), .ZN(new_n813));
  INV_X1    g612(.A(new_n757), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(KEYINPUT120), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n796), .B2(new_n757), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n693), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n672), .B1(new_n818), .B2(new_n724), .ZN(new_n819));
  OAI21_X1  g618(.A(KEYINPUT121), .B1(new_n819), .B2(KEYINPUT57), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n787), .A2(KEYINPUT57), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822));
  INV_X1    g621(.A(new_n724), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n757), .B1(new_n812), .B2(new_n528), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n568), .B1(new_n824), .B2(KEYINPUT120), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(new_n817), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n822), .B(new_n791), .C1(new_n826), .C2(new_n672), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n820), .A2(new_n821), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n800), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n828), .A2(new_n641), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n811), .B1(new_n830), .B2(G148gat), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n641), .B(new_n829), .C1(new_n790), .C2(new_n798), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n832), .A2(new_n811), .A3(G148gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n810), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT122), .B(new_n810), .C1(new_n831), .C2(new_n833), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1345gat));
  AOI21_X1  g637(.A(G155gat), .B1(new_n803), .B2(new_n568), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n568), .A2(G155gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n801), .B2(new_n840), .ZN(G1346gat));
  AOI21_X1  g640(.A(G162gat), .B1(new_n803), .B2(new_n647), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n647), .A2(G162gat), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n801), .B2(new_n843), .ZN(G1347gat));
  NOR2_X1   g643(.A1(new_n413), .A2(new_n607), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n760), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT124), .ZN(new_n847));
  OAI21_X1  g646(.A(G169gat), .B1(new_n847), .B2(new_n601), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n759), .A2(new_n265), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT123), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(new_n378), .A3(new_n407), .A4(new_n362), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n482), .A2(new_n267), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(G1348gat));
  OAI21_X1  g652(.A(G176gat), .B1(new_n847), .B2(new_n596), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n641), .A2(new_n268), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n854), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n856), .B(new_n857), .ZN(G1349gat));
  INV_X1    g657(.A(new_n851), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n568), .A3(new_n285), .ZN(new_n860));
  OAI21_X1  g659(.A(G183gat), .B1(new_n847), .B2(new_n693), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g662(.A1(new_n859), .A2(new_n286), .A3(new_n647), .ZN(new_n864));
  OAI21_X1  g663(.A(G190gat), .B1(new_n847), .B2(new_n528), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n865), .A2(KEYINPUT61), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n865), .A2(KEYINPUT61), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(G1351gat));
  NAND2_X1  g667(.A1(new_n411), .A2(new_n845), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n828), .A2(new_n482), .A3(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT126), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(KEYINPUT126), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(G197gat), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n850), .A2(new_n378), .A3(new_n809), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n601), .A2(G197gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(G1352gat));
  NOR2_X1   g676(.A1(new_n875), .A2(G204gat), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT127), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n878), .A2(new_n641), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n828), .A2(new_n641), .A3(new_n870), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G204gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n881), .A2(new_n882), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n883), .A2(new_n885), .A3(new_n886), .ZN(G1353gat));
  INV_X1    g686(.A(new_n875), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n306), .A3(new_n568), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n828), .A2(new_n870), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n568), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n891), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT63), .B1(new_n891), .B2(G211gat), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n889), .B1(new_n892), .B2(new_n893), .ZN(G1354gat));
  AOI21_X1  g693(.A(G218gat), .B1(new_n888), .B2(new_n647), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n528), .A2(new_n307), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n890), .B2(new_n896), .ZN(G1355gat));
endmodule


