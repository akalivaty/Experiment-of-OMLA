//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(G227gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n209), .B(new_n210), .C1(new_n206), .C2(new_n207), .ZN(new_n211));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT27), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G183gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G190gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT28), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT65), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT28), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT27), .B1(new_n213), .B2(KEYINPUT67), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT67), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(new_n215), .A3(G183gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n224), .A2(new_n225), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n230));
  AND3_X1   g029(.A1(new_n219), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n219), .B2(new_n229), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n211), .B(new_n212), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(G183gat), .B1(new_n221), .B2(new_n223), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n234), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT23), .B1(new_n206), .B2(new_n207), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n208), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT25), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(G169gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n244), .B2(new_n207), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n239), .A2(KEYINPUT66), .A3(new_n241), .A4(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n238), .B1(new_n213), .B2(new_n220), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT64), .B(G176gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n241), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n242), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n241), .B(new_n245), .C1(new_n234), .C2(new_n238), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n246), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(KEYINPUT69), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G120gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n257), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G113gat), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(new_n265), .A3(new_n256), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n259), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G127gat), .ZN(new_n268));
  INV_X1    g067(.A(G127gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n259), .A2(new_n266), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(KEYINPUT70), .A3(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n259), .A2(new_n266), .A3(new_n269), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n259), .B2(new_n266), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n233), .A2(new_n255), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n233), .A2(new_n255), .B1(new_n275), .B2(new_n271), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n205), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT32), .ZN(new_n281));
  INV_X1    g080(.A(new_n205), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n233), .A2(new_n255), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n271), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n282), .B1(new_n285), .B2(new_n276), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT71), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G15gat), .B(G43gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(G71gat), .ZN(new_n290));
  INV_X1    g089(.A(G99gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT33), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n279), .A2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n281), .A2(new_n288), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(KEYINPUT33), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n279), .A2(KEYINPUT32), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n285), .A2(new_n282), .A3(new_n276), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n298), .B(KEYINPUT34), .Z(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n299), .B1(new_n295), .B2(new_n297), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n202), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n295), .A2(new_n297), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(KEYINPUT36), .A3(new_n300), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n303), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT3), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  INV_X1    g109(.A(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G155gat), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G162gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n312), .A2(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n317), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n323), .A2(new_n324), .A3(new_n316), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n321), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g126(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n310), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n310), .A2(KEYINPUT74), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT74), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(G141gat), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n311), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n309), .B(new_n319), .C1(new_n327), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT77), .ZN(new_n337));
  OR2_X1    g136(.A1(KEYINPUT76), .A2(G162gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n338), .A2(G155gat), .A3(new_n322), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n320), .B1(new_n339), .B2(KEYINPUT2), .ZN(new_n340));
  AND2_X1   g139(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT75), .A2(G148gat), .ZN(new_n342));
  OAI21_X1  g141(.A(G141gat), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT74), .B(G141gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(new_n311), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n318), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n309), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT29), .B1(new_n337), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G197gat), .B(G204gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351));
  INV_X1    g150(.A(G211gat), .ZN(new_n352));
  INV_X1    g151(.A(G218gat), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  XOR2_X1   g154(.A(G211gat), .B(G218gat), .Z(new_n356));
  OR2_X1    g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n356), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(KEYINPUT72), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT86), .B1(new_n349), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT29), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n345), .ZN(new_n363));
  AND4_X1   g162(.A1(new_n347), .A2(new_n363), .A3(new_n309), .A4(new_n319), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n347), .B1(new_n346), .B2(new_n309), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT72), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n359), .B(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n366), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n319), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n357), .A2(new_n358), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n372), .A2(KEYINPUT29), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n371), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n361), .A2(new_n370), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n309), .B1(new_n373), .B2(KEYINPUT85), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n359), .A2(KEYINPUT85), .A3(new_n362), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n371), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n376), .C1(new_n359), .C2(new_n349), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n378), .A2(new_n382), .A3(G22gat), .ZN(new_n383));
  AOI21_X1  g182(.A(G22gat), .B1(new_n378), .B2(new_n382), .ZN(new_n384));
  XOR2_X1   g183(.A(G78gat), .B(G106gat), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT84), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n386), .B(KEYINPUT31), .ZN(new_n387));
  INV_X1    g186(.A(G50gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  OAI22_X1  g188(.A1(new_n383), .A2(new_n384), .B1(KEYINPUT87), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n378), .A2(new_n382), .ZN(new_n391));
  INV_X1    g190(.A(G22gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n389), .B(KEYINPUT87), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n382), .A3(G22gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n346), .B1(new_n273), .B2(new_n274), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT81), .ZN(new_n400));
  XOR2_X1   g199(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n275), .A2(new_n271), .A3(new_n346), .A4(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT81), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n404), .A3(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n346), .A2(new_n309), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n337), .B2(new_n348), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n273), .A2(new_n274), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n406), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND3_X1  g218(.A1(new_n371), .A2(new_n268), .A3(new_n270), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n398), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT79), .B1(new_n421), .B2(new_n408), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n423));
  AOI211_X1 g222(.A(new_n423), .B(new_n407), .C1(new_n420), .C2(new_n398), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT5), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n371), .A2(KEYINPUT3), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n411), .B(new_n426), .C1(new_n364), .C2(new_n365), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n407), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n346), .B(new_n429), .C1(new_n273), .C2(new_n274), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n275), .A2(new_n271), .A3(new_n346), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n432), .B2(new_n401), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n414), .B(new_n419), .C1(new_n425), .C2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT82), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI221_X1 g236(.A(KEYINPUT5), .B1(new_n422), .B2(new_n424), .C1(new_n428), .C2(new_n433), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n438), .A2(KEYINPUT82), .A3(new_n419), .A4(new_n414), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n419), .B1(new_n438), .B2(new_n414), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(KEYINPUT6), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n414), .B1(new_n425), .B2(new_n434), .ZN(new_n443));
  INV_X1    g242(.A(new_n419), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(KEYINPUT6), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT83), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT83), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n443), .A2(new_n447), .A3(KEYINPUT6), .A4(new_n444), .ZN(new_n448));
  AOI22_X1  g247(.A1(new_n440), .A2(new_n442), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G226gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n283), .B2(new_n362), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n450), .B1(new_n233), .B2(new_n255), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n360), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n283), .A2(new_n451), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n233), .B2(new_n255), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n455), .B(new_n372), .C1(new_n451), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G8gat), .B(G36gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n459), .B(G64gat), .ZN(new_n460));
  INV_X1    g259(.A(G92gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n458), .A2(KEYINPUT30), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n463), .B1(new_n462), .B2(new_n458), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n458), .A2(new_n466), .A3(new_n462), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n466), .B1(new_n458), .B2(new_n462), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n465), .B1(new_n470), .B2(KEYINPUT30), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n397), .B1(new_n449), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n458), .A2(new_n462), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(new_n467), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n283), .A2(new_n362), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n453), .B1(new_n476), .B2(new_n450), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT91), .B1(new_n477), .B2(new_n359), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n360), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n480), .B(new_n372), .C1(new_n452), .C2(new_n453), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT37), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n462), .B1(new_n458), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT38), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n454), .A2(KEYINPUT37), .A3(new_n457), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n485), .A2(KEYINPUT38), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n475), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n446), .A2(new_n448), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n443), .A2(new_n444), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n437), .A2(new_n439), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n406), .A2(new_n427), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT88), .B(KEYINPUT39), .Z(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n408), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT39), .B1(new_n421), .B2(new_n408), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n407), .B1(new_n406), .B2(new_n427), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n498), .B(new_n419), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT90), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(KEYINPUT40), .ZN(new_n505));
  OR2_X1    g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n441), .B1(new_n505), .B2(new_n503), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT30), .B1(new_n474), .B2(new_n467), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n506), .B(new_n507), .C1(new_n508), .C2(new_n464), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n390), .A2(new_n396), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n308), .B(new_n472), .C1(new_n495), .C2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n306), .A2(new_n300), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n510), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n508), .A2(new_n464), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n494), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n513), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n397), .B2(new_n514), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n510), .A2(KEYINPUT92), .A3(new_n300), .A4(new_n306), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n513), .B1(new_n490), .B2(new_n493), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n521), .A2(new_n517), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n512), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT93), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G29gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n528), .A2(new_n530), .A3(G36gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(G29gat), .B2(G36gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n527), .A2(new_n534), .A3(KEYINPUT14), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n388), .A2(G43gat), .ZN(new_n537));
  INV_X1    g336(.A(G43gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G50gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT15), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n533), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT94), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n535), .A2(new_n533), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT15), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n538), .A2(G50gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n388), .A2(G43gat), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n531), .A3(new_n540), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n542), .B1(new_n547), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g357(.A1(new_n531), .A2(new_n540), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n559), .A2(new_n544), .A3(new_n546), .A4(new_n551), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n555), .A3(new_n556), .A4(new_n542), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G15gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n392), .ZN(new_n564));
  NAND2_X1  g363(.A1(G15gat), .A2(G22gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G1gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT16), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n564), .A2(new_n567), .A3(new_n565), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(G8gat), .B1(new_n570), .B2(KEYINPUT96), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n569), .B(new_n570), .C1(KEYINPUT96), .C2(G8gat), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n562), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(KEYINPUT97), .ZN(new_n578));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n553), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT97), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n562), .A2(new_n581), .A3(new_n576), .ZN(new_n582));
  NAND4_X1  g381(.A1(new_n578), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n526), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n562), .B2(new_n576), .ZN(new_n586));
  AOI211_X1 g385(.A(KEYINPUT97), .B(new_n575), .C1(new_n558), .C2(new_n561), .ZN(new_n587));
  INV_X1    g386(.A(new_n580), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n589), .A2(KEYINPUT98), .A3(KEYINPUT18), .A4(new_n579), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n575), .A2(new_n553), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n579), .B(KEYINPUT13), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n583), .B2(new_n584), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(G197gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT11), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(new_n206), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT12), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n584), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(KEYINPUT99), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n597), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(new_n596), .A3(new_n591), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n609), .A2(KEYINPUT100), .ZN(new_n610));
  XOR2_X1   g409(.A(G57gat), .B(G64gat), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(KEYINPUT100), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G71gat), .B(G78gat), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n610), .A2(new_n611), .A3(new_n614), .A4(new_n612), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(G127gat), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n616), .A2(new_n617), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n575), .B1(KEYINPUT21), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n621), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  XNOR2_X1  g424(.A(G155gat), .B(G183gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n624), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n352), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n628), .B(new_n630), .Z(new_n631));
  AOI21_X1  g430(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G162gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT102), .B1(KEYINPUT101), .B2(KEYINPUT7), .ZN(new_n635));
  AND2_X1   g434(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n636));
  NAND2_X1  g435(.A1(G85gat), .A2(G92gat), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(G99gat), .B(G106gat), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n637), .ZN(new_n641));
  NAND2_X1  g440(.A1(G99gat), .A2(G106gat), .ZN(new_n642));
  INV_X1    g441(.A(G85gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n642), .B1(new_n643), .B2(new_n461), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n638), .A2(new_n640), .A3(new_n641), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n641), .ZN(new_n646));
  NOR3_X1   g445(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n639), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT103), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n562), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n649), .B(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n553), .ZN(new_n654));
  NAND3_X1  g453(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(G134gat), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(G134gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G190gat), .B(G218gat), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n661), .B1(new_n658), .B2(new_n659), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n634), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n633), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AND4_X1   g468(.A1(new_n525), .A2(new_n608), .A3(new_n631), .A4(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G230gat), .A2(G233gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n671), .B(KEYINPUT106), .Z(new_n672));
  NAND2_X1  g471(.A1(new_n618), .A2(new_n649), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n618), .A2(new_n649), .A3(KEYINPUT104), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n645), .A2(new_n648), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n622), .A2(new_n678), .A3(KEYINPUT105), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n618), .B2(new_n649), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT10), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n677), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n653), .A2(KEYINPUT10), .A3(new_n622), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n672), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G120gat), .B(G148gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT107), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(G176gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(G204gat), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n672), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n677), .A2(new_n682), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n687), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n691), .B1(new_n696), .B2(new_n686), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n670), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n494), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n567), .ZN(G1324gat));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n517), .ZN(new_n703));
  INV_X1    g502(.A(G8gat), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT42), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT108), .B(G8gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT16), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g507(.A(KEYINPUT42), .B(new_n705), .S(new_n708), .Z(G1325gat));
  NOR3_X1   g508(.A1(new_n700), .A2(new_n563), .A3(new_n308), .ZN(new_n710));
  INV_X1    g509(.A(new_n700), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n515), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n710), .B1(new_n563), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n700), .A2(new_n510), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  NOR2_X1   g515(.A1(new_n631), .A2(new_n698), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n668), .ZN(new_n718));
  OR2_X1    g517(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(KEYINPUT109), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n719), .A2(new_n525), .A3(new_n608), .A4(new_n720), .ZN(new_n721));
  AOI211_X1 g520(.A(new_n494), .B(new_n721), .C1(new_n528), .C2(new_n530), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT45), .Z(new_n723));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n525), .A2(new_n724), .A3(new_n668), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n525), .A2(new_n724), .A3(KEYINPUT44), .A4(new_n668), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n727), .A2(new_n608), .A3(new_n717), .A4(new_n728), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n528), .B(new_n530), .C1(new_n729), .C2(new_n494), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n723), .A2(new_n730), .ZN(G1328gat));
  OAI21_X1  g530(.A(G36gat), .B1(new_n729), .B2(new_n517), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n721), .A2(G36gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n471), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT46), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n733), .A2(new_n736), .A3(new_n471), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n732), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT111), .ZN(G1329gat));
  OAI21_X1  g538(.A(G43gat), .B1(new_n729), .B2(new_n308), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n515), .A2(new_n538), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n721), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1330gat));
  OAI21_X1  g543(.A(new_n388), .B1(new_n721), .B2(new_n510), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT48), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n397), .A2(G50gat), .ZN(new_n748));
  OAI221_X1 g547(.A(new_n745), .B1(new_n746), .B2(new_n747), .C1(new_n729), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n747), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n749), .B(new_n750), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n525), .A2(new_n698), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n628), .B(new_n630), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n668), .A2(new_n608), .A3(new_n753), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n449), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g556(.A1(new_n752), .A2(new_n754), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n517), .ZN(new_n759));
  NOR2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  AND2_X1   g559(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n760), .ZN(G1333gat));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764));
  INV_X1    g563(.A(new_n308), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n755), .A2(G71gat), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT113), .ZN(new_n767));
  INV_X1    g566(.A(G71gat), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n758), .B2(new_n514), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n767), .B1(new_n766), .B2(new_n769), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n764), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(new_n772), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(KEYINPUT50), .A3(new_n770), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n755), .A2(new_n397), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n631), .A2(new_n608), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n727), .A2(new_n698), .A3(new_n728), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(G85gat), .B1(new_n780), .B2(new_n494), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n525), .A2(new_n668), .A3(new_n779), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT51), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n525), .A2(KEYINPUT51), .A3(new_n668), .A4(new_n779), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n699), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n786), .A2(new_n643), .A3(new_n449), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n788), .B(new_n789), .ZN(G1336gat));
  OAI21_X1  g589(.A(G92gat), .B1(new_n780), .B2(new_n517), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(KEYINPUT115), .A3(new_n785), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n782), .A2(new_n793), .A3(new_n783), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n517), .A2(G92gat), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n792), .A2(new_n698), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT52), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n786), .B2(new_n795), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n791), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1337gat));
  OAI21_X1  g600(.A(G99gat), .B1(new_n780), .B2(new_n308), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n786), .A2(new_n291), .A3(new_n515), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n804), .B(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n510), .A2(new_n699), .A3(G106gat), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n792), .A2(new_n794), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(KEYINPUT117), .ZN(new_n809));
  OAI21_X1  g608(.A(G106gat), .B1(new_n780), .B2(new_n510), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n792), .A2(new_n811), .A3(new_n794), .A4(new_n807), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n510), .A2(G106gat), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n786), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n810), .A2(new_n816), .A3(KEYINPUT118), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT118), .B1(new_n810), .B2(new_n816), .ZN(new_n818));
  OAI22_X1  g617(.A1(new_n813), .A2(new_n814), .B1(new_n817), .B2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n684), .A2(new_n672), .A3(new_n685), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT54), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n822), .A2(new_n686), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n684), .A2(new_n685), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(new_n693), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n691), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n820), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n692), .B1(new_n686), .B2(new_n825), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(KEYINPUT55), .C1(new_n686), .C2(new_n822), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(new_n695), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n607), .B2(new_n605), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n593), .A2(new_n594), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n578), .A2(new_n580), .A3(new_n582), .ZN(new_n834));
  INV_X1    g633(.A(new_n579), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n601), .ZN(new_n837));
  OR3_X1    g636(.A1(new_n836), .A2(KEYINPUT119), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT119), .B1(new_n836), .B2(new_n837), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n591), .A2(new_n602), .A3(new_n596), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n698), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT120), .B1(new_n832), .B2(new_n842), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n828), .A2(new_n695), .A3(new_n830), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n608), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n840), .A2(new_n698), .A3(new_n841), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n848), .A3(new_n669), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n668), .A2(new_n841), .A3(new_n844), .A4(new_n840), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n753), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n754), .A2(new_n699), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n521), .A2(new_n522), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n854), .A2(new_n449), .A3(new_n517), .A4(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n262), .A3(new_n608), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n631), .B1(new_n849), .B2(new_n850), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n754), .A2(new_n699), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(new_n494), .ZN(new_n862));
  INV_X1    g661(.A(new_n516), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n517), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT121), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n866), .A3(new_n517), .A4(new_n863), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n865), .A2(new_n608), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n858), .B1(new_n868), .B2(new_n262), .ZN(G1340gat));
  NAND3_X1  g668(.A1(new_n857), .A2(new_n260), .A3(new_n698), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n865), .A2(new_n698), .A3(new_n867), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n260), .ZN(G1341gat));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n631), .A3(new_n867), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT69), .B(G127gat), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n753), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n856), .B2(new_n876), .ZN(G1342gat));
  NOR3_X1   g676(.A1(new_n856), .A2(G134gat), .A3(new_n669), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n879), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n865), .A2(new_n668), .A3(new_n867), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n880), .B(new_n881), .C1(new_n882), .C2(new_n256), .ZN(G1343gat));
  NOR3_X1   g682(.A1(new_n765), .A2(new_n494), .A3(new_n471), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n885), .B(new_n397), .C1(new_n859), .C2(new_n860), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n669), .B1(new_n832), .B2(new_n842), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n631), .B1(new_n887), .B2(new_n850), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n860), .B1(new_n888), .B2(KEYINPUT122), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n668), .B1(new_n845), .B2(new_n847), .ZN(new_n890));
  AND4_X1   g689(.A1(new_n668), .A2(new_n841), .A3(new_n840), .A4(new_n844), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n753), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n510), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n884), .B(new_n886), .C1(new_n895), .C2(new_n885), .ZN(new_n896));
  INV_X1    g695(.A(new_n608), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n344), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n397), .B(new_n884), .C1(new_n859), .C2(new_n860), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n310), .A3(new_n608), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n900), .A2(KEYINPUT123), .A3(new_n310), .A4(new_n608), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n898), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(KEYINPUT58), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT124), .B1(new_n896), .B2(new_n897), .ZN(new_n907));
  INV_X1    g706(.A(new_n884), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n853), .B1(new_n892), .B2(new_n893), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n397), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n911), .B2(KEYINPUT57), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n608), .A4(new_n886), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n907), .A2(new_n914), .A3(new_n344), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n901), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n906), .A2(new_n918), .ZN(G1344gat));
  NAND2_X1  g718(.A1(new_n328), .A2(new_n329), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n900), .A2(new_n920), .A3(new_n698), .ZN(new_n921));
  INV_X1    g720(.A(new_n896), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT59), .B(new_n920), .C1(new_n922), .C2(new_n698), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT59), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT57), .B1(new_n861), .B2(new_n510), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n885), .B(new_n397), .C1(new_n888), .C2(new_n860), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n925), .A2(new_n698), .A3(new_n884), .A4(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n921), .B1(new_n923), .B2(new_n928), .ZN(G1345gat));
  AOI21_X1  g728(.A(G155gat), .B1(new_n900), .B2(new_n631), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n753), .A2(new_n316), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n922), .B2(new_n931), .ZN(G1346gat));
  NOR2_X1   g731(.A1(new_n323), .A2(new_n324), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n896), .B2(new_n669), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n668), .B1(new_n324), .B2(new_n323), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n899), .B2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n449), .A2(new_n517), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n863), .B(new_n937), .C1(new_n859), .C2(new_n860), .ZN(new_n938));
  OAI21_X1  g737(.A(G169gat), .B1(new_n938), .B2(new_n897), .ZN(new_n939));
  INV_X1    g738(.A(new_n937), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n852), .B2(new_n853), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n855), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n608), .A2(new_n206), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G1348gat));
  OAI21_X1  g743(.A(new_n207), .B1(new_n942), .B2(new_n699), .ZN(new_n945));
  OR3_X1    g744(.A1(new_n938), .A2(new_n699), .A3(new_n248), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n947), .B(new_n948), .ZN(G1349gat));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n941), .A2(new_n953), .A3(new_n863), .A4(new_n631), .ZN(new_n954));
  OAI21_X1  g753(.A(KEYINPUT126), .B1(new_n938), .B2(new_n753), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(G183gat), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n753), .A2(new_n217), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n855), .A3(new_n957), .ZN(new_n958));
  AOI211_X1 g757(.A(new_n951), .B(new_n952), .C1(new_n956), .C2(new_n958), .ZN(new_n959));
  AND4_X1   g758(.A1(new_n950), .A2(new_n956), .A3(KEYINPUT60), .A4(new_n958), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n959), .A2(new_n960), .ZN(G1350gat));
  NAND3_X1  g760(.A1(new_n941), .A2(new_n863), .A3(new_n668), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n962), .A2(new_n963), .A3(G190gat), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n963), .B1(new_n962), .B2(G190gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n668), .A2(new_n224), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n965), .A2(new_n966), .B1(new_n942), .B2(new_n967), .ZN(G1351gat));
  AND2_X1   g767(.A1(new_n925), .A2(new_n926), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n940), .A2(new_n765), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n608), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G197gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n854), .A2(new_n397), .A3(new_n970), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n897), .A2(G197gat), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(G1352gat));
  NAND3_X1  g774(.A1(new_n969), .A2(new_n698), .A3(new_n970), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(G204gat), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n973), .A2(G204gat), .A3(new_n699), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(G1353gat));
  NAND4_X1  g781(.A1(new_n925), .A2(new_n631), .A3(new_n926), .A4(new_n970), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n631), .A2(new_n352), .ZN(new_n986));
  OAI22_X1  g785(.A1(new_n984), .A2(new_n985), .B1(new_n973), .B2(new_n986), .ZN(G1354gat));
  NAND4_X1  g786(.A1(new_n969), .A2(G218gat), .A3(new_n668), .A4(new_n970), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n353), .B1(new_n973), .B2(new_n669), .ZN(new_n989));
  AND2_X1   g788(.A1(new_n988), .A2(new_n989), .ZN(G1355gat));
endmodule


