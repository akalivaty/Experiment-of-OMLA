//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008;
  INV_X1    g000(.A(KEYINPUT90), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g014(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n217));
  NAND2_X1  g016(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n216), .A2(new_n217), .A3(G148gat), .A4(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n207), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n216), .A2(new_n218), .ZN(new_n222));
  OAI211_X1 g021(.A(KEYINPUT75), .B(new_n211), .C1(new_n222), .C2(new_n210), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n215), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT29), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT73), .B(G197gat), .ZN(new_n226));
  INV_X1    g025(.A(G204gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230));
  INV_X1    g029(.A(G211gat), .ZN(new_n231));
  INV_X1    g030(.A(G218gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n228), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n229), .B1(new_n228), .B2(new_n233), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n225), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n224), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n234), .ZN(new_n241));
  AND2_X1   g040(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n242), .A2(new_n243), .A3(new_n210), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT75), .B1(new_n212), .B2(G148gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n219), .B(new_n220), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G141gat), .B(G148gat), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n207), .B(new_n206), .C1(new_n247), .C2(KEYINPUT2), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n238), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n241), .B1(new_n225), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n203), .B1(new_n239), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n252));
  INV_X1    g051(.A(new_n249), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(KEYINPUT29), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n203), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT3), .B1(new_n241), .B2(new_n225), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n255), .C1(new_n256), .C2(new_n224), .ZN(new_n257));
  NAND2_X1  g056(.A1(G228gat), .A2(G233gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G22gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT31), .B(G50gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  AND3_X1   g060(.A1(new_n251), .A2(new_n257), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n261), .B1(new_n251), .B2(new_n257), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT35), .ZN(new_n264));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G183gat), .A2(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G183gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT27), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT27), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n270), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n268), .B1(new_n274), .B2(KEYINPUT28), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n270), .A2(new_n272), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n273), .ZN(new_n278));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT64), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n283), .B1(KEYINPUT26), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT67), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n275), .B(new_n278), .C1(new_n287), .C2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n292));
  MUX2_X1   g091(.A(G183gat), .B(new_n292), .S(G190gat), .Z(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(KEYINPUT24), .B2(new_n268), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n295), .A2(new_n284), .A3(new_n285), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n298), .A2(new_n283), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n294), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n283), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT66), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT24), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n303), .A2(new_n305), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n302), .B1(new_n293), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n291), .B(new_n301), .C1(new_n311), .C2(new_n300), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n266), .B1(new_n312), .B2(new_n225), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n310), .A2(new_n293), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n302), .A2(KEYINPUT25), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n315), .A2(KEYINPUT25), .B1(new_n316), .B2(new_n294), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n265), .B1(new_n317), .B2(new_n291), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n252), .B1(new_n313), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n312), .A2(new_n266), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT29), .B1(new_n317), .B2(new_n291), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n320), .B(new_n241), .C1(new_n321), .C2(new_n266), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(G8gat), .B(G36gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G64gat), .B(G92gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n319), .A2(new_n326), .A3(new_n322), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(KEYINPUT30), .A3(new_n329), .ZN(new_n330));
  OR3_X1    g129(.A1(new_n323), .A2(KEYINPUT30), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(G227gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT69), .ZN(new_n335));
  INV_X1    g134(.A(G134gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G127gat), .ZN(new_n337));
  INV_X1    g136(.A(G127gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G134gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G113gat), .ZN(new_n342));
  AOI21_X1  g141(.A(KEYINPUT68), .B1(new_n342), .B2(G120gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n342), .A2(G120gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n341), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G120gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G113gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n342), .A2(G120gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n351), .A2(new_n340), .B1(new_n337), .B2(new_n339), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n335), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n348), .B2(G113gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n349), .A3(new_n346), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n337), .A2(new_n339), .ZN(new_n359));
  XNOR2_X1  g158(.A(G113gat), .B(G120gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(KEYINPUT1), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n358), .A2(KEYINPUT69), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n353), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n312), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n317), .A2(new_n291), .B1(new_n353), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n334), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT32), .ZN(new_n367));
  XNOR2_X1  g166(.A(G15gat), .B(G43gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT70), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G71gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n368), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G71gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n370), .A2(new_n374), .A3(G99gat), .ZN(new_n375));
  AOI21_X1  g174(.A(G99gat), .B1(new_n370), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n353), .A2(new_n362), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n378), .A2(new_n291), .A3(new_n317), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n312), .A2(new_n363), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n333), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n367), .B(new_n377), .C1(KEYINPUT33), .C2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n377), .B1(new_n381), .B2(KEYINPUT33), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT32), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n379), .A2(new_n333), .A3(new_n380), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT34), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT34), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n379), .A2(new_n380), .A3(new_n389), .A4(new_n333), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n382), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n382), .B2(new_n386), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n264), .B(new_n332), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n219), .A2(new_n220), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n242), .A2(new_n243), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n245), .B1(new_n396), .B2(G148gat), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n248), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n358), .A2(new_n361), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n249), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n351), .A2(new_n340), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n359), .B1(new_n354), .B2(new_n357), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(KEYINPUT76), .A3(new_n249), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n378), .A2(KEYINPUT4), .A3(new_n224), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n246), .A2(new_n248), .A3(new_n361), .A4(new_n358), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n408), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n416), .A2(KEYINPUT77), .A3(new_n412), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n418), .A3(new_n400), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n411), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n420), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT78), .B1(new_n420), .B2(KEYINPUT5), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n415), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n398), .A2(new_n400), .A3(new_n413), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n224), .A2(new_n353), .A3(new_n362), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n425), .B1(new_n413), .B2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n408), .A2(new_n424), .A3(new_n427), .A4(new_n410), .ZN(new_n428));
  XOR2_X1   g227(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT80), .ZN(new_n430));
  XNOR2_X1  g229(.A(G1gat), .B(G29gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G57gat), .B(G85gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n432), .B(new_n433), .Z(new_n434));
  NAND4_X1  g233(.A1(new_n423), .A2(KEYINPUT81), .A3(new_n428), .A4(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n423), .A2(new_n428), .A3(new_n434), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT81), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n434), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n414), .B1(new_n426), .B2(new_n413), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n403), .B2(new_n407), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n420), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n420), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n443), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n428), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n434), .B1(new_n423), .B2(new_n428), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT84), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n437), .A2(new_n440), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n394), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n453), .A2(KEYINPUT82), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n440), .A2(new_n436), .A3(new_n435), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n262), .A2(new_n263), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT71), .B1(new_n388), .B2(new_n390), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n382), .A2(new_n386), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n382), .B2(new_n386), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n463), .A2(new_n469), .A3(new_n332), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n457), .B1(new_n470), .B2(KEYINPUT35), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n392), .A2(new_n393), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n391), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n383), .A2(new_n385), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n379), .A2(new_n380), .ZN(new_n478));
  AOI221_X4 g277(.A(new_n384), .B1(new_n377), .B2(KEYINPUT33), .C1(new_n478), .C2(new_n334), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n382), .A2(new_n386), .A3(new_n465), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT36), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n474), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n464), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n406), .A2(KEYINPUT76), .A3(new_n249), .ZN(new_n487));
  AOI21_X1  g286(.A(KEYINPUT76), .B1(new_n406), .B2(new_n249), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n427), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n411), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT39), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n417), .A2(new_n419), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(new_n410), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n489), .A2(new_n491), .A3(new_n411), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n494), .A2(new_n434), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n330), .A3(new_n331), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n410), .B1(new_n408), .B2(new_n427), .ZN(new_n500));
  INV_X1    g299(.A(new_n493), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n497), .B(new_n434), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n502), .A2(new_n495), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n423), .A2(new_n428), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n505), .B2(new_n441), .ZN(new_n506));
  AOI211_X1 g305(.A(new_n451), .B(new_n434), .C1(new_n423), .C2(new_n428), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n508), .A3(KEYINPUT85), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n452), .A2(new_n454), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n502), .A2(new_n495), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n512), .A2(new_n331), .A3(new_n330), .A4(new_n498), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n486), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n326), .B1(new_n323), .B2(KEYINPUT37), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT38), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT37), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n319), .A2(new_n518), .A3(new_n322), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n516), .B2(new_n519), .ZN(new_n521));
  INV_X1    g320(.A(new_n329), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n523), .B(new_n456), .C1(new_n462), .C2(new_n511), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n485), .B1(new_n515), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n463), .A2(new_n332), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(new_n486), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n471), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT14), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(G29gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT14), .B(G29gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n530), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT86), .B(G43gat), .Z(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT87), .B(G50gat), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n534), .A2(G50gat), .B1(new_n535), .B2(G43gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(G43gat), .A2(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(G43gat), .A2(G50gat), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g340(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n532), .A2(new_n530), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n543), .B2(new_n531), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(G1gat), .B2(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n542), .A2(new_n553), .A3(new_n544), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n546), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT88), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n542), .A2(new_n544), .ZN(new_n558));
  INV_X1    g357(.A(new_n552), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n545), .A2(KEYINPUT88), .A3(new_n552), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n555), .B(new_n556), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT18), .ZN(new_n565));
  OAI22_X1  g364(.A1(new_n560), .A2(new_n561), .B1(new_n558), .B2(new_n559), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n556), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT18), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G113gat), .B(G141gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G197gat), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT11), .B(G169gat), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(new_n575), .B(KEYINPUT12), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n565), .A2(new_n568), .A3(new_n578), .A4(new_n570), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n202), .B1(new_n528), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT85), .B1(new_n504), .B2(new_n508), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n511), .A2(new_n513), .A3(new_n510), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n524), .B(new_n464), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n527), .A3(new_n484), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(KEYINPUT90), .B(new_n580), .C1(new_n587), .C2(new_n471), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G71gat), .A2(G78gat), .ZN(new_n590));
  OR2_X1    g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT91), .ZN(new_n592));
  XNOR2_X1  g391(.A(G57gat), .B(G64gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n593), .A2(KEYINPUT92), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT9), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n593), .B2(KEYINPUT92), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n590), .B(new_n592), .C1(new_n594), .C2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G57gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT93), .B(G57gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n591), .A2(KEYINPUT94), .A3(new_n590), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n591), .A2(new_n590), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT94), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n602), .A2(new_n596), .A3(new_n603), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G127gat), .B(G155gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n612), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G183gat), .B(G211gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n552), .B1(new_n609), .B2(new_n608), .ZN(new_n618));
  XOR2_X1   g417(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  XNOR2_X1  g426(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n628));
  INV_X1    g427(.A(G85gat), .ZN(new_n629));
  INV_X1    g428(.A(G92gat), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT98), .ZN(new_n632));
  XOR2_X1   g431(.A(G99gat), .B(G106gat), .Z(new_n633));
  AOI21_X1  g432(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(G99gat), .A2(G106gat), .ZN(new_n636));
  AOI22_X1  g435(.A1(KEYINPUT8), .A2(new_n636), .B1(new_n629), .B2(new_n630), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n633), .A2(new_n632), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n634), .B(new_n638), .C1(new_n632), .C2(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n546), .A2(new_n644), .A3(new_n554), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n558), .A2(new_n643), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT99), .ZN(new_n647));
  NAND2_X1  g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n650));
  AND3_X1   g449(.A1(new_n646), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n647), .B1(new_n646), .B2(new_n650), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n645), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n649), .A2(KEYINPUT41), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT96), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n655), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n645), .B(new_n657), .C1(new_n651), .C2(new_n652), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n627), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(new_n658), .A3(new_n627), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n624), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G230gat), .ZN(new_n664));
  INV_X1    g463(.A(G233gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n608), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n643), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT10), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n641), .A2(new_n608), .A3(new_n642), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n643), .A2(KEYINPUT10), .A3(new_n667), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n666), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(new_n670), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n666), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G120gat), .B(G148gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT100), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n681), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n676), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n663), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n589), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n463), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g491(.A1(new_n688), .A2(new_n332), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n693), .A2(new_n551), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  INV_X1    g497(.A(G15gat), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n484), .B(KEYINPUT102), .Z(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n688), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n688), .B2(new_n472), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n702), .B1(new_n704), .B2(new_n705), .ZN(G1326gat));
  NOR2_X1   g505(.A1(new_n688), .A2(new_n464), .ZN(new_n707));
  XOR2_X1   g506(.A(KEYINPUT43), .B(G22gat), .Z(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1327gat));
  INV_X1    g508(.A(new_n624), .ZN(new_n710));
  INV_X1    g509(.A(new_n685), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n662), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n713), .B1(new_n582), .B2(new_n588), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(G29gat), .A3(new_n463), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n716), .A2(KEYINPUT45), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n580), .ZN(new_n718));
  INV_X1    g517(.A(new_n662), .ZN(new_n719));
  INV_X1    g518(.A(new_n457), .ZN(new_n720));
  INV_X1    g519(.A(new_n332), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n437), .A2(new_n440), .A3(new_n459), .A4(new_n460), .ZN(new_n722));
  AOI211_X1 g521(.A(new_n721), .B(new_n468), .C1(new_n722), .C2(new_n456), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT35), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n719), .B1(new_n586), .B2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT44), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(KEYINPUT44), .C1(new_n528), .C2(new_n719), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n471), .A2(KEYINPUT104), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n471), .A2(KEYINPUT104), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n586), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n735));
  INV_X1    g534(.A(new_n661), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n736), .B2(new_n659), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n660), .A2(KEYINPUT105), .A3(new_n661), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n718), .B1(new_n731), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G29gat), .B1(new_n744), .B2(new_n463), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n716), .A2(KEYINPUT45), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n717), .A2(new_n745), .A3(new_n746), .ZN(G1328gat));
  NOR3_X1   g546(.A1(new_n715), .A2(G36gat), .A3(new_n332), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G36gat), .B1(new_n744), .B2(new_n332), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n749), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(G1329gat));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n754));
  INV_X1    g553(.A(new_n472), .ZN(new_n755));
  AND2_X1   g554(.A1(new_n755), .A2(new_n534), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n714), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n534), .B1(new_n743), .B2(new_n700), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g559(.A(KEYINPUT106), .B(new_n534), .C1(new_n743), .C2(new_n700), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n754), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n754), .B1(new_n714), .B2(new_n756), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n728), .A2(new_n730), .B1(new_n734), .B2(new_n741), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n764), .A2(new_n484), .A3(new_n718), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n765), .B2(new_n534), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT107), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT107), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n763), .B(new_n768), .C1(new_n765), .C2(new_n534), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n762), .A2(new_n770), .ZN(G1330gat));
  INV_X1    g570(.A(new_n535), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n714), .B2(new_n486), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(KEYINPUT48), .ZN(new_n775));
  OR2_X1    g574(.A1(new_n774), .A2(KEYINPUT48), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n743), .A2(new_n486), .A3(new_n772), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1331gat));
  INV_X1    g579(.A(new_n734), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n663), .A2(new_n581), .A3(new_n711), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n690), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(new_n601), .ZN(G1332gat));
  NOR3_X1   g584(.A1(new_n781), .A2(new_n332), .A3(new_n782), .ZN(new_n786));
  NOR2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  AND2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(G1333gat));
  NAND3_X1  g589(.A1(new_n783), .A2(new_n373), .A3(new_n755), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n781), .A2(new_n701), .A3(new_n782), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n373), .ZN(new_n793));
  XOR2_X1   g592(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n783), .A2(new_n486), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g596(.A1(new_n710), .A2(new_n580), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n711), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT110), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n764), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(KEYINPUT111), .B1(new_n802), .B2(new_n463), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G85gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n802), .A2(KEYINPUT111), .A3(new_n463), .ZN(new_n805));
  INV_X1    g604(.A(new_n798), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n719), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n734), .A2(new_n807), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n690), .A2(new_n629), .A3(new_n711), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n804), .A2(new_n805), .B1(new_n811), .B2(new_n812), .ZN(G1336gat));
  AOI21_X1  g612(.A(new_n630), .B1(new_n801), .B2(new_n721), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n734), .A2(KEYINPUT112), .A3(new_n807), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT51), .B1(new_n815), .B2(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g615(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n817));
  AOI22_X1  g616(.A1(new_n734), .A2(new_n807), .B1(KEYINPUT112), .B2(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n685), .A2(G92gat), .A3(new_n332), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n811), .B2(new_n820), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n814), .B2(new_n824), .ZN(G1337gat));
  OAI21_X1  g624(.A(G99gat), .B1(new_n802), .B2(new_n701), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n685), .A2(G99gat), .A3(new_n472), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n811), .B2(new_n827), .ZN(G1338gat));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n685), .A2(G106gat), .A3(new_n464), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n809), .A2(new_n810), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n801), .A2(new_n832), .A3(new_n486), .ZN(new_n833));
  XOR2_X1   g632(.A(KEYINPUT114), .B(G106gat), .Z(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n832), .B1(new_n801), .B2(new_n486), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n829), .B(new_n831), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n834), .B1(new_n801), .B2(new_n486), .ZN(new_n839));
  INV_X1    g638(.A(new_n830), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n816), .A2(new_n818), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n838), .A2(new_n842), .ZN(G1339gat));
  NOR2_X1   g642(.A1(new_n686), .A2(new_n580), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n671), .A2(new_n672), .A3(new_n666), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n673), .A3(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(KEYINPUT54), .B(new_n666), .C1(new_n671), .C2(new_n672), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n849), .A2(new_n850), .A3(new_n683), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n673), .A2(new_n846), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT116), .B1(new_n852), .B2(new_n681), .ZN(new_n853));
  OAI211_X1 g652(.A(KEYINPUT55), .B(new_n848), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n684), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n850), .B1(new_n849), .B2(new_n683), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(KEYINPUT116), .A3(new_n681), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n847), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(KEYINPUT55), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n560), .A2(new_n561), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n556), .B1(new_n861), .B2(new_n555), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n566), .A2(new_n567), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n575), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n579), .A2(KEYINPUT117), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n579), .A2(new_n864), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n860), .A2(new_n739), .A3(new_n865), .A4(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n866), .A2(new_n685), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n870), .B1(new_n860), .B2(new_n580), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n869), .B1(new_n871), .B2(new_n739), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n844), .B1(new_n872), .B2(new_n624), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n463), .A3(new_n468), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n332), .ZN(new_n875));
  AOI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n580), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n690), .A2(new_n332), .A3(new_n755), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n873), .A2(new_n486), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n581), .A2(new_n342), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(G1340gat));
  AOI21_X1  g679(.A(G120gat), .B1(new_n875), .B2(new_n711), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n685), .A2(new_n348), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n881), .B1(new_n878), .B2(new_n882), .ZN(G1341gat));
  AOI21_X1  g682(.A(new_n338), .B1(new_n878), .B2(new_n710), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n624), .A2(G127gat), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n875), .B2(new_n885), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT118), .Z(G1342gat));
  NAND2_X1  g686(.A1(new_n662), .A2(new_n332), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n888), .B(KEYINPUT119), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n889), .A2(G134gat), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n874), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT56), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n336), .B1(new_n878), .B2(new_n662), .ZN(new_n898));
  XOR2_X1   g697(.A(new_n898), .B(KEYINPUT121), .Z(new_n899));
  NAND3_X1  g698(.A1(new_n893), .A2(KEYINPUT56), .A3(new_n894), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  NOR2_X1   g700(.A1(new_n873), .A2(new_n463), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n700), .A2(new_n464), .ZN(new_n903));
  AND3_X1   g702(.A1(new_n902), .A2(new_n332), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n212), .A3(new_n580), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n869), .B1(new_n871), .B2(new_n662), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n844), .B1(new_n906), .B2(new_n624), .ZN(new_n907));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n907), .B2(new_n464), .ZN(new_n908));
  INV_X1    g707(.A(new_n684), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n858), .B2(KEYINPUT55), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT55), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n868), .A2(new_n910), .A3(new_n913), .A4(new_n865), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n740), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n580), .A3(new_n913), .ZN(new_n916));
  INV_X1    g715(.A(new_n870), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n739), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n624), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n687), .A2(new_n581), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n486), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n485), .A2(new_n463), .A3(new_n721), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n222), .B1(new_n925), .B2(new_n581), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n905), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n927), .B(new_n928), .ZN(G1344gat));
  NOR3_X1   g728(.A1(new_n925), .A2(KEYINPUT59), .A3(new_n685), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n904), .A2(new_n711), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT59), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(new_n210), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n914), .A2(new_n719), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n662), .B1(new_n916), .B2(new_n917), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n624), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n464), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n937), .A2(KEYINPUT123), .A3(KEYINPUT57), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n921), .A2(KEYINPUT57), .A3(new_n486), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT123), .B1(new_n937), .B2(KEYINPUT57), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(new_n711), .A3(new_n924), .ZN(new_n942));
  NAND2_X1  g741(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n933), .B1(new_n942), .B2(new_n943), .ZN(G1345gat));
  NAND3_X1  g743(.A1(new_n904), .A2(new_n204), .A3(new_n710), .ZN(new_n945));
  OAI21_X1  g744(.A(G155gat), .B1(new_n925), .B2(new_n624), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1346gat));
  OAI21_X1  g746(.A(G162gat), .B1(new_n925), .B2(new_n740), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n889), .A2(G162gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n902), .A2(new_n903), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n873), .A2(new_n486), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n690), .A2(new_n332), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n954), .A2(new_n472), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g755(.A(G169gat), .B1(new_n956), .B2(new_n581), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n468), .A2(new_n332), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n960), .B1(new_n873), .B2(new_n690), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n921), .A2(KEYINPUT124), .A3(new_n463), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n580), .A2(new_n284), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT125), .ZN(G1348gat));
  OAI21_X1  g766(.A(G176gat), .B1(new_n956), .B2(new_n685), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n711), .A2(new_n285), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n964), .B2(new_n969), .ZN(G1349gat));
  OAI21_X1  g769(.A(G183gat), .B1(new_n956), .B2(new_n624), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n710), .A2(new_n276), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n963), .A2(KEYINPUT126), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT126), .B1(new_n963), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(KEYINPUT60), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT60), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n977), .B(new_n971), .C1(new_n973), .C2(new_n974), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1350gat));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n273), .A3(new_n739), .ZN(new_n980));
  OAI21_X1  g779(.A(G190gat), .B1(new_n956), .B2(new_n719), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(G1351gat));
  NOR2_X1   g783(.A1(new_n700), .A2(new_n954), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n941), .A2(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(G197gat), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n986), .A2(new_n987), .A3(new_n581), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n961), .A2(new_n962), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n700), .A2(new_n464), .A3(new_n332), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n989), .A2(KEYINPUT127), .A3(new_n990), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n993), .A2(new_n580), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n988), .B1(new_n995), .B2(new_n987), .ZN(G1352gat));
  OAI21_X1  g795(.A(G204gat), .B1(new_n986), .B2(new_n685), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n711), .A2(new_n227), .ZN(new_n998));
  OAI21_X1  g797(.A(KEYINPUT62), .B1(new_n991), .B2(new_n998), .ZN(new_n999));
  OR3_X1    g798(.A1(new_n991), .A2(KEYINPUT62), .A3(new_n998), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(G1353gat));
  NAND4_X1  g800(.A1(new_n993), .A2(new_n231), .A3(new_n710), .A4(new_n994), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n941), .A2(new_n710), .A3(new_n985), .ZN(new_n1003));
  AND3_X1   g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1004));
  AOI21_X1  g803(.A(KEYINPUT63), .B1(new_n1003), .B2(G211gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1354gat));
  OAI21_X1  g805(.A(G218gat), .B1(new_n986), .B2(new_n719), .ZN(new_n1007));
  NAND4_X1  g806(.A1(new_n993), .A2(new_n232), .A3(new_n739), .A4(new_n994), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(G1355gat));
endmodule


