//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT75), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT27), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n190), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G116), .ZN(new_n196));
  INV_X1    g010(.A(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT69), .A3(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n197), .A2(G119), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT2), .B(G113), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n200), .B1(new_n196), .B2(new_n198), .ZN(new_n205));
  INV_X1    g019(.A(new_n203), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT70), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT70), .B1(new_n205), .B2(new_n206), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G143), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n215), .A2(new_n216), .B1(KEYINPUT1), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n220));
  AOI21_X1  g034(.A(KEYINPUT67), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND4_X1   g035(.A1(KEYINPUT67), .A2(new_n220), .A3(new_n212), .A4(new_n214), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G134), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n226), .A2(G134), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G131), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  OAI22_X1  g048(.A1(KEYINPUT64), .A2(new_n233), .B1(new_n234), .B2(G137), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT65), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n236), .B1(new_n226), .B2(G134), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n234), .A2(KEYINPUT65), .A3(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n233), .A2(KEYINPUT64), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n227), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n239), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n232), .B1(new_n244), .B2(new_n231), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT71), .B(new_n218), .C1(new_n221), .C2(new_n222), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n225), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI22_X1  g061(.A1(KEYINPUT65), .A2(new_n229), .B1(new_n227), .B2(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n241), .A2(new_n242), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n228), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(new_n250), .A3(new_n231), .A4(new_n237), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n239), .B2(new_n243), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT66), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n254), .B(G131), .C1(new_n239), .C2(new_n243), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n219), .A2(KEYINPUT0), .A3(G128), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G128), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n219), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n253), .A2(new_n255), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n247), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n210), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n247), .A2(new_n260), .A3(KEYINPUT73), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT28), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n245), .A2(new_n223), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n210), .ZN(new_n269));
  INV_X1    g083(.A(new_n210), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n247), .A2(new_n260), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n266), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n193), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n275), .B(new_n193), .C1(new_n265), .C2(new_n272), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n247), .A2(new_n260), .A3(KEYINPUT30), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT72), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n247), .A2(new_n260), .A3(new_n279), .A4(KEYINPUT30), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n268), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n268), .A2(new_n282), .A3(new_n283), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n281), .B(new_n210), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(new_n192), .A3(new_n271), .ZN(new_n288));
  AOI22_X1  g102(.A1(new_n274), .A2(new_n276), .B1(new_n288), .B2(KEYINPUT31), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n287), .A2(new_n290), .A3(new_n192), .A4(new_n271), .ZN(new_n291));
  AOI21_X1  g105(.A(G902), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G472), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT32), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n274), .A2(new_n276), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n288), .A2(KEYINPUT31), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT32), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n298), .A2(G472), .A3(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n261), .A2(new_n210), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n266), .B1(new_n301), .B2(new_n271), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n265), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n193), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(new_n265), .A2(new_n272), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n304), .B1(new_n307), .B2(new_n193), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n192), .B1(new_n287), .B2(new_n271), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G472), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n300), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n187), .B1(new_n294), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G902), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n297), .A2(new_n293), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n298), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n297), .A2(new_n299), .B1(new_n310), .B2(G472), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(KEYINPUT75), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT22), .B(G137), .ZN(new_n320));
  INV_X1    g134(.A(G953), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n321), .A2(G221), .A3(G234), .ZN(new_n322));
  XOR2_X1   g136(.A(new_n320), .B(new_n322), .Z(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT16), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  OR3_X1    g140(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n211), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n325), .A2(G146), .A3(new_n327), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT23), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n195), .B2(G128), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n333), .B(new_n334), .C1(G119), .C2(new_n216), .ZN(new_n335));
  XNOR2_X1  g149(.A(G119), .B(G128), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  AOI22_X1  g151(.A1(new_n335), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n331), .A2(new_n338), .ZN(new_n339));
  OAI22_X1  g153(.A1(new_n335), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n324), .A2(new_n211), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n330), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n343), .A2(KEYINPUT76), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n339), .B2(new_n342), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n323), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n323), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n348), .B1(new_n343), .B2(KEYINPUT76), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT25), .B1(new_n350), .B2(G902), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n347), .A2(new_n352), .A3(new_n314), .A4(new_n349), .ZN(new_n353));
  INV_X1    g167(.A(G217), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n354), .B1(G234), .B2(new_n314), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n351), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n350), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n350), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT77), .A3(new_n358), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n356), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G221), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT9), .B(G234), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n365), .B1(new_n367), .B2(new_n314), .ZN(new_n368));
  INV_X1    g182(.A(G469), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(new_n314), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT12), .ZN(new_n371));
  INV_X1    g185(.A(G104), .ZN(new_n372));
  OAI21_X1  g186(.A(KEYINPUT3), .B1(new_n372), .B2(G107), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  INV_X1    g188(.A(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(G104), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n372), .A2(G107), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n373), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(KEYINPUT78), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n375), .A2(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n378), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n381), .A2(new_n382), .B1(G101), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(new_n223), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n379), .B(KEYINPUT78), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n223), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT80), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT80), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n385), .A2(new_n392), .A3(new_n223), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n386), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n253), .A2(new_n255), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n371), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n392), .B1(new_n385), .B2(new_n223), .ZN(new_n397));
  AND4_X1   g211(.A1(new_n392), .A2(new_n387), .A3(new_n223), .A4(new_n388), .ZN(new_n398));
  OAI22_X1  g212(.A1(new_n397), .A2(new_n398), .B1(new_n223), .B2(new_n385), .ZN(new_n399));
  INV_X1    g213(.A(new_n395), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(KEYINPUT12), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT10), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n397), .B2(new_n398), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n385), .A2(new_n225), .A3(KEYINPUT10), .A4(new_n246), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n373), .A2(new_n376), .A3(new_n378), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(G101), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n259), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n406), .B2(G101), .ZN(new_n411));
  INV_X1    g225(.A(new_n382), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n410), .B(new_n411), .C1(new_n412), .C2(new_n380), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n410), .B1(new_n387), .B2(new_n411), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n409), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n404), .A2(new_n395), .A3(new_n405), .A4(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G110), .B(G140), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n321), .A2(G227), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n402), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(new_n405), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT10), .B1(new_n391), .B2(new_n393), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n400), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n420), .ZN(new_n427));
  AOI21_X1  g241(.A(G902), .B1(new_n422), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n370), .B1(new_n428), .B2(new_n369), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n421), .B1(new_n402), .B2(new_n417), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n417), .A3(new_n421), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT81), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n423), .A2(new_n424), .ZN(new_n435));
  AOI22_X1  g249(.A1(new_n401), .A2(new_n396), .B1(new_n435), .B2(new_n395), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n431), .C1(new_n436), .C2(new_n421), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n437), .A3(G469), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n368), .B1(new_n429), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n216), .A2(G143), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n213), .A2(G128), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n234), .ZN(new_n444));
  OAI21_X1  g258(.A(G134), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT88), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT88), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n444), .A2(new_n448), .A3(new_n445), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n375), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  XNOR2_X1  g266(.A(G116), .B(G122), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n447), .A2(new_n449), .A3(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n443), .A2(new_n234), .B1(G107), .B2(new_n453), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n441), .A2(KEYINPUT13), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n457), .A2(new_n458), .A3(new_n442), .ZN(new_n459));
  OAI221_X1 g273(.A(new_n456), .B1(G107), .B2(new_n453), .C1(new_n459), .C2(new_n234), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n366), .A2(new_n354), .A3(G953), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(new_n314), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT89), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(KEYINPUT15), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(KEYINPUT15), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n467), .B(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(G113), .B(G122), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(new_n372), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n478));
  AOI21_X1  g292(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n231), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n331), .B1(KEYINPUT17), .B2(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n478), .A2(new_n479), .A3(G131), .ZN(new_n483));
  OR3_X1    g297(.A1(new_n481), .A2(KEYINPUT17), .A3(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n480), .B1(new_n486), .B2(new_n231), .ZN(new_n487));
  OAI211_X1 g301(.A(KEYINPUT18), .B(G131), .C1(new_n478), .C2(new_n479), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n324), .B(new_n211), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n477), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT20), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT19), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  XOR2_X1   g309(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n496));
  MUX2_X1   g310(.A(new_n495), .B(new_n496), .S(new_n324), .Z(new_n497));
  OAI221_X1 g311(.A(new_n330), .B1(new_n481), .B2(new_n483), .C1(new_n497), .C2(G146), .ZN(new_n498));
  INV_X1    g312(.A(new_n477), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n498), .A2(new_n499), .A3(new_n490), .ZN(new_n500));
  NOR2_X1   g314(.A1(G475), .A2(G902), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n492), .A2(new_n493), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n491), .B1(new_n482), .B2(new_n484), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n500), .B(new_n501), .C1(new_n503), .C2(new_n499), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT20), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(G234), .A2(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(G952), .A3(new_n321), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT90), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT21), .B(G898), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(G902), .A3(G953), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n503), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n503), .B2(new_n516), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G475), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n475), .A2(new_n506), .A3(new_n515), .A4(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G214), .B1(G237), .B2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G110), .B(G122), .ZN(new_n523));
  XOR2_X1   g337(.A(KEYINPUT82), .B(KEYINPUT5), .Z(new_n524));
  OR2_X1    g338(.A1(new_n202), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G113), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n524), .B2(new_n200), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n528), .B1(new_n202), .B2(new_n203), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n525), .A2(new_n527), .B1(new_n529), .B2(new_n207), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n385), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n414), .A2(new_n415), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n210), .A2(new_n408), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n523), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n256), .B(G125), .C1(new_n219), .C2(new_n257), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n326), .B2(new_n223), .ZN(new_n537));
  INV_X1    g351(.A(G224), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G953), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT83), .B(KEYINPUT7), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(KEYINPUT84), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n223), .A2(new_n326), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n539), .A3(new_n535), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n535), .A3(new_n540), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT84), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(new_n523), .B(KEYINPUT8), .Z(new_n548));
  INV_X1    g362(.A(KEYINPUT5), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n527), .B1(new_n549), .B2(new_n202), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n208), .B2(new_n209), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n548), .B1(new_n551), .B2(new_n385), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n530), .A2(new_n389), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n539), .B1(new_n542), .B2(new_n535), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n552), .A2(new_n553), .B1(new_n554), .B2(KEYINPUT7), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n534), .A2(new_n547), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n314), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT85), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n523), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n387), .A2(new_n411), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(KEYINPUT79), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n533), .B1(new_n562), .B2(new_n413), .ZN(new_n563));
  INV_X1    g377(.A(new_n531), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(KEYINPUT6), .A3(new_n534), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT6), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(new_n560), .C1(new_n563), .C2(new_n564), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n537), .B(new_n539), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n556), .A2(KEYINPUT85), .A3(new_n314), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n559), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G210), .B1(G237), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n559), .A2(new_n570), .A3(new_n573), .A4(new_n571), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n522), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n440), .A2(new_n520), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n319), .A2(new_n364), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(KEYINPUT91), .B(G101), .Z(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(G3));
  NAND2_X1  g396(.A1(new_n297), .A2(new_n314), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n315), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n585), .A2(new_n440), .A3(new_n363), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT92), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n577), .A2(new_n515), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n468), .A2(new_n314), .ZN(new_n589));
  INV_X1    g403(.A(new_n467), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(new_n468), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT33), .B1(new_n462), .B2(KEYINPUT93), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n466), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n592), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n464), .B2(new_n465), .ZN(new_n595));
  OAI21_X1  g409(.A(G478), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n506), .A2(new_n519), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n588), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n587), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT94), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G6));
  INV_X1    g418(.A(KEYINPUT95), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n502), .A2(new_n505), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n504), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(new_n519), .A3(new_n474), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n588), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n587), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT35), .B(G107), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  AOI211_X1 g427(.A(new_n368), .B(new_n520), .C1(new_n429), .C2(new_n438), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n575), .A2(new_n576), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n343), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n358), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n356), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n615), .A2(new_n521), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n614), .A2(new_n620), .A3(new_n315), .A4(new_n584), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT37), .B(G110), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G12));
  INV_X1    g437(.A(G900), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n510), .B1(new_n624), .B2(new_n513), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n518), .B2(G475), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n606), .A2(new_n626), .A3(new_n474), .A4(new_n607), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT96), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n577), .A2(new_n619), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n316), .A2(KEYINPUT75), .A3(new_n317), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT75), .B1(new_n316), .B2(new_n317), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n439), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  XOR2_X1   g449(.A(new_n625), .B(KEYINPUT39), .Z(new_n636));
  NAND2_X1  g450(.A1(new_n439), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT40), .ZN(new_n638));
  OR2_X1    g452(.A1(new_n638), .A2(KEYINPUT98), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(KEYINPUT98), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n287), .A2(new_n271), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n192), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n301), .A2(new_n271), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(G902), .B1(new_n644), .B2(new_n193), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n293), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n297), .B2(new_n299), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n316), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n619), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n615), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n598), .A2(new_n474), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n522), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n639), .A2(new_n640), .A3(new_n650), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  INV_X1    g470(.A(new_n625), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n597), .A2(new_n598), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n630), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n439), .B(new_n659), .C1(new_n632), .C2(new_n633), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G146), .ZN(G48));
  NAND2_X1  g475(.A1(new_n422), .A2(new_n427), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n314), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT99), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n369), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n428), .B1(new_n664), .B2(new_n369), .ZN(new_n667));
  INV_X1    g481(.A(new_n368), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n666), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n588), .A2(new_n669), .A3(new_n599), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n364), .B(new_n670), .C1(new_n632), .C2(new_n633), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT100), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n363), .B1(new_n313), .B2(new_n318), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT100), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT41), .B(G113), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G15));
  NOR3_X1   g492(.A1(new_n588), .A2(new_n669), .A3(new_n609), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n364), .B(new_n679), .C1(new_n632), .C2(new_n633), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G116), .ZN(G18));
  INV_X1    g495(.A(new_n619), .ZN(new_n682));
  NOR4_X1   g496(.A1(new_n578), .A2(new_n669), .A3(new_n520), .A4(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n632), .B2(new_n633), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT101), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT101), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n319), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT102), .B(G119), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G21));
  OAI21_X1  g504(.A(KEYINPUT105), .B1(new_n292), .B2(new_n293), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n583), .A2(new_n692), .A3(G472), .ZN(new_n693));
  NOR2_X1   g507(.A1(G472), .A2(G902), .ZN(new_n694));
  INV_X1    g508(.A(new_n302), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n263), .A2(new_n264), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n695), .B(new_n696), .C1(new_n697), .C2(KEYINPUT28), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT103), .B1(new_n265), .B2(new_n302), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n699), .A3(new_n193), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n296), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT104), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n296), .A2(new_n700), .A3(KEYINPUT104), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n703), .A2(new_n291), .A3(new_n704), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n691), .A2(new_n693), .B1(new_n694), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n669), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n363), .B(KEYINPUT106), .Z(new_n708));
  NOR3_X1   g522(.A1(new_n578), .A2(new_n514), .A3(new_n653), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND2_X1  g525(.A1(new_n707), .A2(new_n577), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n658), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n706), .A2(new_n713), .A3(new_n619), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n431), .B1(new_n436), .B2(new_n421), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n429), .B1(new_n369), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n668), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n575), .A2(new_n521), .A3(new_n576), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n364), .B(new_n722), .C1(new_n632), .C2(new_n633), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n717), .B1(new_n723), .B2(new_n658), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n720), .A2(new_n658), .A3(new_n721), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n300), .B(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n316), .A3(new_n311), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n726), .A2(new_n708), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n724), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G131), .ZN(G33));
  NAND3_X1  g546(.A1(new_n673), .A2(new_n628), .A3(new_n722), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(new_n370), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n433), .B2(new_n437), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n718), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  OR2_X1    g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n739), .A2(new_n740), .B1(new_n369), .B2(new_n428), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n368), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n636), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n598), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n597), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT43), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n749), .A3(new_n597), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n585), .A2(new_n619), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n721), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n745), .B(new_n754), .C1(new_n753), .C2(new_n752), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n741), .A2(new_n742), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n368), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n743), .A2(KEYINPUT47), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR4_X1   g575(.A1(new_n319), .A2(new_n364), .A3(new_n658), .A4(new_n721), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT108), .B(G140), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G42));
  NOR2_X1   g579(.A1(G952), .A2(G953), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n680), .A2(new_n710), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n676), .A2(new_n688), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n721), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n475), .A2(new_n626), .ZN(new_n772));
  AND4_X1   g586(.A1(new_n608), .A2(new_n771), .A3(new_n619), .A4(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(new_n773), .B(new_n439), .C1(new_n632), .C2(new_n633), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n725), .A2(new_n706), .A3(new_n619), .ZN(new_n775));
  AND2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n598), .A2(new_n474), .ZN(new_n777));
  AOI22_X1  g591(.A1(new_n506), .A2(new_n519), .B1(new_n591), .B2(new_n596), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n577), .A2(new_n515), .A3(new_n779), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n368), .B(new_n363), .C1(new_n429), .C2(new_n438), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n315), .A4(new_n584), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n621), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n673), .B2(new_n579), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n784), .A3(new_n733), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n673), .A2(new_n714), .A3(new_n722), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n729), .A2(new_n708), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n786), .A2(new_n717), .B1(new_n787), .B2(new_n726), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n770), .A2(new_n785), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT52), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n634), .A2(new_n715), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n440), .B1(new_n313), .B2(new_n318), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n577), .A2(new_n598), .A3(new_n474), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n720), .A2(new_n794), .A3(new_n625), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n793), .A2(new_n659), .B1(new_n650), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n791), .B1(new_n792), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n648), .A3(new_n682), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n634), .A2(new_n660), .A3(new_n715), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n790), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n792), .A2(new_n796), .A3(new_n791), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT52), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n789), .A2(new_n801), .A3(KEYINPUT53), .A4(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n799), .A2(KEYINPUT111), .A3(new_n790), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n790), .B1(new_n799), .B2(KEYINPUT111), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n774), .B(new_n775), .C1(new_n723), .C2(new_n629), .ZN(new_n810));
  INV_X1    g624(.A(new_n783), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n580), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n768), .B1(new_n687), .B2(new_n685), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n676), .A4(new_n731), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n806), .B1(new_n809), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n767), .B1(new_n805), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n809), .A2(new_n815), .A3(new_n806), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n789), .A2(new_n801), .A3(new_n804), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n818), .B1(new_n806), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n817), .B1(new_n820), .B2(new_n767), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n691), .A2(new_n693), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n705), .A2(new_n694), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n708), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n669), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n652), .A2(new_n510), .A3(new_n522), .A4(new_n751), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n827), .A3(KEYINPUT50), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n830), .B2(new_n826), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT114), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n828), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  NOR4_X1   g649(.A1(new_n669), .A2(new_n721), .A3(new_n363), .A4(new_n509), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n597), .A2(new_n598), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n649), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n748), .A2(new_n510), .A3(new_n750), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n669), .A3(new_n721), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n706), .A2(new_n619), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT115), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n706), .A2(new_n844), .A3(new_n841), .A4(new_n619), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n839), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n833), .A2(new_n835), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n833), .A2(new_n849), .A3(new_n835), .A4(new_n846), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n666), .A2(new_n667), .ZN(new_n851));
  OR2_X1    g665(.A1(new_n851), .A2(KEYINPUT113), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(KEYINPUT113), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n852), .A2(new_n368), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n759), .A2(new_n760), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n824), .A2(new_n721), .A3(new_n840), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n848), .A2(new_n850), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT120), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n787), .B2(new_n841), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT48), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n787), .A2(new_n861), .A3(new_n841), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n864), .A2(KEYINPUT48), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n863), .A2(new_n865), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n321), .A2(G952), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT119), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n649), .A2(new_n836), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n599), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n824), .A2(new_n712), .A3(new_n840), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n866), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n862), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n868), .B(new_n874), .C1(new_n876), .C2(new_n865), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n879), .B(new_n839), .C1(new_n843), .C2(new_n845), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n857), .A2(KEYINPUT51), .A3(new_n832), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n878), .A2(new_n880), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n857), .A2(KEYINPUT51), .A3(new_n832), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT118), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n877), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n860), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n766), .B1(new_n821), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n747), .A2(new_n368), .A3(new_n522), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n708), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(KEYINPUT49), .B2(new_n851), .ZN(new_n893));
  OR2_X1    g707(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(KEYINPUT109), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT110), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n894), .A2(new_n652), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n648), .ZN(new_n899));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n890), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT122), .ZN(new_n901));
  INV_X1    g715(.A(new_n899), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n860), .A2(new_n888), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n785), .A2(new_n788), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n676), .A2(new_n688), .A3(new_n769), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n804), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT52), .B1(new_n802), .B2(new_n803), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n806), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n789), .B(KEYINPUT53), .C1(new_n808), .C2(new_n807), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n908), .A2(new_n767), .A3(new_n909), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n903), .A2(new_n910), .A3(new_n817), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n901), .B(new_n902), .C1(new_n911), .C2(new_n766), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n900), .A2(new_n912), .ZN(G75));
  NAND2_X1  g727(.A1(new_n566), .A2(new_n568), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(new_n569), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n915), .B(new_n916), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n908), .A2(new_n909), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n918), .A2(G210), .A3(G902), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n917), .B1(new_n919), .B2(KEYINPUT56), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n321), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n919), .A2(KEYINPUT56), .A3(new_n917), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G51));
  XNOR2_X1  g739(.A(new_n918), .B(new_n767), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n370), .B(KEYINPUT57), .Z(new_n927));
  OAI21_X1  g741(.A(new_n662), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n820), .A2(new_n314), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n736), .A2(new_n738), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n921), .B1(new_n928), .B2(new_n931), .ZN(G54));
  NAND2_X1  g746(.A1(new_n492), .A2(new_n500), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(KEYINPUT58), .A2(G475), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n929), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n929), .B2(new_n935), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n936), .A2(new_n937), .A3(new_n921), .ZN(G60));
  NOR2_X1   g752(.A1(new_n593), .A2(new_n595), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n589), .B(KEYINPUT59), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n922), .B1(new_n926), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n821), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n939), .B1(new_n943), .B2(new_n940), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT61), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(G217), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT60), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n908), .B2(new_n909), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n617), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n922), .B1(new_n952), .B2(new_n361), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n946), .B(new_n949), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n951), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n918), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n921), .B1(new_n957), .B2(new_n350), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n952), .A2(new_n617), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n947), .A3(new_n948), .A4(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n955), .A2(new_n960), .ZN(G66));
  OAI21_X1  g775(.A(G953), .B1(new_n511), .B2(new_n538), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n770), .A2(new_n812), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(G953), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n914), .B1(G898), .B2(new_n321), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(G69));
  NAND2_X1  g780(.A1(new_n763), .A2(new_n755), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n578), .A2(new_n653), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n745), .A2(new_n968), .A3(new_n787), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(new_n660), .A3(new_n733), .A4(new_n792), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n967), .A2(new_n970), .A3(new_n788), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n321), .ZN(new_n972));
  INV_X1    g786(.A(new_n284), .ZN(new_n973));
  AOI22_X1  g787(.A1(new_n973), .A2(new_n285), .B1(new_n280), .B2(new_n278), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(new_n497), .Z(new_n975));
  OAI211_X1 g789(.A(new_n972), .B(new_n975), .C1(new_n624), .C2(new_n321), .ZN(new_n976));
  INV_X1    g790(.A(new_n673), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n771), .A2(new_n779), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n977), .A2(new_n637), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n655), .A2(new_n660), .A3(new_n792), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n984));
  AOI211_X1 g798(.A(new_n967), .B(new_n979), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT126), .ZN(new_n987));
  AOI21_X1  g801(.A(G953), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n975), .B(KEYINPUT125), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n976), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n321), .B1(G227), .B2(G900), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n991), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n993), .B(new_n976), .C1(new_n988), .C2(new_n989), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n994), .ZN(G72));
  NAND3_X1  g809(.A1(new_n985), .A2(new_n963), .A3(new_n987), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT63), .Z(new_n998));
  AOI21_X1  g812(.A(new_n642), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n998), .ZN(new_n1000));
  INV_X1    g814(.A(new_n309), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n288), .ZN(new_n1002));
  AOI211_X1 g816(.A(new_n1000), .B(new_n1002), .C1(new_n805), .C2(new_n816), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1000), .B1(new_n971), .B2(new_n963), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n287), .A2(new_n193), .A3(new_n271), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n922), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g820(.A1(new_n999), .A2(new_n1003), .A3(new_n1006), .ZN(G57));
endmodule


