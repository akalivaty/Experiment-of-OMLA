//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(G155gat), .ZN(new_n211));
  INV_X1    g010(.A(G162gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G141gat), .B(G148gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n210), .B(new_n213), .C1(new_n214), .C2(KEYINPUT2), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(KEYINPUT81), .A3(new_n210), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n216), .A2(new_n220), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n228));
  AND2_X1   g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229));
  NOR2_X1   g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n228), .B1(new_n231), .B2(new_n224), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n209), .B(new_n215), .C1(new_n227), .C2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(G155gat), .B2(G162gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n237), .B1(new_n214), .B2(KEYINPUT80), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n238), .A2(new_n216), .A3(new_n226), .A4(new_n220), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n239), .A2(KEYINPUT83), .A3(new_n209), .A4(new_n215), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n235), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n215), .B1(new_n227), .B2(new_n232), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G120gat), .ZN(new_n246));
  INV_X1    g045(.A(G120gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G113gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G134gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(G127gat), .ZN(new_n251));
  INV_X1    g050(.A(G127gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G134gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n249), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n251), .A2(new_n253), .A3(new_n244), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n257), .B1(new_n245), .B2(G120gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n245), .A2(G120gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n247), .A2(KEYINPUT68), .A3(G113gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n249), .A2(new_n254), .B1(new_n256), .B2(new_n261), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT82), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n241), .A2(new_n243), .A3(new_n265), .A4(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n213), .A2(new_n210), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n231), .B2(new_n236), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n216), .A2(new_n220), .A3(new_n226), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(new_n238), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT4), .A3(new_n266), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n274), .B1(new_n242), .B2(new_n263), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n273), .A2(KEYINPUT5), .A3(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n208), .B1(new_n268), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n274), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n266), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(new_n242), .B2(new_n263), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n243), .A2(new_n265), .A3(new_n267), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n282), .B1(new_n241), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n277), .B1(KEYINPUT5), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n267), .A3(new_n242), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT85), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n266), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n265), .A2(new_n267), .A3(KEYINPUT85), .A4(new_n242), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n207), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n288), .A2(new_n289), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n206), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n202), .B1(new_n294), .B2(KEYINPUT6), .ZN(new_n295));
  INV_X1    g094(.A(new_n293), .ZN(new_n296));
  INV_X1    g095(.A(new_n282), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n268), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n291), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n296), .B1(new_n299), .B2(new_n277), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n301));
  NOR4_X1   g100(.A1(new_n300), .A2(KEYINPUT87), .A3(new_n301), .A4(new_n206), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT6), .B1(new_n300), .B2(new_n206), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n206), .B2(new_n300), .ZN(new_n305));
  AND2_X1   g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  INV_X1    g106(.A(G176gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(G169gat), .B2(G176gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT24), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(G190gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT65), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n314), .A2(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n327));
  NAND3_X1  g126(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(KEYINPUT66), .A2(KEYINPUT24), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n319), .A2(new_n320), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND4_X1   g131(.A1(KEYINPUT25), .A2(new_n309), .A3(new_n311), .A4(new_n312), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n322), .A2(new_n324), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n307), .A2(new_n308), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n336), .A3(new_n312), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT26), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(new_n314), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n340));
  AOI21_X1  g139(.A(G190gat), .B1(new_n340), .B2(KEYINPUT27), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT27), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n343));
  AOI21_X1  g142(.A(KEYINPUT28), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT28), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n342), .A2(G183gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n317), .A2(KEYINPUT27), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n339), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n306), .B1(new_n334), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n333), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n316), .A2(new_n319), .A3(new_n320), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n324), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g157(.A1(new_n338), .A2(new_n314), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n337), .B(new_n359), .C1(new_n344), .C2(new_n350), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n353), .B1(new_n361), .B2(new_n306), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND2_X1   g163(.A1(G211gat), .A2(G218gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(G211gat), .A2(G218gat), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT74), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g170(.A1(G211gat), .A2(G218gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT76), .ZN(new_n375));
  AND2_X1   g174(.A1(G197gat), .A2(G204gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(G197gat), .A2(G204gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n377), .A2(new_n379), .B1(new_n380), .B2(new_n372), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n374), .A2(new_n375), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n374), .B2(new_n381), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI22_X1  g184(.A1(new_n378), .A2(new_n376), .B1(new_n365), .B2(KEYINPUT22), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n386), .A2(new_n367), .A3(new_n373), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT75), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n386), .A2(KEYINPUT75), .A3(new_n367), .A4(new_n373), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n385), .A2(new_n391), .A3(KEYINPUT77), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT77), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n389), .A2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n374), .A2(new_n381), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n382), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n393), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n392), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT78), .B1(new_n361), .B2(new_n306), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n364), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n402), .B(KEYINPUT79), .ZN(new_n403));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n398), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n394), .A2(new_n397), .A3(new_n393), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n362), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n401), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n401), .A2(new_n410), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n405), .B1(new_n412), .B2(KEYINPUT37), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n364), .A3(new_n400), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT37), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n399), .B2(new_n362), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT38), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(new_n414), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n401), .B2(new_n410), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT38), .B1(new_n413), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n303), .A2(new_n305), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n406), .B1(new_n401), .B2(new_n410), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT30), .ZN(new_n424));
  NOR3_X1   g223(.A1(new_n411), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n412), .A2(KEYINPUT30), .A3(new_n405), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n288), .A2(new_n289), .A3(new_n207), .A4(new_n290), .ZN(new_n428));
  OAI211_X1 g227(.A(KEYINPUT39), .B(new_n428), .C1(new_n284), .C2(new_n207), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n206), .ZN(new_n431));
  NOR3_X1   g230(.A1(new_n284), .A2(KEYINPUT39), .A3(new_n207), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n294), .B1(new_n433), .B2(KEYINPUT40), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n427), .B(new_n434), .C1(KEYINPUT40), .C2(new_n433), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n241), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n392), .B2(new_n398), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT88), .B1(new_n383), .B2(new_n384), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n396), .A2(new_n441), .A3(new_n382), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n442), .A3(new_n387), .ZN(new_n443));
  AOI21_X1  g242(.A(KEYINPUT3), .B1(new_n443), .B2(new_n437), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n439), .B1(new_n444), .B2(new_n272), .ZN(new_n445));
  AND2_X1   g244(.A1(G228gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n437), .B1(new_n385), .B2(new_n391), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n209), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(new_n242), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n445), .A2(new_n447), .B1(new_n450), .B2(new_n439), .ZN(new_n451));
  INV_X1    g250(.A(G22gat), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n436), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G78gat), .B(G106gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT31), .B(G50gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n445), .A2(new_n447), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n450), .A2(new_n439), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n458), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n452), .B1(new_n458), .B2(new_n459), .ZN(new_n461));
  OAI22_X1  g260(.A1(new_n453), .A2(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n459), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(G22gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n451), .A2(new_n452), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n464), .A2(new_n436), .A3(new_n465), .A4(new_n456), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n422), .A2(new_n435), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT86), .B1(new_n300), .B2(new_n206), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n268), .A2(new_n276), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n207), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT5), .B1(new_n268), .B2(new_n297), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n293), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT86), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(new_n474), .A3(new_n431), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n469), .A2(new_n304), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n294), .A2(new_n202), .A3(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n431), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT87), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n425), .A2(new_n426), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n462), .A2(new_n466), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT36), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n309), .A2(new_n311), .A3(KEYINPUT25), .A4(new_n312), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n486), .B1(new_n331), .B2(new_n330), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n323), .B1(new_n313), .B2(new_n321), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n360), .B(new_n266), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT69), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n358), .A2(KEYINPUT69), .A3(new_n266), .A4(new_n360), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n263), .B1(new_n334), .B2(new_n352), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT71), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT71), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n499), .A3(new_n496), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n495), .A2(KEYINPUT34), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n504));
  INV_X1    g303(.A(new_n492), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT32), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT33), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G15gat), .B(G43gat), .Z(new_n510));
  XNOR2_X1  g309(.A(G71gat), .B(G99gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n512), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n506), .B(KEYINPUT32), .C1(new_n508), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n498), .A2(new_n501), .A3(new_n517), .A4(new_n500), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n503), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n516), .B1(new_n518), .B2(new_n503), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n485), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n516), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n495), .A2(KEYINPUT34), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n523), .B1(KEYINPUT71), .B2(new_n497), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n517), .B1(new_n524), .B2(new_n500), .ZN(new_n525));
  INV_X1    g324(.A(new_n518), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT73), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n528), .A3(new_n518), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n522), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT36), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n521), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n468), .A2(new_n484), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT35), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n301), .B1(new_n473), .B2(new_n431), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n479), .B(new_n477), .C1(new_n537), .C2(new_n294), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n536), .A2(new_n538), .A3(new_n481), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n535), .B1(new_n539), .B2(new_n483), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n427), .B1(new_n303), .B2(new_n476), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n520), .B1(new_n462), .B2(new_n466), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n503), .A2(new_n528), .A3(new_n518), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n528), .B1(new_n503), .B2(new_n518), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n516), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT35), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n534), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G15gat), .B(G22gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT16), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n549), .B1(new_n550), .B2(G1gat), .ZN(new_n551));
  NAND2_X1  g350(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n551), .B(new_n552), .C1(G1gat), .C2(new_n549), .ZN(new_n553));
  NOR2_X1   g352(.A1(KEYINPUT93), .A2(G8gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT14), .ZN(new_n559));
  INV_X1    g358(.A(G29gat), .ZN(new_n560));
  INV_X1    g359(.A(G36gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT15), .ZN(new_n565));
  INV_X1    g364(.A(G43gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G50gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n567), .B2(KEYINPUT92), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n558), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G43gat), .B(G50gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n563), .ZN(new_n572));
  NOR3_X1   g371(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n556), .A2(new_n557), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT91), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  OAI22_X1  g374(.A1(new_n572), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI22_X1  g375(.A1(new_n569), .A2(new_n571), .B1(new_n565), .B2(new_n576), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n558), .A2(new_n568), .A3(new_n570), .A4(new_n564), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n555), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n577), .A2(KEYINPUT17), .A3(new_n578), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT17), .B1(new_n577), .B2(new_n578), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n555), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT18), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n555), .A2(KEYINPUT94), .A3(new_n579), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n555), .A2(new_n579), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT94), .B1(new_n555), .B2(new_n579), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n584), .B(KEYINPUT13), .Z(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n586), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n587), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G197gat), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT11), .B(G169gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT90), .B(KEYINPUT12), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n593), .A3(new_n601), .A4(new_n594), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n548), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608));
  OR2_X1    g407(.A1(G99gat), .A2(G106gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT100), .B(G92gat), .ZN(new_n613));
  INV_X1    g412(.A(G85gat), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n613), .A2(new_n614), .B1(KEYINPUT8), .B2(new_n610), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT99), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(G85gat), .A3(G92gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT7), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT7), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n616), .A2(new_n619), .A3(G85gat), .A4(G92gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI211_X1 g420(.A(new_n608), .B(new_n612), .C1(new_n615), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n611), .A2(KEYINPUT101), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n609), .A2(new_n608), .A3(new_n610), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n615), .A2(new_n623), .A3(new_n621), .A4(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(KEYINPUT102), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n615), .A2(new_n621), .A3(new_n624), .ZN(new_n628));
  INV_X1    g427(.A(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n631), .A3(new_n625), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n627), .B(new_n632), .C1(new_n581), .C2(new_n582), .ZN(new_n633));
  INV_X1    g432(.A(new_n579), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n625), .ZN(new_n635));
  NAND2_X1  g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n636), .B(KEYINPUT97), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n634), .A2(new_n635), .B1(KEYINPUT41), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n633), .B2(new_n639), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(KEYINPUT103), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n633), .A2(new_n639), .A3(new_n645), .A4(new_n641), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT98), .ZN(new_n649));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n647), .A2(KEYINPUT104), .A3(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n659));
  XNOR2_X1  g458(.A(G57gat), .B(G64gat), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n659), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G71gat), .B(G78gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT21), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g465(.A(G127gat), .B(G155gat), .Z(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n555), .B1(new_n665), .B2(new_n664), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(G231gat), .A2(G233gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT96), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G183gat), .B(G211gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n670), .B(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n643), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n651), .A2(new_n678), .A3(new_n642), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n657), .A2(new_n658), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(KEYINPUT104), .B1(new_n647), .B2(new_n652), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n654), .B(new_n651), .C1(new_n644), .C2(new_n646), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n677), .B(new_n679), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT105), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(G230gat), .A2(G233gat), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n662), .B(new_n663), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n635), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT10), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n664), .A2(new_n630), .A3(new_n625), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n635), .A2(new_n688), .A3(KEYINPUT10), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n687), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n689), .A2(new_n691), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n687), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n695), .A2(new_n697), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n685), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n607), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n480), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G1gat), .ZN(G1324gat));
  INV_X1    g510(.A(G8gat), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n712), .B1(new_n708), .B2(new_n427), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT16), .B(G8gat), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n707), .A2(new_n481), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT42), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(KEYINPUT42), .B2(new_n715), .ZN(G1325gat));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n521), .B(new_n718), .C1(new_n530), .C2(new_n532), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n520), .A2(new_n485), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n545), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(new_n521), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(G15gat), .B1(new_n707), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n536), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(G15gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n707), .B2(new_n727), .ZN(G1326gat));
  OR3_X1    g527(.A1(new_n707), .A2(KEYINPUT107), .A3(new_n467), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT107), .B1(new_n707), .B2(new_n467), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(KEYINPUT43), .B(G22gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1327gat));
  NAND2_X1  g532(.A1(new_n657), .A2(new_n679), .ZN(new_n734));
  INV_X1    g533(.A(new_n677), .ZN(new_n735));
  INV_X1    g534(.A(new_n705), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT108), .ZN(new_n738));
  AND2_X1   g537(.A1(new_n607), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(new_n560), .A3(new_n709), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT45), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n468), .A2(new_n484), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n547), .B1(new_n724), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n734), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n742), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n534), .B2(new_n547), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n705), .B(KEYINPUT109), .Z(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(new_n606), .A3(new_n677), .ZN(new_n751));
  NAND4_X1  g550(.A1(new_n746), .A2(new_n747), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n533), .A2(KEYINPUT106), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n753), .A2(new_n484), .A3(new_n468), .A4(new_n719), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n467), .A2(new_n545), .A3(new_n531), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n480), .A2(KEYINPUT35), .A3(new_n481), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n467), .A2(new_n536), .A3(new_n481), .A4(new_n538), .ZN(new_n757));
  AOI22_X1  g556(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n535), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n745), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n749), .B(new_n751), .C1(new_n759), .C2(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT110), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n752), .A2(new_n709), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n741), .B1(new_n560), .B2(new_n762), .ZN(G1328gat));
  NAND3_X1  g562(.A1(new_n752), .A2(new_n427), .A3(new_n761), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(G36gat), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n607), .A2(new_n561), .A3(new_n427), .A4(new_n738), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n765), .A2(new_n768), .A3(KEYINPUT111), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(G1329gat));
  NOR2_X1   g572(.A1(new_n726), .A2(G43gat), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n739), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(G43gat), .B1(new_n760), .B2(new_n724), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(KEYINPUT47), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n724), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n752), .A2(new_n778), .A3(new_n761), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n779), .A2(G43gat), .B1(new_n739), .B2(new_n774), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n777), .B1(new_n780), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g580(.A1(new_n467), .A2(G50gat), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n739), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(G50gat), .B1(new_n760), .B2(new_n467), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n739), .A2(KEYINPUT112), .A3(new_n782), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n785), .A2(KEYINPUT48), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n752), .A2(new_n483), .A3(new_n761), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n789), .A2(G50gat), .B1(new_n739), .B2(new_n782), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n790), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g590(.A1(new_n754), .A2(new_n758), .ZN(new_n792));
  INV_X1    g591(.A(new_n750), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n685), .A2(new_n605), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n709), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g597(.A1(new_n795), .A2(new_n481), .ZN(new_n799));
  NOR2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  AND2_X1   g599(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n802), .B1(new_n799), .B2(new_n800), .ZN(G1333gat));
  INV_X1    g602(.A(G71gat), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n795), .A2(new_n804), .A3(new_n724), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT113), .ZN(new_n806));
  XOR2_X1   g605(.A(new_n536), .B(KEYINPUT114), .Z(new_n807));
  NOR2_X1   g606(.A1(new_n795), .A2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n808), .A2(KEYINPUT115), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n804), .B1(new_n808), .B2(KEYINPUT115), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT50), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n806), .B(new_n813), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1334gat));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n483), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G78gat), .ZN(G1335gat));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n605), .A2(new_n677), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n746), .A2(new_n705), .A3(new_n749), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n820), .B2(new_n480), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G85gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n820), .A2(new_n818), .A3(new_n480), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n759), .A2(new_n819), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(KEYINPUT51), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(KEYINPUT51), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n709), .A2(new_n614), .A3(new_n705), .ZN(new_n828));
  OAI22_X1  g627(.A1(new_n822), .A2(new_n823), .B1(new_n827), .B2(new_n828), .ZN(G1336gat));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n830));
  INV_X1    g629(.A(new_n613), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n820), .B2(new_n481), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n793), .A2(G92gat), .A3(new_n481), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n827), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OAI221_X1 g637(.A(new_n832), .B1(new_n833), .B2(new_n830), .C1(new_n827), .C2(new_n836), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1337gat));
  OAI21_X1  g639(.A(G99gat), .B1(new_n820), .B2(new_n724), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n726), .A2(G99gat), .A3(new_n736), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n827), .B2(new_n842), .ZN(G1338gat));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  OAI21_X1  g643(.A(G106gat), .B1(new_n820), .B2(new_n467), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n793), .A2(G106gat), .A3(new_n467), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n827), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  OAI221_X1 g650(.A(new_n845), .B1(new_n846), .B2(new_n844), .C1(new_n827), .C2(new_n849), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(G1339gat));
  NOR2_X1   g652(.A1(new_n480), .A2(new_n427), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n680), .A2(new_n684), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n856), .A2(new_n857), .A3(new_n606), .A4(new_n736), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n680), .A2(new_n684), .A3(new_n606), .A4(new_n736), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n591), .A2(new_n592), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n584), .B1(new_n580), .B2(new_n583), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n599), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n604), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n705), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT122), .B1(new_n736), .B2(new_n865), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n692), .A2(new_n693), .A3(new_n687), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n692), .A2(KEYINPUT120), .A3(new_n693), .A4(new_n687), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n694), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n701), .B1(new_n694), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(KEYINPUT55), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n704), .ZN(new_n882));
  AOI21_X1  g681(.A(KEYINPUT55), .B1(new_n878), .B2(new_n880), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n605), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n734), .B1(new_n870), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n734), .A2(new_n884), .A3(new_n866), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n735), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n855), .B1(new_n861), .B2(new_n889), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n890), .A2(new_n755), .ZN(new_n891));
  AOI21_X1  g690(.A(G113gat), .B1(new_n891), .B2(new_n605), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n861), .A2(new_n889), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n467), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(new_n726), .A3(new_n855), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n606), .A2(new_n245), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(G1340gat));
  AOI21_X1  g696(.A(G120gat), .B1(new_n891), .B2(new_n705), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n793), .A2(new_n247), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n895), .B2(new_n899), .ZN(G1341gat));
  NAND3_X1  g699(.A1(new_n891), .A2(new_n252), .A3(new_n677), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n895), .A2(new_n677), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n252), .ZN(G1342gat));
  NAND3_X1  g702(.A1(new_n891), .A2(new_n250), .A3(new_n734), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(KEYINPUT56), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n895), .A2(new_n734), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n905), .B(new_n906), .C1(new_n250), .C2(new_n907), .ZN(G1343gat));
  OAI21_X1  g707(.A(KEYINPUT123), .B1(new_n882), .B2(new_n883), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n878), .A2(new_n880), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT55), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT123), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n912), .A2(new_n913), .A3(new_n704), .A4(new_n881), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n909), .A2(new_n914), .A3(new_n605), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n866), .A2(new_n705), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n745), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n677), .B1(new_n918), .B2(new_n887), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n860), .B2(new_n858), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT57), .B1(new_n920), .B2(new_n467), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n467), .B1(new_n861), .B2(new_n889), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT57), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n778), .A2(new_n855), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n606), .A2(new_n221), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n921), .A2(new_n924), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  NOR2_X1   g726(.A1(KEYINPUT124), .A2(KEYINPUT58), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n778), .A2(new_n467), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n890), .A2(new_n605), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n930), .B2(new_n221), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(KEYINPUT124), .A2(KEYINPUT58), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n932), .B(new_n933), .ZN(G1344gat));
  NAND2_X1  g733(.A1(new_n890), .A2(new_n929), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n936), .A2(new_n222), .A3(new_n705), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n467), .A2(KEYINPUT57), .ZN(new_n940));
  INV_X1    g739(.A(new_n859), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n919), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n705), .A3(new_n925), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n938), .B1(new_n945), .B2(G148gat), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n938), .A2(G148gat), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n705), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n937), .B1(new_n946), .B2(new_n949), .ZN(G1345gat));
  NAND3_X1  g749(.A1(new_n936), .A2(new_n211), .A3(new_n677), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n948), .A2(new_n677), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n211), .ZN(G1346gat));
  AOI21_X1  g752(.A(G162gat), .B1(new_n936), .B2(new_n734), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n745), .A2(new_n212), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n948), .B2(new_n955), .ZN(G1347gat));
  NOR2_X1   g755(.A1(new_n709), .A2(new_n481), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n893), .A2(new_n755), .A3(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(G169gat), .B1(new_n959), .B2(new_n605), .ZN(new_n960));
  INV_X1    g759(.A(new_n957), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n807), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n894), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n606), .A2(new_n307), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1348gat));
  NAND3_X1  g764(.A1(new_n959), .A2(new_n308), .A3(new_n705), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n894), .A2(new_n793), .A3(new_n962), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n966), .B1(new_n967), .B2(new_n308), .ZN(G1349gat));
  NAND4_X1  g767(.A1(new_n959), .A2(new_n348), .A3(new_n349), .A4(new_n677), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n894), .A2(new_n735), .A3(new_n962), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n317), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n959), .A2(new_n318), .A3(new_n734), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n963), .A2(new_n734), .ZN(new_n974));
  XNOR2_X1  g773(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n974), .A2(G190gat), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n974), .B2(G190gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(G1351gat));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(new_n939), .B2(new_n943), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n778), .A2(new_n961), .ZN(new_n981));
  OAI211_X1 g780(.A(new_n942), .B(KEYINPUT126), .C1(new_n922), .C2(new_n923), .ZN(new_n982));
  INV_X1    g781(.A(G197gat), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n606), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n922), .A2(new_n981), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n983), .B1(new_n986), .B2(new_n606), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n985), .A2(new_n987), .ZN(G1352gat));
  NOR3_X1   g787(.A1(new_n986), .A2(G204gat), .A3(new_n736), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT62), .ZN(new_n990));
  AND4_X1   g789(.A1(new_n750), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n991));
  INV_X1    g790(.A(G204gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(G1353gat));
  NOR3_X1   g792(.A1(new_n778), .A2(new_n735), .A3(new_n961), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n922), .A2(new_n368), .A3(new_n994), .ZN(new_n995));
  OAI211_X1 g794(.A(new_n942), .B(new_n994), .C1(new_n922), .C2(new_n923), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n995), .B(KEYINPUT127), .C1(new_n997), .C2(new_n998), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(G1354gat));
  NOR2_X1   g802(.A1(new_n745), .A2(new_n369), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n369), .B1(new_n986), .B2(new_n745), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1355gat));
endmodule


