//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n213), .B1(new_n203), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n212), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  NOR2_X1   g0022(.A1(new_n212), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n225));
  XNOR2_X1  g0025(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n206), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n210), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n226), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT13), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT3), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(G226), .ZN(new_n257));
  OR2_X1    g0057(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n258), .B(new_n259), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(new_n255), .B(new_n256), .C1(new_n257), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  INV_X1    g0066(.A(G45), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(G1), .A3(G13), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n270), .A3(G274), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n271), .B1(new_n214), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n249), .B1(new_n265), .B2(new_n275), .ZN(new_n276));
  AOI211_X1 g0076(.A(KEYINPUT13), .B(new_n274), .C1(new_n263), .C2(new_n264), .ZN(new_n277));
  OAI21_X1  g0077(.A(G169), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT14), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n265), .A2(new_n275), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n265), .A2(new_n249), .A3(new_n275), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(G179), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT14), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n284), .B(G169), .C1(new_n276), .C2(new_n277), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n279), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G50), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT74), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n288), .B(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n251), .A2(G20), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n291), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n229), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT11), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(KEYINPUT11), .A3(new_n295), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  OR3_X1    g0102(.A1(new_n302), .A2(KEYINPUT12), .A3(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n295), .B1(new_n209), .B2(G20), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n303), .A2(new_n304), .B1(G68), .B2(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n298), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n286), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT8), .B(G58), .ZN(new_n310));
  INV_X1    g0110(.A(new_n287), .ZN(new_n311));
  INV_X1    g0111(.A(G77), .ZN(new_n312));
  OAI22_X1  g0112(.A1(new_n310), .A2(new_n311), .B1(new_n210), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  INV_X1    g0114(.A(new_n291), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n295), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n305), .A2(G77), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(G77), .C2(new_n302), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n252), .B2(new_n253), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G238), .ZN(new_n325));
  INV_X1    g0125(.A(G232), .ZN(new_n326));
  INV_X1    g0126(.A(G107), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G107), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n325), .B1(new_n262), .B2(new_n326), .C1(new_n254), .C2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(new_n264), .ZN(new_n334));
  INV_X1    g0134(.A(G244), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n271), .B1(new_n335), .B2(new_n273), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n321), .B(new_n322), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  OR2_X1    g0139(.A1(new_n334), .A2(new_n336), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n340), .A2(G179), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n319), .B1(new_n337), .B2(G169), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT71), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n281), .A2(G190), .A3(new_n282), .ZN(new_n350));
  OAI21_X1  g0150(.A(G200), .B1(new_n276), .B2(new_n277), .ZN(new_n351));
  AND3_X1   g0151(.A1(new_n350), .A2(new_n351), .A3(new_n307), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT71), .B1(new_n343), .B2(new_n346), .ZN(new_n354));
  AND4_X1   g0154(.A1(new_n309), .A2(new_n349), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT68), .ZN(new_n357));
  MUX2_X1   g0157(.A(new_n356), .B(new_n310), .S(new_n357), .Z(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n305), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n359), .B1(new_n358), .B2(new_n302), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT76), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n260), .A2(new_n261), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT7), .B1(new_n362), .B2(new_n210), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n252), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n253), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G58), .A2(G68), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n204), .A2(new_n205), .A3(new_n367), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT16), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n361), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI211_X1 g0172(.A(KEYINPUT76), .B(KEYINPUT16), .C1(new_n366), .C2(new_n369), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n295), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(G20), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n287), .A2(G159), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT75), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n364), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n254), .B2(G20), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n362), .A2(KEYINPUT75), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n384), .B2(G68), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n375), .B1(new_n385), .B2(KEYINPUT16), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n360), .B1(new_n374), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  OAI211_X1 g0188(.A(G226), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  INV_X1    g0190(.A(G223), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n389), .B(new_n390), .C1(new_n262), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n264), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n270), .A2(G232), .A3(new_n272), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n271), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n388), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G179), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n398), .B(new_n395), .C1(new_n392), .C2(new_n264), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n387), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n203), .B1(new_n382), .B2(new_n364), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n371), .B1(new_n402), .B2(new_n378), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT76), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n384), .A2(G68), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(KEYINPUT16), .A3(new_n369), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n361), .B(new_n371), .C1(new_n402), .C2(new_n378), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n295), .A4(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n360), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n400), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT18), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n395), .B1(new_n392), .B2(new_n264), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n414), .A2(G190), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n338), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n408), .A2(new_n417), .A3(KEYINPUT17), .A4(new_n409), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n401), .A2(new_n413), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n271), .ZN(new_n424));
  INV_X1    g0224(.A(new_n273), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n424), .B1(G226), .B2(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n324), .A2(G223), .B1(new_n362), .B2(G77), .ZN(new_n427));
  AND2_X1   g0227(.A1(new_n258), .A2(new_n259), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(G222), .A3(new_n254), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n426), .B1(new_n430), .B2(new_n270), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT10), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n302), .A2(G50), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(G50), .B2(new_n305), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n440));
  INV_X1    g0240(.A(G150), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n440), .B1(new_n441), .B2(new_n311), .C1(new_n358), .C2(new_n315), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n442), .B2(new_n295), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT72), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT9), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n443), .B2(KEYINPUT9), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI221_X1 g0248(.A(new_n432), .B1(new_n341), .B2(new_n431), .C1(new_n443), .C2(KEYINPUT9), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n436), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n447), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n445), .ZN(new_n452));
  INV_X1    g0252(.A(new_n449), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n435), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n443), .B1(new_n388), .B2(new_n431), .ZN(new_n456));
  OR2_X1    g0256(.A1(new_n431), .A2(G179), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n355), .A2(new_n423), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n209), .A2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n375), .A2(new_n302), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n314), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n302), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n314), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n291), .A2(G97), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n254), .A2(new_n210), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n203), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT78), .ZN(new_n475));
  NOR2_X1   g0275(.A1(G87), .A2(G97), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n328), .A2(new_n330), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT77), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n478), .A2(new_n479), .A3(new_n210), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n478), .B2(new_n210), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n482), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n484), .A2(KEYINPUT78), .A3(new_n477), .A4(new_n480), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n474), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n295), .B1(new_n486), .B2(KEYINPUT79), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT79), .ZN(new_n488));
  AOI211_X1 g0288(.A(new_n488), .B(new_n474), .C1(new_n483), .C2(new_n485), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n467), .B(new_n469), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n267), .A2(G1), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n216), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n270), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n270), .A2(G274), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n209), .A2(G45), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n254), .A2(G244), .A3(G1698), .ZN(new_n497));
  NAND2_X1  g0297(.A1(G33), .A2(G116), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n497), .B(new_n498), .C1(new_n214), .C2(new_n262), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n496), .B1(new_n499), .B2(new_n264), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(G169), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n398), .B2(new_n500), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n490), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n483), .A2(new_n485), .ZN(new_n504));
  INV_X1    g0304(.A(new_n474), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n488), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n486), .A2(KEYINPUT79), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n507), .A2(new_n295), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n465), .A2(G87), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n499), .A2(new_n264), .ZN(new_n511));
  INV_X1    g0311(.A(new_n496), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n341), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(G200), .B2(new_n500), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n509), .A2(new_n469), .A3(new_n510), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n262), .B2(new_n335), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n324), .A2(G250), .B1(G33), .B2(G283), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n428), .A2(KEYINPUT4), .A3(G244), .A4(new_n254), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n264), .ZN(new_n521));
  INV_X1    g0321(.A(new_n494), .ZN(new_n522));
  OR2_X1    g0322(.A1(KEYINPUT5), .A2(G41), .ZN(new_n523));
  NAND2_X1  g0323(.A1(KEYINPUT5), .A2(G41), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n495), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n491), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n528), .A2(G257), .A3(new_n270), .ZN(new_n529));
  INV_X1    g0329(.A(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n521), .A2(new_n398), .A3(new_n526), .A4(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  INV_X1    g0332(.A(G97), .ZN(new_n533));
  NOR3_X1   g0333(.A1(new_n532), .A2(new_n533), .A3(G107), .ZN(new_n534));
  XNOR2_X1  g0334(.A(G97), .B(G107), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n534), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n536), .A2(new_n210), .B1(new_n312), .B2(new_n311), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n332), .B1(new_n382), .B2(new_n364), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n295), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n468), .A2(new_n533), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n465), .A2(G97), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n526), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n529), .B(new_n543), .C1(new_n520), .C2(new_n264), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n531), .B(new_n542), .C1(new_n544), .C2(G169), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n529), .B1(new_n520), .B2(new_n264), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n547), .A2(G190), .A3(new_n526), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n548), .C1(new_n338), .C2(new_n544), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n503), .A2(new_n515), .A3(new_n545), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(G20), .B1(G33), .B2(G283), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G33), .B2(new_n533), .ZN(new_n552));
  INV_X1    g0352(.A(G116), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G20), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n295), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(KEYINPUT80), .A2(KEYINPUT20), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(KEYINPUT80), .A2(KEYINPUT20), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n552), .A2(new_n295), .A3(new_n554), .A4(new_n556), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n375), .A2(new_n302), .A3(G116), .A4(new_n463), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n468), .A2(new_n553), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(G1698), .C1(new_n260), .C2(new_n261), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n362), .A2(G303), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n254), .A2(G257), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n258), .A2(new_n259), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n264), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n525), .A2(new_n264), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(G270), .B1(new_n522), .B2(new_n525), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n563), .B1(new_n572), .B2(G200), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n341), .B2(new_n572), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(G169), .A3(new_n563), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT21), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n569), .A2(G179), .A3(new_n571), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n563), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n572), .A2(KEYINPUT21), .A3(G169), .A4(new_n563), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n574), .A2(new_n577), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n210), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(KEYINPUT22), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT22), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n254), .A2(new_n584), .A3(new_n210), .A4(G87), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(KEYINPUT23), .B1(new_n331), .B2(new_n210), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(KEYINPUT81), .B(KEYINPUT23), .C1(new_n331), .C2(new_n210), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT23), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n210), .A2(G107), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n591), .A2(new_n592), .B1(new_n291), .B2(G116), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n586), .A2(new_n589), .A3(new_n590), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT24), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n590), .A2(new_n593), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT24), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n586), .A3(new_n597), .A4(new_n589), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n295), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n464), .A2(new_n327), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n301), .A2(new_n592), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT25), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n254), .A2(G257), .A3(G1698), .ZN(new_n605));
  NAND2_X1  g0405(.A1(G33), .A2(G294), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n605), .B(new_n606), .C1(new_n216), .C2(new_n262), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n264), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n528), .A2(G264), .A3(new_n270), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n526), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n608), .A2(new_n610), .A3(G190), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G200), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n600), .A2(new_n604), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n608), .A2(new_n610), .A3(new_n398), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n388), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n375), .B1(new_n595), .B2(new_n598), .ZN(new_n617));
  INV_X1    g0417(.A(new_n604), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n614), .A2(new_n619), .ZN(new_n620));
  NOR4_X1   g0420(.A1(new_n462), .A2(new_n550), .A3(new_n581), .A4(new_n620), .ZN(G372));
  AOI21_X1  g0421(.A(new_n412), .B1(new_n410), .B2(new_n411), .ZN(new_n622));
  AOI211_X1 g0422(.A(KEYINPUT18), .B(new_n400), .C1(new_n408), .C2(new_n409), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n346), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n309), .B1(new_n626), .B2(new_n352), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n420), .A2(new_n421), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n455), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n459), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT82), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n545), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n547), .A2(new_n526), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n388), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(KEYINPUT82), .A3(new_n531), .A4(new_n542), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n503), .A3(new_n637), .A4(new_n515), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n545), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n503), .A2(new_n515), .A3(new_n641), .A4(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n503), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n503), .A2(new_n515), .A3(new_n545), .A4(new_n549), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n609), .A2(new_n526), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n264), .B2(new_n607), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n611), .B1(new_n647), .B2(new_n338), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n617), .A2(new_n648), .A3(new_n618), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n649), .B1(new_n651), .B2(new_n619), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n644), .B1(new_n645), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n643), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n632), .B1(new_n462), .B2(new_n655), .ZN(G369));
  NAND2_X1  g0456(.A1(new_n301), .A2(new_n210), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(KEYINPUT27), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(G213), .A3(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G343), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n662), .A2(new_n563), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n650), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n581), .B2(new_n663), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n665), .A2(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n662), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n667), .B1(new_n600), .B2(new_n604), .ZN(new_n668));
  OAI22_X1  g0468(.A1(new_n620), .A2(new_n668), .B1(new_n619), .B2(new_n667), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n614), .A2(new_n619), .A3(new_n650), .A4(new_n667), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n616), .A2(new_n615), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n600), .B2(new_n604), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n667), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT83), .B1(new_n671), .B2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n671), .A2(KEYINPUT83), .A3(new_n674), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n670), .B1(new_n675), .B2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n223), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n477), .A2(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n227), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT28), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n662), .B1(new_n643), .B2(new_n653), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n578), .A2(new_n500), .A3(new_n547), .A4(new_n647), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n647), .A2(new_n500), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n691), .A2(new_n398), .A3(new_n635), .A4(new_n572), .ZN(new_n692));
  AND3_X1   g0492(.A1(new_n500), .A2(new_n608), .A3(new_n610), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n547), .A4(new_n578), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n690), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n662), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  XOR2_X1   g0497(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(KEYINPUT31), .B2(new_n697), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n620), .A2(new_n581), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n645), .A3(new_n667), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(G330), .B1(new_n701), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n638), .A2(KEYINPUT26), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n503), .A2(new_n515), .A3(new_n641), .A4(new_n639), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n614), .B1(new_n673), .B2(new_n650), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n503), .B1(new_n709), .B2(new_n550), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n667), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n687), .A2(new_n705), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n684), .B1(new_n714), .B2(G1), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT85), .ZN(G364));
  NOR2_X1   g0516(.A1(new_n300), .A2(G20), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n209), .B1(new_n717), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n679), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n666), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(G330), .B2(new_n665), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n223), .A2(new_n254), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n723), .B1(KEYINPUT86), .B2(G355), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(KEYINPUT86), .B2(G355), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G116), .B2(new_n223), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n244), .A2(new_n267), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n223), .A2(new_n362), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n728), .B1(new_n228), .B2(new_n267), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(G13), .A2(G33), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G20), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n229), .B1(G20), .B2(new_n388), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n720), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n338), .A2(G179), .ZN(new_n738));
  XNOR2_X1  g0538(.A(new_n738), .B(KEYINPUT88), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n210), .A2(G190), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT87), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT87), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n327), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n210), .A2(new_n341), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n398), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n202), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n740), .A2(new_n746), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n254), .B1(new_n749), .B2(new_n312), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n744), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n739), .A2(new_n745), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n215), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G179), .A2(G200), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n210), .B1(new_n754), .B2(G190), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n533), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n341), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G50), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n757), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n758), .A2(G190), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n762), .B1(G68), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n741), .A2(new_n742), .A3(new_n754), .ZN(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  OR3_X1    g0566(.A1(new_n765), .A2(KEYINPUT32), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT32), .B1(new_n765), .B2(new_n766), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n764), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n752), .ZN(new_n770));
  INV_X1    g0570(.A(new_n765), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n770), .A2(G303), .B1(new_n771), .B2(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n362), .B1(new_n749), .B2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n747), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G322), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G283), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n772), .B(new_n776), .C1(new_n777), .C2(new_n743), .ZN(new_n778));
  NOR2_X1   g0578(.A1(KEYINPUT33), .A2(G317), .ZN(new_n779));
  AND2_X1   g0579(.A1(KEYINPUT33), .A2(G317), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n763), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G294), .ZN(new_n782));
  INV_X1    g0582(.A(G326), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n781), .B1(new_n782), .B2(new_n755), .C1(new_n783), .C2(new_n760), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n753), .A2(new_n769), .B1(new_n778), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n737), .B1(new_n785), .B2(new_n734), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n733), .B(KEYINPUT89), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n665), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n722), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(G396));
  NAND2_X1  g0590(.A1(new_n347), .A2(new_n667), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n642), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n639), .B2(new_n638), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n792), .B1(new_n794), .B2(new_n710), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n319), .A2(new_n662), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n343), .A2(new_n796), .B1(new_n344), .B2(new_n345), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n346), .A2(new_n667), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n795), .B1(new_n685), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n720), .B1(new_n800), .B2(new_n705), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n705), .B2(new_n800), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n734), .A2(new_n731), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n719), .B(new_n679), .C1(new_n312), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n734), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n743), .A2(new_n215), .B1(new_n752), .B2(new_n327), .ZN(new_n806));
  INV_X1    g0606(.A(new_n763), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n757), .B1(new_n807), .B2(new_n777), .C1(new_n808), .C2(new_n760), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n765), .A2(new_n773), .ZN(new_n810));
  OAI221_X1 g0610(.A(new_n362), .B1(new_n749), .B2(new_n553), .C1(new_n782), .C2(new_n747), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n806), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n749), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G143), .A2(new_n775), .B1(new_n813), .B2(G159), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n814), .B1(new_n807), .B2(new_n441), .C1(new_n815), .C2(new_n760), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT90), .Z(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n770), .A2(G50), .B1(new_n771), .B2(G132), .ZN(new_n819));
  INV_X1    g0619(.A(new_n743), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G68), .ZN(new_n821));
  INV_X1    g0621(.A(new_n755), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n362), .B1(new_n822), .B2(G58), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n824), .B1(new_n817), .B2(KEYINPUT34), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n812), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n804), .B1(new_n805), .B2(new_n826), .C1(new_n799), .C2(new_n732), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n802), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(G384));
  INV_X1    g0629(.A(new_n536), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(KEYINPUT35), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(KEYINPUT35), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n831), .A2(G116), .A3(new_n230), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT36), .Z(new_n834));
  NAND3_X1  g0634(.A1(new_n228), .A2(G77), .A3(new_n367), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n761), .A2(G68), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n209), .B(G13), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT39), .ZN(new_n839));
  INV_X1    g0639(.A(new_n660), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n410), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n422), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n410), .A2(new_n411), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT37), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n844), .A2(new_n841), .A3(new_n845), .A4(new_n418), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n844), .A2(new_n841), .A3(new_n418), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT37), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n843), .A2(KEYINPUT95), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n841), .B1(new_n628), .B2(new_n624), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT95), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT38), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n386), .B1(KEYINPUT16), .B2(new_n385), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n660), .B1(new_n854), .B2(new_n409), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n422), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n854), .A2(new_n409), .B1(new_n400), .B2(new_n660), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n845), .B1(new_n858), .B2(new_n418), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT93), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n418), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n862), .B2(new_n857), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n846), .A3(KEYINPUT93), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n856), .A2(new_n861), .A3(new_n864), .A4(KEYINPUT38), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n839), .B1(new_n853), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n286), .A2(new_n308), .A3(new_n667), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT94), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n856), .A2(new_n861), .A3(new_n864), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n865), .A3(KEYINPUT39), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n867), .A2(new_n869), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT91), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n795), .A2(new_n875), .A3(new_n798), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n791), .B1(new_n643), .B2(new_n653), .ZN(new_n877));
  INV_X1    g0677(.A(new_n798), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT91), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n865), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n307), .A2(new_n667), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n286), .B2(new_n352), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(KEYINPUT92), .ZN(new_n884));
  INV_X1    g0684(.A(new_n882), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n309), .A2(new_n353), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT92), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n887), .B(new_n882), .C1(new_n286), .C2(new_n352), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n880), .A2(new_n881), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n625), .A2(new_n660), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n874), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n462), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n687), .A2(new_n712), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n631), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n892), .B(new_n895), .Z(new_n896));
  AND3_X1   g0696(.A1(new_n695), .A2(KEYINPUT31), .A3(new_n662), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n699), .B1(new_n695), .B2(new_n662), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n703), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n900), .A2(new_n901), .A3(new_n889), .A4(new_n799), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n865), .B2(new_n872), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n799), .A3(new_n889), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n853), .B2(new_n866), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n903), .B1(new_n906), .B2(KEYINPUT40), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n899), .A2(new_n703), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n462), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n881), .A2(new_n905), .A3(new_n901), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n848), .A2(new_n846), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n850), .B2(new_n851), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n843), .A2(KEYINPUT95), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n871), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n904), .B1(new_n914), .B2(new_n865), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n910), .B1(new_n915), .B2(new_n901), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n916), .A2(new_n893), .A3(new_n900), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n909), .A2(new_n917), .A3(G330), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n896), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n209), .B2(new_n717), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n896), .A2(new_n918), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n838), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT96), .Z(G367));
  OAI221_X1 g0723(.A(new_n735), .B1(new_n223), .B2(new_n314), .C1(new_n240), .C2(new_n728), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n720), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT101), .Z(new_n926));
  NAND2_X1  g0726(.A1(new_n770), .A2(G116), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT46), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n771), .A2(G317), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n820), .A2(G97), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n254), .B1(new_n763), .B2(G294), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(G283), .A2(new_n813), .B1(new_n822), .B2(new_n331), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT102), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n775), .A2(G303), .B1(G311), .B2(new_n759), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT103), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n755), .A2(new_n203), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n759), .B2(G143), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n766), .B2(new_n807), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n254), .B1(new_n749), .B2(new_n761), .C1(new_n441), .C2(new_n747), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n770), .B2(G58), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n771), .A2(G137), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n820), .A2(G77), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n932), .A2(new_n937), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT47), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n734), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n503), .A2(new_n515), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n509), .A2(new_n469), .A3(new_n510), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n662), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT97), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n503), .A2(new_n952), .A3(new_n662), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n955), .B1(new_n954), .B2(new_n956), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n926), .B1(new_n948), .B2(new_n950), .C1(new_n960), .C2(new_n787), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT100), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n549), .B(new_n545), .C1(new_n546), .C2(new_n667), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n641), .A2(new_n662), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(KEYINPUT45), .B(new_n965), .C1(new_n676), .C2(new_n675), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n965), .B1(new_n676), .B2(new_n675), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n671), .A2(new_n674), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT83), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n671), .A2(KEYINPUT83), .A3(new_n674), .ZN(new_n973));
  INV_X1    g0773(.A(new_n965), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT44), .A4(new_n974), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n966), .A2(new_n969), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n962), .B1(new_n979), .B2(new_n670), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n969), .A2(new_n966), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n978), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n670), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(KEYINPUT100), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n650), .A2(new_n667), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n671), .B1(new_n669), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(new_n666), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n989), .A2(new_n712), .A3(new_n687), .A4(new_n705), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n979), .A2(new_n670), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n980), .A2(new_n985), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n714), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n679), .B(KEYINPUT41), .Z(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n719), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n670), .A2(new_n974), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n671), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT42), .B1(new_n965), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n965), .A2(new_n1000), .A3(KEYINPUT42), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n545), .B1(new_n963), .B2(new_n619), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n1002), .A2(new_n1003), .B1(new_n667), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n959), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT43), .B1(new_n1006), .B2(new_n957), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT98), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1004), .A2(new_n667), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1003), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n1001), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT43), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n958), .B2(new_n959), .ZN(new_n1014));
  OAI21_X1  g0814(.A(KEYINPUT98), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1009), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT99), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1018), .A2(new_n1014), .A3(new_n1012), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1017), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n999), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT99), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(new_n998), .A3(new_n1020), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n961), .B1(new_n997), .B2(new_n1027), .ZN(G387));
  NOR2_X1   g0828(.A1(new_n237), .A2(new_n267), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n1029), .A2(new_n728), .B1(new_n681), .B2(new_n723), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n310), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g0832(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n681), .A3(new_n1033), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1030), .A2(new_n1034), .B1(new_n327), .B2(new_n678), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n720), .B1(new_n1035), .B2(new_n736), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G317), .A2(new_n775), .B1(new_n813), .B2(G303), .ZN(new_n1037));
  INV_X1    g0837(.A(G322), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n1037), .B1(new_n807), .B2(new_n773), .C1(new_n1038), .C2(new_n760), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT48), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n777), .B2(new_n755), .C1(new_n782), .C2(new_n752), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n1044), .A2(KEYINPUT49), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n362), .B1(new_n765), .B2(new_n783), .C1(new_n743), .C2(new_n553), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(KEYINPUT49), .B2(new_n1044), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n358), .A2(new_n807), .B1(new_n203), .B2(new_n749), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT105), .Z(new_n1050));
  NAND2_X1  g0850(.A1(new_n822), .A2(new_n466), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n362), .B1(new_n775), .B2(G50), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n930), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n752), .A2(new_n312), .B1(new_n765), .B2(new_n441), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n759), .A2(G159), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT104), .Z(new_n1056));
  OR3_X1    g0856(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1048), .B1(new_n1050), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1036), .B1(new_n1058), .B2(new_n734), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n669), .A2(new_n787), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n719), .B2(new_n989), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n714), .A2(new_n989), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n990), .A2(new_n679), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT106), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT106), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1061), .B(new_n1066), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1067), .ZN(G393));
  INV_X1    g0868(.A(new_n993), .ZN(new_n1069));
  AND3_X1   g0869(.A1(new_n981), .A2(new_n982), .A3(new_n670), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n670), .B1(new_n981), .B2(new_n982), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n679), .B1(new_n1072), .B2(new_n991), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT108), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1071), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n992), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n680), .B1(new_n1076), .B2(new_n990), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT108), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1077), .A2(new_n1078), .A3(new_n993), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n974), .A2(new_n733), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n735), .B1(new_n533), .B2(new_n223), .C1(new_n247), .C2(new_n728), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n720), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT107), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n755), .A2(new_n312), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n254), .B1(new_n749), .B2(new_n310), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G50), .C2(new_n763), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n775), .A2(G159), .B1(G150), .B2(new_n759), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT51), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT51), .ZN(new_n1090));
  AND3_X1   g0890(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n820), .A2(G87), .B1(G143), .B2(new_n771), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n203), .C2(new_n752), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n254), .B1(new_n813), .B2(G294), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n1094), .B1(new_n553), .B2(new_n755), .C1(new_n807), .C2(new_n808), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT52), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n759), .A2(G317), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n773), .B2(new_n747), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n744), .B1(G283), .B2(new_n770), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1038), .B2(new_n765), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1093), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1084), .B1(new_n1103), .B2(new_n734), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1072), .A2(new_n719), .B1(new_n1081), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1080), .A2(new_n1105), .ZN(G390));
  INV_X1    g0906(.A(KEYINPUT111), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT109), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n900), .A2(G330), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n889), .A2(new_n799), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n875), .B1(new_n795), .B2(new_n798), .ZN(new_n1112));
  NOR3_X1   g0912(.A1(new_n877), .A2(KEYINPUT91), .A3(new_n878), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n889), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n869), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1114), .A2(new_n1115), .B1(new_n867), .B2(new_n873), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n849), .A2(new_n852), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n866), .B1(new_n1117), .B2(new_n871), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n889), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n667), .B(new_n797), .C1(new_n708), .C2(new_n710), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n798), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1118), .A2(new_n1121), .A3(new_n869), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1108), .B(new_n1111), .C1(new_n1116), .C2(new_n1122), .ZN(new_n1123));
  OR3_X1    g0923(.A1(new_n1118), .A2(new_n869), .A3(new_n1121), .ZN(new_n1124));
  INV_X1    g0924(.A(G330), .ZN(new_n1125));
  MUX2_X1   g0925(.A(new_n698), .B(KEYINPUT31), .S(new_n696), .Z(new_n1126));
  AOI21_X1  g0926(.A(new_n1125), .B1(new_n1126), .B2(new_n703), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n799), .A3(new_n889), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n867), .A2(new_n873), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n869), .B1(new_n880), .B2(new_n889), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1124), .B(new_n1128), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1108), .B1(new_n1133), .B2(new_n1111), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1107), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n867), .A2(new_n873), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1122), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1111), .ZN(new_n1139));
  OAI21_X1  g0939(.A(KEYINPUT109), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1140), .A2(KEYINPUT111), .A3(new_n1131), .A4(new_n1123), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1109), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n893), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n895), .A2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1109), .A2(KEYINPUT110), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n799), .B1(new_n1109), .B2(KEYINPUT110), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1119), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n798), .A3(new_n1120), .A4(new_n1128), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n889), .B1(new_n1127), .B2(new_n799), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n880), .B1(new_n1149), .B2(new_n1111), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1144), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1135), .A2(new_n1141), .A3(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1140), .A2(new_n1151), .A3(new_n1131), .A4(new_n1123), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT112), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1135), .A2(KEYINPUT112), .A3(new_n1141), .A4(new_n1152), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1156), .A2(new_n679), .A3(new_n1157), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1140), .A2(new_n719), .A3(new_n1131), .A4(new_n1123), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n358), .A2(new_n803), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n720), .A2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n820), .A2(G50), .B1(G125), .B2(new_n771), .ZN(new_n1162));
  INV_X1    g0962(.A(G132), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n254), .B1(new_n747), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G128), .B2(new_n759), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1162), .B(new_n1165), .C1(new_n766), .C2(new_n755), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT54), .B(G143), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n813), .A2(new_n1168), .B1(G137), .B2(new_n763), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OR2_X1    g0970(.A1(new_n1170), .A2(KEYINPUT113), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1172));
  NAND3_X1  g0972(.A1(new_n770), .A2(G150), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1172), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n752), .B2(new_n441), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1170), .A2(KEYINPUT113), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1171), .A2(new_n1173), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n821), .B1(new_n215), .B2(new_n752), .C1(new_n782), .C2(new_n765), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n813), .A2(G97), .B1(new_n331), .B2(new_n763), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1180), .A2(KEYINPUT115), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(KEYINPUT115), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n759), .A2(G283), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n254), .B(new_n1085), .C1(G116), .C2(new_n775), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1166), .A2(new_n1177), .B1(new_n1178), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1161), .B1(new_n1186), .B2(new_n734), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1129), .B2(new_n732), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1159), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT116), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1159), .A2(KEYINPUT116), .A3(new_n1188), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1158), .A2(new_n1194), .ZN(G378));
  INV_X1    g0995(.A(new_n1144), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n892), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n443), .A2(new_n660), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n460), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1198), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n455), .A2(new_n459), .A3(new_n1200), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1202), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1200), .B1(new_n455), .B2(new_n459), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n458), .B(new_n1198), .C1(new_n450), .C2(new_n454), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1203), .A2(new_n1207), .A3(KEYINPUT120), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT120), .B1(new_n1203), .B2(new_n1207), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n907), .A2(new_n1210), .A3(new_n1125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n916), .B2(G330), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1197), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1212), .B1(new_n907), .B2(new_n1125), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT120), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1203), .A2(new_n1207), .A3(KEYINPUT120), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n916), .A2(G330), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1216), .A2(new_n1221), .A3(new_n892), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1154), .A2(new_n1196), .B1(new_n1215), .B2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n679), .B1(new_n1223), .B2(KEYINPUT57), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1154), .A2(new_n1196), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1215), .A2(new_n1222), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1225), .A2(KEYINPUT57), .A3(new_n1226), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1216), .A2(new_n892), .A3(new_n1221), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n892), .B1(new_n1216), .B2(new_n1221), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n719), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n803), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n720), .B1(G50), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n820), .A2(G58), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT117), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n938), .B1(new_n763), .B2(G97), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n553), .B2(new_n760), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n362), .A2(new_n266), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n749), .A2(new_n314), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1238), .B(new_n1239), .C1(G107), .C2(new_n775), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1240), .B1(new_n312), .B2(new_n752), .C1(new_n777), .C2(new_n765), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1235), .A2(new_n1237), .A3(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT58), .Z(new_n1243));
  OAI211_X1 g1043(.A(new_n1238), .B(new_n761), .C1(G33), .C2(G41), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n752), .A2(new_n1167), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1246), .A2(KEYINPUT118), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1246), .A2(KEYINPUT118), .ZN(new_n1248));
  INV_X1    g1048(.A(G128), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n747), .A2(new_n1249), .B1(new_n749), .B2(new_n815), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n807), .A2(new_n1163), .B1(new_n755), .B2(new_n441), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(G125), .C2(new_n759), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1247), .A2(new_n1248), .A3(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(KEYINPUT59), .ZN(new_n1255));
  OAI211_X1 g1055(.A(new_n251), .B(new_n266), .C1(new_n743), .C2(new_n766), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(G124), .B2(new_n771), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1243), .B(new_n1244), .C1(new_n1254), .C2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT119), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n805), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1232), .B(new_n1263), .C1(new_n731), .C2(new_n1220), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT121), .B1(new_n1230), .B2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n718), .B1(new_n1215), .B2(new_n1222), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT121), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1264), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1224), .A2(new_n1227), .B1(new_n1266), .B2(new_n1269), .ZN(G375));
  NAND2_X1  g1070(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1119), .A2(new_n731), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n720), .B1(G68), .B2(new_n1231), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n770), .A2(G159), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n1163), .A2(new_n760), .B1(new_n807), .B2(new_n1167), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G50), .B2(new_n822), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n771), .A2(G128), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n254), .B1(new_n749), .B2(new_n441), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(G137), .B2(new_n775), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1274), .A2(new_n1276), .A3(new_n1277), .A4(new_n1279), .ZN(new_n1280));
  OAI221_X1 g1080(.A(new_n1051), .B1(new_n807), .B2(new_n553), .C1(new_n782), .C2(new_n760), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n770), .A2(G97), .B1(new_n771), .B2(G303), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n362), .B1(new_n332), .B2(new_n749), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G283), .B2(new_n775), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n944), .A3(new_n1284), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1235), .A2(new_n1280), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1273), .B1(new_n1286), .B2(new_n734), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1271), .A2(new_n719), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1288));
  XOR2_X1   g1088(.A(new_n995), .B(KEYINPUT122), .Z(new_n1289));
  NAND2_X1  g1089(.A1(new_n1152), .A2(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1271), .A2(new_n1196), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1288), .B1(new_n1290), .B2(new_n1291), .ZN(G381));
  NOR2_X1   g1092(.A1(new_n1269), .A2(new_n1266), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT57), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n680), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1223), .A2(KEYINPUT57), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1293), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n680), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1189), .B1(new_n1299), .B2(new_n1157), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1105), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n828), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1065), .A2(new_n789), .A3(new_n1067), .ZN(new_n1304));
  NOR4_X1   g1104(.A1(new_n1303), .A2(G381), .A3(G387), .A4(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1298), .A2(new_n1300), .A3(new_n1305), .ZN(G407));
  NAND2_X1  g1106(.A1(new_n661), .A2(G213), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1298), .A2(new_n1300), .A3(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(G407), .A2(new_n1309), .A3(G213), .ZN(G409));
  NAND2_X1  g1110(.A1(new_n1152), .A2(KEYINPUT60), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1291), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT60), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1151), .A2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n680), .B1(new_n1315), .B2(new_n1291), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1316), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1317), .A2(G384), .A3(new_n1288), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G384), .B1(new_n1317), .B2(new_n1288), .ZN(new_n1319));
  OAI211_X1 g1119(.A(G2897), .B(new_n1308), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1319), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1317), .A2(G384), .A3(new_n1288), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1308), .A2(G2897), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1189), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1267), .A2(new_n1264), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1289), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1327), .B1(new_n1294), .B2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1158), .A2(new_n1326), .A3(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1193), .B1(new_n1299), .B2(new_n1157), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1330), .B1(new_n1331), .B2(G375), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1325), .B1(new_n1332), .B2(new_n1307), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1332), .A2(new_n1307), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  AOI22_X1  g1136(.A1(KEYINPUT123), .A2(new_n1333), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G387), .A2(new_n1302), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(G387), .A2(new_n1302), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT124), .B1(G387), .B2(new_n1302), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(G393), .A2(G396), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1304), .ZN(new_n1343));
  OAI22_X1  g1143(.A1(new_n1339), .A2(new_n1340), .B1(new_n1341), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  OR2_X1    g1145(.A1(new_n997), .A2(new_n1027), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(G390), .A2(new_n1346), .A3(new_n961), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1343), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1347), .A2(new_n1348), .A3(KEYINPUT124), .A4(new_n1338), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1344), .A2(new_n1345), .A3(new_n1349), .ZN(new_n1350));
  XNOR2_X1  g1150(.A(new_n1350), .B(KEYINPUT125), .ZN(new_n1351));
  AND2_X1   g1151(.A1(new_n1320), .A2(new_n1324), .ZN(new_n1352));
  AOI22_X1  g1152(.A1(new_n1298), .A2(G378), .B1(new_n1300), .B2(new_n1329), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1352), .B1(new_n1353), .B2(new_n1308), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT123), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1351), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1298), .A2(G378), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1308), .B1(new_n1357), .B2(new_n1330), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(KEYINPUT63), .A3(new_n1334), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1337), .A2(new_n1356), .A3(new_n1359), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1344), .A2(KEYINPUT126), .A3(new_n1349), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(KEYINPUT126), .B1(new_n1344), .B2(new_n1349), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT62), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1332), .A2(new_n1365), .A3(new_n1334), .A4(new_n1307), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1354), .A2(new_n1366), .A3(new_n1345), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1365), .B1(new_n1358), .B2(new_n1334), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1364), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1360), .A2(new_n1369), .ZN(G405));
  INV_X1    g1170(.A(new_n1334), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(G375), .A2(new_n1300), .ZN(new_n1372));
  AND3_X1   g1172(.A1(new_n1357), .A2(new_n1371), .A3(new_n1372), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1371), .B1(new_n1357), .B2(new_n1372), .ZN(new_n1374));
  NOR2_X1   g1174(.A1(new_n1373), .A2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(KEYINPUT127), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1376), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1377));
  INV_X1    g1177(.A(new_n1363), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1378), .A2(KEYINPUT127), .A3(new_n1361), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1377), .A2(new_n1379), .ZN(new_n1380));
  XNOR2_X1  g1180(.A(new_n1375), .B(new_n1380), .ZN(G402));
endmodule


