

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  XNOR2_X1 U326 ( .A(n392), .B(n319), .ZN(n320) );
  XNOR2_X1 U327 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U328 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U329 ( .A(n329), .B(n328), .ZN(n331) );
  INV_X1 U330 ( .A(G190GAT), .ZN(n457) );
  XNOR2_X1 U331 ( .A(n334), .B(KEYINPUT64), .ZN(n555) );
  XOR2_X1 U332 ( .A(n455), .B(n454), .Z(n532) );
  XNOR2_X1 U333 ( .A(n457), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(G218GAT), .ZN(n393) );
  XOR2_X1 U336 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n295) );
  XNOR2_X1 U337 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U339 ( .A(n393), .B(n296), .ZN(n300) );
  XOR2_X1 U340 ( .A(G134GAT), .B(G162GAT), .Z(n396) );
  XOR2_X1 U341 ( .A(G92GAT), .B(G85GAT), .Z(n298) );
  XNOR2_X1 U342 ( .A(G99GAT), .B(G106GAT), .ZN(n297) );
  XNOR2_X1 U343 ( .A(n298), .B(n297), .ZN(n312) );
  XNOR2_X1 U344 ( .A(n396), .B(n312), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT11), .B(KEYINPUT79), .Z(n302) );
  NAND2_X1 U347 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n311) );
  XOR2_X1 U350 ( .A(G29GAT), .B(KEYINPUT8), .Z(n306) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(G36GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U353 ( .A(G50GAT), .B(KEYINPUT7), .Z(n307) );
  XOR2_X1 U354 ( .A(n308), .B(n307), .Z(n345) );
  INV_X1 U355 ( .A(n345), .ZN(n309) );
  XOR2_X1 U356 ( .A(n309), .B(KEYINPUT10), .Z(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n560) );
  XOR2_X1 U358 ( .A(KEYINPUT80), .B(n560), .Z(n544) );
  XOR2_X1 U359 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n348) );
  XOR2_X1 U360 ( .A(G71GAT), .B(KEYINPUT13), .Z(n355) );
  XNOR2_X1 U361 ( .A(n312), .B(KEYINPUT32), .ZN(n316) );
  INV_X1 U362 ( .A(n316), .ZN(n314) );
  AND2_X1 U363 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  INV_X1 U364 ( .A(n315), .ZN(n313) );
  NAND2_X1 U365 ( .A1(n314), .A2(n313), .ZN(n318) );
  NAND2_X1 U366 ( .A1(n316), .A2(n315), .ZN(n317) );
  NAND2_X1 U367 ( .A1(n318), .A2(n317), .ZN(n321) );
  XOR2_X1 U368 ( .A(G176GAT), .B(G64GAT), .Z(n392) );
  XOR2_X1 U369 ( .A(KEYINPUT72), .B(KEYINPUT75), .Z(n319) );
  XOR2_X1 U370 ( .A(n355), .B(n322), .Z(n329) );
  XOR2_X1 U371 ( .A(G204GAT), .B(G78GAT), .Z(n429) );
  XNOR2_X1 U372 ( .A(G120GAT), .B(G148GAT), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n323), .B(G57GAT), .ZN(n397) );
  XNOR2_X1 U374 ( .A(n429), .B(n397), .ZN(n327) );
  XOR2_X1 U375 ( .A(KEYINPUT33), .B(KEYINPUT74), .Z(n325) );
  XNOR2_X1 U376 ( .A(KEYINPUT31), .B(KEYINPUT73), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  INV_X1 U378 ( .A(n331), .ZN(n372) );
  NAND2_X1 U379 ( .A1(n372), .A2(KEYINPUT41), .ZN(n333) );
  INV_X1 U380 ( .A(KEYINPUT41), .ZN(n330) );
  NAND2_X1 U381 ( .A1(n331), .A2(n330), .ZN(n332) );
  NAND2_X1 U382 ( .A1(n333), .A2(n332), .ZN(n334) );
  XOR2_X1 U383 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n336) );
  XNOR2_X1 U384 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G22GAT), .Z(n356) );
  XNOR2_X1 U387 ( .A(n337), .B(n356), .ZN(n341) );
  XOR2_X1 U388 ( .A(G113GAT), .B(G1GAT), .Z(n410) );
  XOR2_X1 U389 ( .A(KEYINPUT70), .B(n410), .Z(n339) );
  NAND2_X1 U390 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n388) );
  XOR2_X1 U394 ( .A(n342), .B(n388), .Z(n344) );
  XNOR2_X1 U395 ( .A(G141GAT), .B(G197GAT), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n346) );
  XOR2_X1 U397 ( .A(n346), .B(n345), .Z(n578) );
  NAND2_X1 U398 ( .A1(n555), .A2(n578), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n370) );
  XOR2_X1 U400 ( .A(G211GAT), .B(G155GAT), .Z(n350) );
  XNOR2_X1 U401 ( .A(G183GAT), .B(G127GAT), .ZN(n349) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U403 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n352) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U406 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U408 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U409 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n360) );
  NAND2_X1 U410 ( .A1(G231GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U412 ( .A(n362), .B(n361), .Z(n367) );
  XOR2_X1 U413 ( .A(G64GAT), .B(G57GAT), .Z(n364) );
  XNOR2_X1 U414 ( .A(G1GAT), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U416 ( .A(n365), .B(KEYINPUT82), .ZN(n366) );
  XOR2_X1 U417 ( .A(n367), .B(n366), .Z(n587) );
  INV_X1 U418 ( .A(n587), .ZN(n573) );
  INV_X1 U419 ( .A(n560), .ZN(n368) );
  AND2_X1 U420 ( .A1(n573), .A2(n368), .ZN(n369) );
  NAND2_X1 U421 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n371), .B(KEYINPUT47), .ZN(n377) );
  INV_X1 U423 ( .A(n372), .ZN(n583) );
  XNOR2_X1 U424 ( .A(KEYINPUT36), .B(n544), .ZN(n590) );
  NOR2_X1 U425 ( .A1(n573), .A2(n590), .ZN(n373) );
  XNOR2_X1 U426 ( .A(n373), .B(KEYINPUT45), .ZN(n374) );
  XNOR2_X1 U427 ( .A(n578), .B(KEYINPUT71), .ZN(n564) );
  NAND2_X1 U428 ( .A1(n374), .A2(n564), .ZN(n375) );
  NOR2_X1 U429 ( .A1(n583), .A2(n375), .ZN(n376) );
  NOR2_X1 U430 ( .A1(n377), .A2(n376), .ZN(n378) );
  XOR2_X1 U431 ( .A(KEYINPUT48), .B(n378), .Z(n531) );
  XOR2_X1 U432 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n380) );
  NAND2_X1 U433 ( .A1(G226GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U435 ( .A(n381), .B(G204GAT), .Z(n386) );
  XOR2_X1 U436 ( .A(G183GAT), .B(KEYINPUT17), .Z(n383) );
  XNOR2_X1 U437 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n437) );
  XNOR2_X1 U439 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n384), .B(G211GAT), .ZN(n428) );
  XNOR2_X1 U441 ( .A(n437), .B(n428), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U443 ( .A(n387), .B(G92GAT), .Z(n390) );
  XNOR2_X1 U444 ( .A(G36GAT), .B(n388), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U447 ( .A(n394), .B(n393), .Z(n483) );
  AND2_X1 U448 ( .A1(n531), .A2(n483), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n395), .B(KEYINPUT54), .ZN(n417) );
  XOR2_X1 U450 ( .A(n397), .B(n396), .Z(n404) );
  XOR2_X1 U451 ( .A(KEYINPUT0), .B(G127GAT), .Z(n449) );
  XOR2_X1 U452 ( .A(G155GAT), .B(KEYINPUT3), .Z(n399) );
  XNOR2_X1 U453 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n423) );
  XOR2_X1 U455 ( .A(n423), .B(KEYINPUT6), .Z(n401) );
  NAND2_X1 U456 ( .A1(G225GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n449), .B(n402), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n416) );
  XOR2_X1 U460 ( .A(KEYINPUT95), .B(KEYINPUT93), .Z(n406) );
  XNOR2_X1 U461 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n414) );
  XOR2_X1 U463 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n408) );
  XNOR2_X1 U464 ( .A(KEYINPUT92), .B(KEYINPUT1), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U466 ( .A(n409), .B(G85GAT), .Z(n412) );
  XNOR2_X1 U467 ( .A(G29GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U469 ( .A(n414), .B(n413), .Z(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n472) );
  XNOR2_X1 U471 ( .A(KEYINPUT96), .B(n472), .ZN(n518) );
  NAND2_X1 U472 ( .A1(n417), .A2(n518), .ZN(n418) );
  XNOR2_X1 U473 ( .A(n418), .B(KEYINPUT65), .ZN(n576) );
  XOR2_X1 U474 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n420) );
  XNOR2_X1 U475 ( .A(G162GAT), .B(G106GAT), .ZN(n419) );
  XNOR2_X1 U476 ( .A(n420), .B(n419), .ZN(n435) );
  XOR2_X1 U477 ( .A(G148GAT), .B(KEYINPUT23), .Z(n422) );
  XNOR2_X1 U478 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n421) );
  XNOR2_X1 U479 ( .A(n422), .B(n421), .ZN(n427) );
  XOR2_X1 U480 ( .A(n423), .B(KEYINPUT90), .Z(n425) );
  NAND2_X1 U481 ( .A1(G228GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n431) );
  XNOR2_X1 U485 ( .A(G50GAT), .B(G218GAT), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n465) );
  NAND2_X1 U489 ( .A1(n576), .A2(n465), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n436), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U491 ( .A(n437), .B(G176GAT), .Z(n439) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n455) );
  XOR2_X1 U494 ( .A(G71GAT), .B(KEYINPUT20), .Z(n441) );
  XNOR2_X1 U495 ( .A(KEYINPUT88), .B(KEYINPUT85), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U497 ( .A(G120GAT), .B(G113GAT), .Z(n443) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(G15GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n453) );
  XOR2_X1 U501 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n447) );
  XNOR2_X1 U502 ( .A(G99GAT), .B(G190GAT), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U504 ( .A(n448), .B(G134GAT), .Z(n451) );
  XNOR2_X1 U505 ( .A(G43GAT), .B(n449), .ZN(n450) );
  XNOR2_X1 U506 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n454) );
  INV_X1 U508 ( .A(n532), .ZN(n466) );
  NAND2_X1 U509 ( .A1(n456), .A2(n466), .ZN(n572) );
  NOR2_X1 U510 ( .A1(n544), .A2(n572), .ZN(n459) );
  NOR2_X1 U511 ( .A1(n583), .A2(n564), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT76), .ZN(n494) );
  XNOR2_X1 U513 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n461) );
  XOR2_X1 U514 ( .A(n461), .B(n465), .Z(n526) );
  INV_X1 U515 ( .A(n526), .ZN(n535) );
  NOR2_X1 U516 ( .A1(n466), .A2(n535), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT27), .B(n483), .Z(n468) );
  NOR2_X1 U518 ( .A1(n518), .A2(n468), .ZN(n530) );
  NAND2_X1 U519 ( .A1(n462), .A2(n530), .ZN(n475) );
  NAND2_X1 U520 ( .A1(n483), .A2(n466), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n465), .A2(n463), .ZN(n464) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT25), .ZN(n470) );
  NOR2_X1 U523 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U524 ( .A(KEYINPUT26), .B(n467), .ZN(n577) );
  INV_X1 U525 ( .A(n577), .ZN(n549) );
  NOR2_X1 U526 ( .A1(n468), .A2(n549), .ZN(n469) );
  NOR2_X1 U527 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U528 ( .A(KEYINPUT99), .B(n471), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n473), .A2(n472), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n489) );
  XOR2_X1 U531 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n477) );
  NAND2_X1 U532 ( .A1(n544), .A2(n587), .ZN(n476) );
  XNOR2_X1 U533 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n489), .A2(n478), .ZN(n479) );
  XOR2_X1 U535 ( .A(KEYINPUT100), .B(n479), .Z(n508) );
  NAND2_X1 U536 ( .A1(n494), .A2(n508), .ZN(n487) );
  NOR2_X1 U537 ( .A1(n518), .A2(n487), .ZN(n481) );
  XNOR2_X1 U538 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G1GAT), .B(n482), .ZN(G1324GAT) );
  INV_X1 U541 ( .A(n483), .ZN(n520) );
  NOR2_X1 U542 ( .A1(n520), .A2(n487), .ZN(n484) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n484), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n532), .A2(n487), .ZN(n486) );
  XNOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U547 ( .A1(n526), .A2(n487), .ZN(n488) );
  XOR2_X1 U548 ( .A(G22GAT), .B(n488), .Z(G1327GAT) );
  NAND2_X1 U549 ( .A1(n573), .A2(n489), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT102), .B(n490), .ZN(n491) );
  NOR2_X1 U551 ( .A1(n590), .A2(n491), .ZN(n493) );
  XNOR2_X1 U552 ( .A(KEYINPUT103), .B(KEYINPUT37), .ZN(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(n517) );
  NAND2_X1 U554 ( .A1(n494), .A2(n517), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(KEYINPUT38), .ZN(n496) );
  XNOR2_X1 U556 ( .A(KEYINPUT104), .B(n496), .ZN(n506) );
  NOR2_X1 U557 ( .A1(n506), .A2(n518), .ZN(n500) );
  XOR2_X1 U558 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n498) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U562 ( .A1(n520), .A2(n506), .ZN(n501) );
  XOR2_X1 U563 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n503) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n502) );
  XNOR2_X1 U566 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U567 ( .A1(n532), .A2(n506), .ZN(n504) );
  XOR2_X1 U568 ( .A(n505), .B(n504), .Z(G1330GAT) );
  NOR2_X1 U569 ( .A1(n526), .A2(n506), .ZN(n507) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  XNOR2_X1 U571 ( .A(n555), .B(KEYINPUT109), .ZN(n567) );
  NOR2_X1 U572 ( .A1(n578), .A2(n567), .ZN(n516) );
  NAND2_X1 U573 ( .A1(n516), .A2(n508), .ZN(n513) );
  NOR2_X1 U574 ( .A1(n518), .A2(n513), .ZN(n509) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n509), .Z(n510) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n510), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n520), .A2(n513), .ZN(n511) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n532), .A2(n513), .ZN(n512) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n513), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n517), .A2(n516), .ZN(n525) );
  NOR2_X1 U585 ( .A1(n518), .A2(n525), .ZN(n519) );
  XOR2_X1 U586 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U587 ( .A1(n520), .A2(n525), .ZN(n521) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(n521), .Z(n522) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U590 ( .A1(n532), .A2(n525), .ZN(n524) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U596 ( .A(G106GAT), .B(n529), .Z(G1339GAT) );
  NAND2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n548) );
  NOR2_X1 U598 ( .A1(n532), .A2(n548), .ZN(n533) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(n533), .Z(n534) );
  NOR2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U601 ( .A(KEYINPUT115), .B(n536), .ZN(n543) );
  NOR2_X1 U602 ( .A1(n564), .A2(n543), .ZN(n537) );
  XOR2_X1 U603 ( .A(G113GAT), .B(n537), .Z(G1340GAT) );
  NOR2_X1 U604 ( .A1(n567), .A2(n543), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NOR2_X1 U607 ( .A1(n573), .A2(n543), .ZN(n541) );
  XNOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U610 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U614 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT118), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n578), .A2(n561), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n553) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT53), .B(n554), .Z(n557) );
  NAND2_X1 U623 ( .A1(n561), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  XOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT121), .Z(n559) );
  NAND2_X1 U626 ( .A1(n561), .A2(n587), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NOR2_X1 U631 ( .A1(n564), .A2(n572), .ZN(n566) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XNOR2_X1 U634 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n572), .A2(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1350GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n589) );
  INV_X1 U643 ( .A(n589), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(KEYINPUT126), .Z(n580) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U647 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

