

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n407) );
  XNOR2_X1 U324 ( .A(n406), .B(n405), .ZN(n535) );
  NOR2_X1 U325 ( .A1(n536), .A2(n448), .ZN(n572) );
  XNOR2_X1 U326 ( .A(n386), .B(KEYINPUT31), .ZN(n387) );
  XNOR2_X1 U327 ( .A(n388), .B(n387), .ZN(n391) );
  XNOR2_X1 U328 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n405) );
  XNOR2_X1 U329 ( .A(n408), .B(n407), .ZN(n579) );
  INV_X1 U330 ( .A(G183GAT), .ZN(n450) );
  XNOR2_X1 U331 ( .A(n450), .B(KEYINPUT124), .ZN(n451) );
  XNOR2_X1 U332 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  XOR2_X1 U333 ( .A(G22GAT), .B(G155GAT), .Z(n421) );
  XOR2_X1 U334 ( .A(G64GAT), .B(n421), .Z(n292) );
  XOR2_X1 U335 ( .A(G15GAT), .B(G127GAT), .Z(n317) );
  XNOR2_X1 U336 ( .A(n317), .B(G78GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U338 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n294) );
  NAND2_X1 U339 ( .A1(G231GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n296), .B(n295), .Z(n298) );
  XOR2_X1 U342 ( .A(KEYINPUT72), .B(G1GAT), .Z(n360) );
  XNOR2_X1 U343 ( .A(n360), .B(KEYINPUT81), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U345 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n300) );
  XNOR2_X1 U346 ( .A(KEYINPUT14), .B(KEYINPUT82), .ZN(n299) );
  XNOR2_X1 U347 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U348 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U349 ( .A(G57GAT), .B(KEYINPUT73), .Z(n304) );
  XNOR2_X1 U350 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n304), .B(n303), .ZN(n381) );
  XNOR2_X1 U352 ( .A(G8GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n305), .B(G211GAT), .ZN(n338) );
  XNOR2_X1 U354 ( .A(n381), .B(n338), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n307), .B(n306), .ZN(n482) );
  XNOR2_X1 U356 ( .A(n482), .B(KEYINPUT112), .ZN(n545) );
  XOR2_X1 U357 ( .A(G120GAT), .B(KEYINPUT0), .Z(n309) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G134GAT), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n434) );
  XOR2_X1 U360 ( .A(G71GAT), .B(G183GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(G190GAT), .B(KEYINPUT20), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n434), .B(n312), .ZN(n322) );
  XOR2_X1 U364 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n314) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n332) );
  XOR2_X1 U367 ( .A(n332), .B(G176GAT), .Z(n316) );
  NAND2_X1 U368 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n318) );
  XOR2_X1 U370 ( .A(n318), .B(n317), .Z(n320) );
  XNOR2_X1 U371 ( .A(G43GAT), .B(G99GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n536) );
  XOR2_X1 U374 ( .A(G36GAT), .B(G190GAT), .Z(n351) );
  INV_X1 U375 ( .A(G197GAT), .ZN(n326) );
  XOR2_X1 U376 ( .A(G218GAT), .B(KEYINPUT85), .Z(n324) );
  XNOR2_X1 U377 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n425) );
  XOR2_X1 U380 ( .A(G176GAT), .B(G64GAT), .Z(n385) );
  XNOR2_X1 U381 ( .A(n425), .B(n385), .ZN(n328) );
  XOR2_X1 U382 ( .A(KEYINPUT91), .B(G92GAT), .Z(n327) );
  XNOR2_X1 U383 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U384 ( .A(n351), .B(n329), .Z(n331) );
  NAND2_X1 U385 ( .A1(G226GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n333) );
  NAND2_X1 U387 ( .A1(n332), .A2(n333), .ZN(n337) );
  INV_X1 U388 ( .A(n332), .ZN(n335) );
  INV_X1 U389 ( .A(n333), .ZN(n334) );
  NAND2_X1 U390 ( .A1(n335), .A2(n334), .ZN(n336) );
  AND2_X1 U391 ( .A1(n337), .A2(n336), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n463) );
  XOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT78), .Z(n341) );
  XNOR2_X1 U394 ( .A(G218GAT), .B(KEYINPUT77), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n347) );
  XOR2_X1 U396 ( .A(G29GAT), .B(G43GAT), .Z(n343) );
  XNOR2_X1 U397 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n361) );
  XOR2_X1 U399 ( .A(G106GAT), .B(n361), .Z(n345) );
  NAND2_X1 U400 ( .A1(G232GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n357) );
  XOR2_X1 U403 ( .A(KEYINPUT65), .B(KEYINPUT11), .Z(n349) );
  XNOR2_X1 U404 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n348) );
  XNOR2_X1 U405 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U406 ( .A(n351), .B(n350), .Z(n355) );
  XOR2_X1 U407 ( .A(G50GAT), .B(G162GAT), .Z(n422) );
  XOR2_X1 U408 ( .A(G85GAT), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U409 ( .A(G99GAT), .B(KEYINPUT76), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n389) );
  XNOR2_X1 U411 ( .A(n422), .B(n389), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U413 ( .A(n357), .B(n356), .ZN(n571) );
  XOR2_X1 U414 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n359) );
  XNOR2_X1 U415 ( .A(KEYINPUT29), .B(KEYINPUT69), .ZN(n358) );
  XNOR2_X1 U416 ( .A(n359), .B(n358), .ZN(n365) );
  XOR2_X1 U417 ( .A(n360), .B(G36GAT), .Z(n363) );
  XNOR2_X1 U418 ( .A(n361), .B(G50GAT), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n378) );
  XOR2_X1 U421 ( .A(G15GAT), .B(G197GAT), .Z(n367) );
  XNOR2_X1 U422 ( .A(G141GAT), .B(G22GAT), .ZN(n366) );
  XNOR2_X1 U423 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U424 ( .A(KEYINPUT30), .B(G8GAT), .Z(n369) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(G113GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U427 ( .A(n371), .B(n370), .Z(n376) );
  XOR2_X1 U428 ( .A(KEYINPUT68), .B(KEYINPUT67), .Z(n373) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U431 ( .A(KEYINPUT66), .B(n374), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n582) );
  XOR2_X1 U434 ( .A(G78GAT), .B(G148GAT), .Z(n380) );
  XNOR2_X1 U435 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n414) );
  XNOR2_X1 U437 ( .A(n414), .B(n381), .ZN(n393) );
  XOR2_X1 U438 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n383) );
  XNOR2_X1 U439 ( .A(G120GAT), .B(G204GAT), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U441 ( .A(n385), .B(n384), .Z(n388) );
  NAND2_X1 U442 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XOR2_X1 U443 ( .A(n389), .B(KEYINPUT74), .Z(n390) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U445 ( .A(n393), .B(n392), .ZN(n399) );
  XNOR2_X1 U446 ( .A(n399), .B(KEYINPUT41), .ZN(n566) );
  NAND2_X1 U447 ( .A1(n582), .A2(n566), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n394), .B(KEYINPUT46), .ZN(n395) );
  NAND2_X1 U449 ( .A1(n395), .A2(n545), .ZN(n396) );
  NOR2_X1 U450 ( .A1(n571), .A2(n396), .ZN(n397) );
  XNOR2_X1 U451 ( .A(KEYINPUT47), .B(n397), .ZN(n404) );
  INV_X1 U452 ( .A(n571), .ZN(n483) );
  XNOR2_X1 U453 ( .A(KEYINPUT36), .B(n483), .ZN(n591) );
  NOR2_X1 U454 ( .A1(n591), .A2(n482), .ZN(n398) );
  XNOR2_X1 U455 ( .A(KEYINPUT45), .B(n398), .ZN(n400) );
  NAND2_X1 U456 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n401), .B(KEYINPUT113), .ZN(n402) );
  INV_X1 U458 ( .A(n582), .ZN(n504) );
  NAND2_X1 U459 ( .A1(n402), .A2(n504), .ZN(n403) );
  NAND2_X1 U460 ( .A1(n404), .A2(n403), .ZN(n406) );
  NAND2_X1 U461 ( .A1(n463), .A2(n535), .ZN(n408) );
  XOR2_X1 U462 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n410) );
  NAND2_X1 U463 ( .A1(G228GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U465 ( .A(n411), .B(G211GAT), .Z(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n413) );
  XNOR2_X1 U467 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n433) );
  XNOR2_X1 U469 ( .A(n433), .B(n414), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U471 ( .A(KEYINPUT84), .B(KEYINPUT87), .Z(n418) );
  XNOR2_X1 U472 ( .A(KEYINPUT88), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U474 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U477 ( .A(n426), .B(n425), .Z(n465) );
  XOR2_X1 U478 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n428) );
  XNOR2_X1 U479 ( .A(G1GAT), .B(G57GAT), .ZN(n427) );
  XNOR2_X1 U480 ( .A(n428), .B(n427), .ZN(n444) );
  XOR2_X1 U481 ( .A(G155GAT), .B(G162GAT), .Z(n430) );
  XNOR2_X1 U482 ( .A(G127GAT), .B(G148GAT), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U484 ( .A(G29GAT), .B(G85GAT), .Z(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n440) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U487 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n436) );
  XNOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U491 ( .A(n440), .B(n439), .ZN(n442) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n578) );
  INV_X1 U495 ( .A(n578), .ZN(n445) );
  NOR2_X1 U496 ( .A1(n465), .A2(n445), .ZN(n446) );
  AND2_X1 U497 ( .A1(n579), .A2(n446), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  INV_X1 U499 ( .A(n572), .ZN(n449) );
  NOR2_X1 U500 ( .A1(n545), .A2(n449), .ZN(n452) );
  XNOR2_X1 U501 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n479) );
  XNOR2_X1 U502 ( .A(n465), .B(KEYINPUT28), .ZN(n539) );
  XOR2_X1 U503 ( .A(KEYINPUT27), .B(n463), .Z(n461) );
  NOR2_X1 U504 ( .A1(n461), .A2(n578), .ZN(n453) );
  NAND2_X1 U505 ( .A1(n453), .A2(KEYINPUT92), .ZN(n457) );
  INV_X1 U506 ( .A(n453), .ZN(n455) );
  INV_X1 U507 ( .A(KEYINPUT92), .ZN(n454) );
  NAND2_X1 U508 ( .A1(n455), .A2(n454), .ZN(n456) );
  NAND2_X1 U509 ( .A1(n457), .A2(n456), .ZN(n534) );
  NAND2_X1 U510 ( .A1(n534), .A2(n536), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n539), .A2(n458), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT93), .ZN(n471) );
  NAND2_X1 U513 ( .A1(n465), .A2(n536), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n460), .B(KEYINPUT26), .ZN(n581) );
  NOR2_X1 U515 ( .A1(n581), .A2(n461), .ZN(n462) );
  XOR2_X1 U516 ( .A(KEYINPUT94), .B(n462), .Z(n468) );
  INV_X1 U517 ( .A(n463), .ZN(n525) );
  NOR2_X1 U518 ( .A1(n536), .A2(n525), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT25), .B(n466), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U522 ( .A1(n469), .A2(n578), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n471), .A2(n470), .ZN(n486) );
  INV_X1 U524 ( .A(n591), .ZN(n472) );
  AND2_X1 U525 ( .A1(n472), .A2(n482), .ZN(n473) );
  NAND2_X1 U526 ( .A1(n486), .A2(n473), .ZN(n475) );
  XOR2_X1 U527 ( .A(KEYINPUT37), .B(KEYINPUT98), .Z(n474) );
  XNOR2_X1 U528 ( .A(n475), .B(n474), .ZN(n521) );
  NAND2_X1 U529 ( .A1(n582), .A2(n399), .ZN(n488) );
  NOR2_X1 U530 ( .A1(n521), .A2(n488), .ZN(n476) );
  XNOR2_X1 U531 ( .A(n476), .B(KEYINPUT38), .ZN(n477) );
  XNOR2_X1 U532 ( .A(n477), .B(KEYINPUT99), .ZN(n502) );
  NOR2_X1 U533 ( .A1(n536), .A2(n502), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n481) );
  INV_X1 U535 ( .A(G43GAT), .ZN(n480) );
  XNOR2_X1 U536 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  INV_X1 U537 ( .A(n482), .ZN(n587) );
  NAND2_X1 U538 ( .A1(n587), .A2(n483), .ZN(n484) );
  XNOR2_X1 U539 ( .A(n484), .B(KEYINPUT83), .ZN(n485) );
  XNOR2_X1 U540 ( .A(n485), .B(KEYINPUT16), .ZN(n487) );
  NAND2_X1 U541 ( .A1(n487), .A2(n486), .ZN(n506) );
  OR2_X1 U542 ( .A1(n488), .A2(n506), .ZN(n497) );
  NOR2_X1 U543 ( .A1(n578), .A2(n497), .ZN(n489) );
  XOR2_X1 U544 ( .A(n489), .B(KEYINPUT34), .Z(n490) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n490), .ZN(G1324GAT) );
  NOR2_X1 U546 ( .A1(n525), .A2(n497), .ZN(n492) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(KEYINPUT95), .ZN(n491) );
  XNOR2_X1 U548 ( .A(n492), .B(n491), .ZN(G1325GAT) );
  NOR2_X1 U549 ( .A1(n497), .A2(n536), .ZN(n496) );
  XOR2_X1 U550 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n494) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  INV_X1 U554 ( .A(n539), .ZN(n530) );
  NOR2_X1 U555 ( .A1(n530), .A2(n497), .ZN(n498) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n498), .Z(G1327GAT) );
  NOR2_X1 U557 ( .A1(n502), .A2(n578), .ZN(n500) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U560 ( .A1(n502), .A2(n525), .ZN(n501) );
  XOR2_X1 U561 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  NOR2_X1 U562 ( .A1(n530), .A2(n502), .ZN(n503) );
  XOR2_X1 U563 ( .A(G50GAT), .B(n503), .Z(G1331GAT) );
  NAND2_X1 U564 ( .A1(n566), .A2(n504), .ZN(n505) );
  XOR2_X1 U565 ( .A(KEYINPUT101), .B(n505), .Z(n520) );
  NOR2_X1 U566 ( .A1(n520), .A2(n506), .ZN(n507) );
  XOR2_X1 U567 ( .A(KEYINPUT102), .B(n507), .Z(n516) );
  NOR2_X1 U568 ( .A1(n516), .A2(n578), .ZN(n509) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n510), .ZN(G1332GAT) );
  XNOR2_X1 U572 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n512) );
  NOR2_X1 U573 ( .A1(n525), .A2(n516), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U576 ( .A1(n536), .A2(n516), .ZN(n514) );
  XOR2_X1 U577 ( .A(KEYINPUT106), .B(n514), .Z(n515) );
  XNOR2_X1 U578 ( .A(G71GAT), .B(n515), .ZN(G1334GAT) );
  XNOR2_X1 U579 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n518) );
  NOR2_X1 U580 ( .A1(n530), .A2(n516), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n519), .Z(G1335GAT) );
  OR2_X1 U583 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X1 U584 ( .A1(n578), .A2(n529), .ZN(n523) );
  XNOR2_X1 U585 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n529), .ZN(n526) );
  XOR2_X1 U589 ( .A(KEYINPUT110), .B(n526), .Z(n527) );
  XNOR2_X1 U590 ( .A(G92GAT), .B(n527), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n536), .A2(n529), .ZN(n528) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n528), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U594 ( .A(KEYINPUT44), .B(KEYINPUT111), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n552) );
  NOR2_X1 U598 ( .A1(n536), .A2(n552), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT114), .B(n537), .Z(n538) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n582), .A2(n549), .ZN(n540) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U604 ( .A1(n549), .A2(n566), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n543), .Z(G1341GAT) );
  INV_X1 U607 ( .A(n549), .ZN(n544) );
  NOR2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U609 ( .A(KEYINPUT50), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n571), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n581), .A2(n552), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n582), .A2(n562), .ZN(n553) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT119), .B(KEYINPUT53), .Z(n555) );
  XNOR2_X1 U619 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(n559) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n562), .A2(n566), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n587), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(KEYINPUT120), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n561), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n571), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n582), .A2(n572), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n568) );
  NAND2_X1 U634 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U636 ( .A(G176GAT), .B(KEYINPUT56), .Z(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(n575), .ZN(G1351GAT) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(KEYINPUT60), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT126), .B(n577), .Z(n584) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n588), .A2(n582), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n586) );
  INV_X1 U650 ( .A(n588), .ZN(n590) );
  OR2_X1 U651 ( .A1(n590), .A2(n399), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G211GAT), .B(n589), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

