//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1254, new_n1255, new_n1256, new_n1257,
    new_n1258, new_n1259;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT0), .Z(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n222), .B1(new_n203), .B2(new_n223), .C1(new_n206), .C2(new_n224), .ZN(new_n225));
  AOI211_X1 g0025(.A(new_n221), .B(new_n225), .C1(G58), .C2(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n212), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n211), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n217), .B(new_n228), .C1(new_n230), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n220), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  INV_X1    g0044(.A(G87), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n206), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n247), .B(new_n251), .ZN(G351));
  OR2_X1    g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G222), .ZN(new_n258));
  OAI21_X1  g0058(.A(KEYINPUT67), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n256), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT68), .B(G223), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n262), .A2(G77), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT67), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n255), .A2(new_n267), .A3(G222), .A4(new_n256), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n259), .A2(new_n265), .A3(new_n266), .A4(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n210), .B(G274), .C1(G41), .C2(G45), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT66), .B(G1), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(new_n270), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n271), .A2(new_n272), .A3(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G169), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n229), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT69), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n273), .A2(G20), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G50), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n204), .A2(G20), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  INV_X1    g0088(.A(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n211), .A2(new_n289), .A3(KEYINPUT71), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT71), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G20), .B2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT8), .ZN(new_n295));
  OAI21_X1  g0095(.A(KEYINPUT70), .B1(new_n295), .B2(G58), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(KEYINPUT8), .B2(new_n202), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(KEYINPUT70), .A3(G58), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n211), .A2(G33), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n287), .B1(new_n288), .B2(new_n294), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n283), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n286), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n273), .A2(G13), .A3(G20), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(new_n201), .ZN(new_n306));
  AND2_X1   g0106(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n279), .A2(new_n307), .A3(KEYINPUT72), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n278), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT72), .B1(new_n279), .B2(new_n307), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT73), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT85), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n260), .A2(new_n261), .A3(G20), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT83), .B(KEYINPUT7), .Z(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT7), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(G68), .C1(new_n318), .C2(new_n315), .ZN(new_n319));
  XNOR2_X1  g0119(.A(G58), .B(G68), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n293), .A2(G159), .B1(new_n320), .B2(G20), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n319), .A2(KEYINPUT16), .A3(new_n321), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n253), .A2(new_n318), .A3(new_n211), .A4(new_n254), .ZN(new_n323));
  OAI211_X1 g0123(.A(G68), .B(new_n323), .C1(new_n315), .C2(new_n316), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n321), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT16), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n327), .A3(new_n281), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT84), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n299), .B1(G20), .B2(new_n273), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n283), .B1(new_n305), .B2(new_n299), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n280), .A2(new_n229), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n325), .B2(new_n326), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT84), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n322), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n255), .A2(G223), .A3(new_n256), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n255), .A2(G226), .A3(G1698), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n337), .B(new_n338), .C1(new_n289), .C2(new_n245), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n270), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n276), .A2(G232), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n272), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G169), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n309), .B2(new_n342), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n336), .A2(KEYINPUT18), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT18), .B1(new_n336), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n314), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n333), .A2(new_n334), .A3(new_n322), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n334), .B1(new_n333), .B2(new_n322), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n330), .A2(new_n283), .ZN(new_n351));
  INV_X1    g0151(.A(new_n299), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n304), .B2(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n349), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n342), .A2(new_n309), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(G169), .B2(new_n342), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n348), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n336), .A2(KEYINPUT18), .A3(new_n344), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(KEYINPUT85), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT17), .ZN(new_n360));
  INV_X1    g0160(.A(new_n342), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(G190), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n354), .A2(new_n360), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(new_n329), .A3(new_n331), .A4(new_n335), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT17), .B1(new_n367), .B2(new_n363), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n347), .A2(new_n359), .A3(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n313), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n307), .A2(KEYINPUT9), .B1(G190), .B2(new_n278), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n278), .A2(new_n362), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT76), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n303), .A2(new_n306), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT9), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT76), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n378), .B1(new_n278), .B2(new_n362), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n372), .A2(new_n374), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  XNOR2_X1  g0180(.A(new_n380), .B(KEYINPUT10), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G20), .A2(G77), .ZN(new_n382));
  XOR2_X1   g0182(.A(KEYINPUT15), .B(G87), .Z(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(KEYINPUT8), .B(G58), .ZN(new_n385));
  XNOR2_X1  g0185(.A(new_n385), .B(KEYINPUT75), .ZN(new_n386));
  OAI221_X1 g0186(.A(new_n382), .B1(new_n300), .B2(new_n384), .C1(new_n386), .C2(new_n294), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n281), .B1(new_n250), .B2(new_n305), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n284), .A2(new_n332), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n250), .B2(new_n389), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n263), .A2(G238), .B1(G107), .B2(new_n262), .ZN(new_n391));
  INV_X1    g0191(.A(G232), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(new_n257), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n270), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n276), .A2(G244), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n272), .A3(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G190), .ZN(new_n397));
  OR3_X1    g0197(.A1(new_n396), .A2(KEYINPUT74), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT74), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n390), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n396), .A2(G200), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n396), .A2(G179), .ZN(new_n403));
  INV_X1    g0203(.A(G169), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n396), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n390), .A3(new_n405), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n381), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n289), .A2(new_n206), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n253), .A2(new_n254), .B1(new_n392), .B2(G1698), .ZN(new_n409));
  OR2_X1    g0209(.A1(G226), .A2(G1698), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n411), .A2(new_n275), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT13), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n274), .A2(G238), .A3(new_n275), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .A4(new_n272), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n272), .C1(new_n411), .C2(new_n275), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT78), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(KEYINPUT78), .A3(KEYINPUT13), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G190), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n211), .A2(G33), .A3(G77), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n293), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n283), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n425), .A2(KEYINPUT11), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n305), .A2(new_n203), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n425), .A2(KEYINPUT11), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n284), .A2(G68), .A3(new_n332), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n430), .B(KEYINPUT79), .Z(new_n431));
  NAND4_X1  g0231(.A1(new_n426), .A2(new_n428), .A3(new_n429), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n415), .A2(new_n417), .A3(KEYINPUT77), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n416), .A2(KEYINPUT77), .A3(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n422), .A2(new_n433), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(KEYINPUT80), .A2(G169), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n434), .A2(new_n435), .A3(new_n442), .A4(new_n439), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT81), .B1(new_n421), .B2(G179), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT81), .ZN(new_n445));
  AOI211_X1 g0245(.A(new_n445), .B(new_n309), .C1(new_n419), .C2(new_n420), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n441), .B(new_n443), .C1(new_n444), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n438), .B1(new_n447), .B2(new_n432), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n448), .A2(KEYINPUT82), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n371), .A2(new_n407), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n273), .A2(G33), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n304), .A2(new_n453), .A3(G116), .A4(new_n332), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n455), .B(new_n211), .C1(G33), .C2(new_n206), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(new_n281), .C1(new_n211), .C2(G116), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT20), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  OAI221_X1 g0260(.A(new_n454), .B1(G116), .B2(new_n304), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G264), .A2(G1698), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(new_n224), .B2(G1698), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n255), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G303), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n255), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT95), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n255), .A2(new_n463), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT95), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n468), .B(new_n469), .C1(new_n465), .C2(new_n255), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n270), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G41), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT66), .A2(G1), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT66), .A2(G1), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(G45), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n472), .A2(G41), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n275), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G270), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n273), .A2(KEYINPUT89), .A3(G45), .A4(new_n473), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n270), .A2(new_n477), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(G274), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n471), .A2(new_n480), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n461), .B1(new_n486), .B2(G200), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n487), .B1(new_n397), .B2(new_n486), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n461), .A3(G169), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT21), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n480), .A2(new_n485), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n461), .A2(new_n492), .A3(G179), .A4(new_n471), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n486), .A2(new_n461), .A3(KEYINPUT21), .A4(G169), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT23), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(new_n207), .A3(G20), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n496), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT96), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n496), .A2(new_n498), .A3(new_n499), .A4(KEYINPUT96), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(G20), .B1(new_n253), .B2(new_n254), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT22), .A3(G87), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n211), .B(G87), .C1(new_n260), .C2(new_n261), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT22), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT24), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n502), .A2(new_n503), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n513), .A3(new_n509), .A4(new_n506), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n332), .A2(KEYINPUT69), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n281), .A2(new_n282), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n304), .B(new_n453), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n515), .A2(new_n281), .B1(G107), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n304), .A2(G107), .ZN(new_n521));
  XNOR2_X1  g0321(.A(new_n521), .B(KEYINPUT25), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n263), .A2(G257), .ZN(new_n523));
  INV_X1    g0323(.A(G250), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(new_n257), .ZN(new_n525));
  INV_X1    g0325(.A(G294), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n289), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n270), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n479), .A2(G264), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n485), .A3(new_n529), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n520), .A2(new_n522), .B1(new_n404), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g0331(.A1(new_n530), .A2(G179), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n495), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n528), .A2(new_n529), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n535), .A2(G190), .A3(new_n485), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n530), .A2(G200), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n520), .A3(new_n522), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n255), .A2(G244), .A3(G1698), .ZN(new_n539));
  OAI221_X1 g0339(.A(new_n539), .B1(new_n289), .B2(new_n219), .C1(new_n257), .C2(new_n223), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n270), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT90), .ZN(new_n542));
  INV_X1    g0342(.A(new_n273), .ZN(new_n543));
  INV_X1    g0343(.A(G45), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n542), .B(G250), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n542), .A2(new_n524), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n273), .B(G45), .C1(G274), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n541), .B1(new_n270), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n404), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n541), .B(new_n309), .C1(new_n270), .C2(new_n548), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT93), .B1(new_n518), .B2(new_n384), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n304), .A2(new_n453), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT93), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n283), .A4(new_n383), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n211), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n245), .A2(new_n206), .A3(new_n207), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT91), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n255), .A2(new_n211), .A3(G68), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n211), .A2(G33), .A3(G97), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT19), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n559), .A2(KEYINPUT91), .A3(new_n560), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n563), .A2(new_n564), .A3(new_n567), .A4(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n281), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n304), .A2(new_n383), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT92), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT92), .ZN(new_n574));
  AOI211_X1 g0374(.A(new_n574), .B(new_n571), .C1(new_n569), .C2(new_n281), .ZN(new_n575));
  OAI211_X1 g0375(.A(KEYINPUT94), .B(new_n557), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n559), .A2(KEYINPUT91), .A3(new_n560), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT91), .B1(new_n559), .B2(new_n560), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n505), .A2(G68), .B1(new_n566), .B2(new_n565), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n332), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n574), .B1(new_n582), .B2(new_n571), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n570), .A2(KEYINPUT92), .A3(new_n572), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT94), .B1(new_n585), .B2(new_n557), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n552), .B1(new_n577), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n540), .A2(new_n270), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n270), .B1(new_n545), .B2(new_n547), .ZN(new_n589));
  OAI21_X1  g0389(.A(G200), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n541), .B(G190), .C1(new_n270), .C2(new_n548), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n573), .A2(new_n575), .B1(new_n245), .B2(new_n518), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT87), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n206), .A2(KEYINPUT6), .ZN(new_n598));
  NAND2_X1  g0398(.A1(G97), .A2(G107), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n208), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n208), .A2(new_n599), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n597), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G20), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT86), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n293), .A2(new_n604), .A3(G77), .ZN(new_n605));
  OAI211_X1 g0405(.A(G107), .B(new_n323), .C1(new_n315), .C2(new_n316), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT86), .B1(new_n294), .B2(new_n250), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n603), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n281), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n519), .A2(G97), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n304), .A2(G97), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(KEYINPUT88), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n485), .B1(new_n224), .B2(new_n478), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT4), .ZN(new_n615));
  OAI211_X1 g0415(.A(G244), .B(new_n256), .C1(new_n260), .C2(new_n261), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n524), .B2(new_n256), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n615), .A2(new_n616), .B1(new_n618), .B2(new_n255), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n275), .B1(new_n619), .B2(new_n455), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n309), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n404), .B1(new_n614), .B2(new_n620), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n613), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n620), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n479), .A2(G257), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n625), .A2(G190), .A3(new_n485), .A4(new_n626), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n608), .A2(new_n281), .B1(G97), .B2(new_n519), .ZN(new_n628));
  OAI21_X1  g0428(.A(G200), .B1(new_n614), .B2(new_n620), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n627), .A2(new_n628), .A3(new_n612), .A4(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  AND4_X1   g0431(.A1(new_n538), .A2(new_n587), .A3(new_n595), .A4(new_n631), .ZN(new_n632));
  AND4_X1   g0432(.A1(new_n452), .A2(new_n488), .A3(new_n533), .A4(new_n632), .ZN(G372));
  NAND2_X1  g0433(.A1(new_n550), .A2(new_n551), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n557), .B1(new_n573), .B2(new_n575), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT94), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n637), .B2(new_n576), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NOR4_X1   g0439(.A1(new_n638), .A2(new_n594), .A3(new_n639), .A4(new_n624), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n638), .A2(new_n594), .A3(new_n624), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT97), .B1(new_n641), .B2(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n624), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n587), .A2(new_n595), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT97), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n639), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n640), .B1(new_n642), .B2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n587), .A2(new_n631), .A3(new_n538), .A4(new_n595), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n587), .B1(new_n649), .B2(new_n533), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n452), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n357), .A2(new_n358), .ZN(new_n654));
  INV_X1    g0454(.A(new_n406), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n447), .A2(new_n432), .B1(new_n437), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n369), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n381), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT98), .ZN(new_n660));
  INV_X1    g0460(.A(new_n313), .ZN(new_n661));
  AND3_X1   g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n653), .B1(new_n662), .B2(new_n663), .ZN(G369));
  NOR2_X1   g0464(.A1(new_n213), .A2(G20), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n273), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(G343), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n461), .A2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n495), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n495), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n488), .A2(new_n672), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT99), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n520), .A2(new_n522), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n671), .ZN(new_n679));
  AOI22_X1  g0479(.A1(new_n679), .A2(new_n538), .B1(new_n531), .B2(new_n532), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n530), .A2(new_n404), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(new_n681), .A3(new_n532), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n671), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n677), .A2(G330), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n671), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n495), .A2(new_n687), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n680), .A2(new_n688), .B1(new_n682), .B2(new_n671), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n686), .A2(new_n689), .ZN(G399));
  NOR2_X1   g0490(.A1(new_n214), .A2(G41), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n560), .A2(G116), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G1), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n231), .B2(new_n692), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT28), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n652), .A2(new_n697), .A3(new_n687), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT101), .B1(new_n649), .B2(new_n533), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n624), .A2(new_n630), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n638), .A2(new_n594), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT101), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n674), .A2(new_n682), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n701), .A2(new_n702), .A3(new_n703), .A4(new_n538), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n637), .A2(new_n576), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n594), .B1(new_n706), .B2(new_n552), .ZN(new_n707));
  AOI21_X1  g0507(.A(KEYINPUT26), .B1(new_n707), .B2(new_n643), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n587), .B1(new_n708), .B2(new_n640), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n687), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n698), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n632), .A2(new_n488), .A3(new_n533), .A4(new_n687), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n486), .A2(new_n309), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT100), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n534), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n492), .A2(G179), .A3(new_n471), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n549), .B1(new_n717), .B2(KEYINPUT100), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(new_n718), .A3(new_n621), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n716), .A2(new_n718), .A3(KEYINPUT30), .A4(new_n621), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n621), .B1(new_n535), .B2(new_n485), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n723), .A2(new_n309), .A3(new_n486), .A4(new_n549), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n671), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n726), .A2(KEYINPUT31), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(new_n728), .A3(G330), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n712), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n696), .B1(new_n731), .B2(G1), .ZN(G364));
  NAND2_X1  g0532(.A1(new_n665), .A2(G45), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n692), .A2(G1), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n735), .B1(new_n677), .B2(G330), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n677), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n229), .B1(G20), .B2(new_n404), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT103), .Z(new_n743));
  NAND2_X1  g0543(.A1(new_n215), .A2(new_n262), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n251), .A2(new_n544), .ZN(new_n745));
  AOI211_X1 g0545(.A(new_n744), .B(new_n745), .C1(new_n544), .C2(new_n232), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n215), .A2(G355), .A3(new_n255), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G116), .B2(new_n215), .ZN(new_n748));
  XOR2_X1   g0548(.A(new_n748), .B(KEYINPUT102), .Z(new_n749));
  OAI21_X1  g0549(.A(new_n743), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n211), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n752), .A2(G179), .A3(new_n362), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT106), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n309), .A2(new_n362), .A3(KEYINPUT105), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT105), .B1(new_n309), .B2(new_n362), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n752), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n757), .A2(G283), .B1(new_n761), .B2(G329), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n211), .A2(new_n309), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(G190), .A3(G200), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G326), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n397), .A3(G200), .ZN(new_n767));
  XOR2_X1   g0567(.A(KEYINPUT33), .B(G317), .Z(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(new_n397), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(G179), .A3(new_n362), .ZN(new_n771));
  INV_X1    g0571(.A(G322), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n770), .A2(new_n309), .A3(G200), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n262), .B1(new_n771), .B2(new_n772), .C1(new_n465), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n751), .A2(G179), .A3(new_n362), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n769), .B(new_n774), .C1(G311), .C2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n760), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n211), .B1(new_n778), .B2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G294), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n762), .A2(new_n766), .A3(new_n777), .A4(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n756), .A2(new_n207), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n776), .A2(KEYINPUT104), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n776), .A2(KEYINPUT104), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n783), .B1(G77), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n788), .B(new_n255), .C1(new_n245), .C2(new_n773), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n767), .A2(new_n203), .B1(new_n764), .B2(new_n201), .ZN(new_n790));
  INV_X1    g0590(.A(new_n771), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G58), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g0592(.A1(new_n761), .A2(KEYINPUT32), .A3(G159), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT32), .B1(new_n761), .B2(G159), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n206), .B2(new_n779), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n782), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n734), .B1(new_n796), .B2(new_n741), .ZN(new_n797));
  INV_X1    g0597(.A(new_n740), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n750), .B(new_n797), .C1(new_n677), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n737), .A2(new_n799), .ZN(G396));
  NAND2_X1  g0600(.A1(new_n652), .A2(new_n687), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n406), .A2(new_n671), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n400), .A2(new_n401), .B1(new_n390), .B2(new_n671), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n804), .B2(new_n655), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n801), .B(new_n806), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n807), .A2(new_n730), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n730), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n808), .A2(new_n734), .A3(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n761), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n756), .A2(new_n245), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(G116), .C2(new_n787), .ZN(new_n815));
  INV_X1    g0615(.A(G283), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n767), .A2(new_n816), .B1(new_n764), .B2(new_n465), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n262), .B1(new_n771), .B2(new_n526), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n817), .B(new_n818), .C1(new_n780), .C2(G97), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n815), .B(new_n819), .C1(new_n207), .C2(new_n773), .ZN(new_n820));
  INV_X1    g0620(.A(new_n767), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n821), .A2(G150), .B1(new_n765), .B2(G137), .ZN(new_n822));
  INV_X1    g0622(.A(G143), .ZN(new_n823));
  INV_X1    g0623(.A(G159), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n822), .B1(new_n823), .B2(new_n771), .C1(new_n786), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT34), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n255), .B1(new_n779), .B2(new_n202), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n756), .A2(new_n203), .B1(new_n201), .B2(new_n773), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT107), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n826), .B(new_n830), .C1(new_n829), .C2(new_n828), .ZN(new_n831));
  INV_X1    g0631(.A(G132), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n811), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n820), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n741), .A2(new_n738), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n834), .A2(new_n741), .B1(new_n250), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n735), .B(new_n836), .C1(new_n806), .C2(new_n739), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n810), .A2(new_n837), .ZN(G384));
  INV_X1    g0638(.A(new_n669), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n319), .A2(new_n321), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n326), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n841), .A2(new_n302), .A3(new_n322), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n331), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n370), .A2(new_n839), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n843), .B1(new_n344), .B2(new_n839), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n363), .B2(new_n367), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(KEYINPUT110), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n354), .A2(new_n364), .A3(new_n365), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n336), .A2(new_n344), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n336), .A2(new_n839), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT110), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n846), .A2(new_n854), .A3(KEYINPUT37), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n848), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  AND3_X1   g0656(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT38), .B1(new_n844), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n432), .A2(new_n671), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n448), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n432), .B(new_n671), .C1(new_n447), .C2(new_n438), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n805), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n727), .A3(new_n728), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n859), .A2(KEYINPUT40), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n863), .A2(new_n727), .A3(new_n728), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n844), .A2(KEYINPUT38), .A3(new_n856), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(new_n850), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n852), .B1(new_n369), .B2(new_n654), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n866), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(G330), .B1(new_n865), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n451), .A2(new_n729), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n879), .B(KEYINPUT111), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n727), .A2(new_n728), .ZN(new_n881));
  INV_X1    g0681(.A(new_n874), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT40), .B1(new_n882), .B2(new_n864), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n844), .A2(new_n856), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(new_n869), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n868), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n886), .A2(new_n867), .A3(new_n866), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n881), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n880), .B1(new_n452), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(KEYINPUT39), .B1(new_n857), .B2(new_n858), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n868), .A2(new_n873), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n447), .A2(new_n432), .A3(new_n687), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n357), .A2(new_n358), .A3(new_n669), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n861), .A2(new_n862), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n687), .B(new_n806), .C1(new_n647), .C2(new_n650), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n898), .B1(new_n899), .B2(new_n803), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n886), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n451), .B1(new_n698), .B2(new_n711), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n662), .A2(new_n663), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n902), .B(new_n905), .Z(new_n906));
  XNOR2_X1  g0706(.A(new_n889), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n273), .B2(new_n665), .ZN(new_n908));
  OAI21_X1  g0708(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n909));
  OAI22_X1  g0709(.A1(new_n909), .A2(new_n231), .B1(G50), .B2(new_n203), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n910), .A2(new_n213), .A3(new_n543), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT109), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n219), .B1(new_n602), .B2(KEYINPUT35), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n230), .C1(KEYINPUT35), .C2(new_n602), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT108), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT36), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n908), .A2(new_n912), .A3(new_n916), .ZN(G367));
  OAI22_X1  g0717(.A1(new_n786), .A2(new_n816), .B1(new_n812), .B2(new_n764), .ZN(new_n918));
  INV_X1    g0718(.A(new_n773), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(KEYINPUT46), .A3(G116), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT46), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n773), .B2(new_n219), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n920), .B(new_n922), .C1(new_n526), .C2(new_n767), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n207), .B2(new_n779), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT115), .ZN(new_n926));
  INV_X1    g0726(.A(G317), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n262), .B1(new_n927), .B2(new_n811), .C1(new_n756), .C2(new_n206), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n925), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  OAI221_X1 g0729(.A(new_n929), .B1(new_n926), .B2(new_n928), .C1(new_n465), .C2(new_n771), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n786), .A2(new_n201), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n756), .A2(new_n250), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n931), .B(new_n932), .C1(G137), .C2(new_n761), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n767), .A2(new_n824), .B1(new_n764), .B2(new_n823), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n255), .B1(new_n773), .B2(new_n202), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n934), .B(new_n935), .C1(new_n780), .C2(G68), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n933), .B(new_n936), .C1(new_n288), .C2(new_n771), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT47), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n741), .ZN(new_n940));
  OAI221_X1 g0740(.A(new_n742), .B1(new_n215), .B2(new_n384), .C1(new_n241), .C2(new_n744), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n735), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT116), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n593), .A2(new_n671), .ZN(new_n944));
  MUX2_X1   g0744(.A(new_n707), .B(new_n638), .S(new_n944), .Z(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n798), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n613), .A2(new_n671), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n631), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n643), .A2(new_n671), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n685), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n688), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n684), .A2(new_n955), .ZN(new_n956));
  OR3_X1    g0756(.A1(new_n956), .A2(KEYINPUT42), .A3(new_n951), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n624), .B1(new_n948), .B2(new_n682), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n687), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT42), .B1(new_n956), .B2(new_n951), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n953), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n953), .B1(new_n961), .B2(new_n954), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n962), .A2(new_n963), .B1(KEYINPUT43), .B2(new_n945), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n733), .A2(G1), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT114), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n689), .A2(new_n951), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT44), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n689), .A2(new_n951), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n686), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(new_n685), .A3(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n684), .ZN(new_n980));
  AOI21_X1  g0780(.A(KEYINPUT112), .B1(new_n980), .B2(new_n688), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(new_n956), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n677), .A2(G330), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT113), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n982), .B(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n731), .B1(new_n979), .B2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n691), .B(KEYINPUT41), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n971), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n946), .B1(new_n968), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(KEYINPUT117), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n990), .A2(KEYINPUT117), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n693), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n386), .A2(G50), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n998), .A2(KEYINPUT50), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n996), .B(new_n999), .C1(G68), .C2(G77), .ZN(new_n1000));
  AOI21_X1  g0800(.A(G45), .B1(new_n998), .B2(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n744), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n238), .A2(G45), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1002), .A2(new_n1003), .B1(new_n207), .B2(new_n214), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n996), .A2(new_n215), .A3(new_n255), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n743), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n684), .B2(new_n798), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n761), .A2(G326), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n786), .A2(new_n465), .B1(new_n927), .B2(new_n771), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT118), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n1010), .A2(new_n1011), .B1(new_n812), .B2(new_n767), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n772), .B2(new_n764), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n816), .B2(new_n779), .C1(new_n526), .C2(new_n773), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT49), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n255), .B(new_n1009), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n1017), .B2(new_n1016), .C1(new_n219), .C2(new_n756), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n756), .A2(new_n206), .B1(new_n288), .B2(new_n811), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n352), .B2(new_n821), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n764), .A2(new_n824), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n255), .B1(new_n775), .B2(new_n203), .C1(new_n250), .C2(new_n773), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(new_n780), .C2(new_n383), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(new_n201), .C2(new_n771), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1019), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1008), .B1(new_n1026), .B2(new_n741), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n986), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1027), .A2(new_n735), .B1(new_n1028), .B2(new_n971), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n731), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n986), .B1(new_n730), .B2(new_n712), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n691), .B(KEYINPUT119), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1031), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1029), .A2(new_n1034), .ZN(G393));
  AND2_X1   g0835(.A1(new_n1030), .A2(new_n979), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1033), .B1(new_n1030), .B2(new_n979), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n977), .A2(new_n978), .A3(new_n971), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n262), .B1(new_n773), .B2(new_n816), .C1(new_n465), .C2(new_n767), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1040), .B(new_n783), .C1(G322), .C2(new_n761), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n780), .A2(G116), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n776), .A2(G294), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n771), .A2(new_n812), .B1(new_n764), .B2(new_n927), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n771), .A2(new_n824), .B1(new_n764), .B2(new_n288), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT51), .Z(new_n1048));
  OAI221_X1 g0848(.A(new_n255), .B1(new_n203), .B2(new_n773), .C1(new_n811), .C2(new_n823), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n779), .A2(new_n250), .ZN(new_n1050));
  OR4_X1    g0850(.A1(new_n814), .A2(new_n1048), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n786), .A2(new_n386), .B1(new_n201), .B2(new_n767), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT120), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n1046), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n734), .B1(new_n1054), .B2(new_n741), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n742), .B1(new_n206), .B2(new_n215), .C1(new_n247), .C2(new_n744), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1055), .B(new_n1056), .C1(new_n798), .C2(new_n950), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1039), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1038), .A2(new_n1058), .ZN(G390));
  AOI22_X1  g0859(.A1(new_n757), .A2(G68), .B1(new_n761), .B2(G294), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n787), .A2(G97), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n767), .A2(new_n207), .B1(new_n764), .B2(new_n816), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1050), .A2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n262), .B1(new_n771), .B2(new_n219), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G87), .B2(new_n919), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(KEYINPUT54), .B(G143), .ZN(new_n1067));
  INV_X1    g0867(.A(G125), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n786), .A2(new_n1067), .B1(new_n811), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G50), .B2(new_n757), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n773), .A2(new_n288), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT53), .ZN(new_n1072));
  INV_X1    g0872(.A(G128), .ZN(new_n1073));
  INV_X1    g0873(.A(G137), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n255), .B1(new_n764), .B2(new_n1073), .C1(new_n1074), .C2(new_n767), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n780), .B2(G159), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1070), .A2(new_n1072), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n771), .A2(new_n832), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1066), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(new_n741), .B1(new_n299), .B2(new_n835), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n735), .B(new_n1080), .C1(new_n893), .C2(new_n739), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n804), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n406), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n687), .B(new_n1083), .C1(new_n705), .C2(new_n709), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n803), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n897), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n894), .B1(new_n868), .B2(new_n873), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n899), .A2(new_n803), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n894), .B1(new_n1089), .B2(new_n897), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1088), .B1(new_n1090), .B2(new_n893), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n863), .A2(new_n727), .A3(G330), .A4(new_n728), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1088), .B(new_n1092), .C1(new_n1090), .C2(new_n893), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1081), .B1(new_n1096), .B2(new_n970), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n727), .A2(new_n728), .A3(G330), .A4(new_n806), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n898), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1092), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1089), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1085), .B2(new_n1100), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n903), .A2(new_n904), .A3(new_n877), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1032), .B1(new_n1096), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1094), .A2(new_n1095), .A3(new_n1103), .A4(new_n1102), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1097), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(G378));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1103), .ZN(new_n1109));
  INV_X1    g0909(.A(G330), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n883), .B2(new_n887), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n902), .A2(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n893), .A2(new_n894), .B1(new_n886), .B2(new_n900), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n876), .A2(new_n1113), .A3(new_n896), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n307), .A2(new_n669), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n381), .A2(new_n312), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n381), .B2(new_n312), .ZN(new_n1118));
  OR3_X1    g0918(.A1(new_n1117), .A2(new_n1118), .A3(KEYINPUT55), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT55), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(new_n1121), .B(KEYINPUT56), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1112), .A2(new_n1114), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1122), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1109), .B(KEYINPUT57), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n1033), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(KEYINPUT123), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT57), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1109), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT123), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1125), .A2(new_n1132), .A3(new_n1033), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1127), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1122), .A2(new_n738), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n835), .A2(new_n201), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G41), .B(new_n255), .C1(new_n919), .C2(G77), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT121), .Z(new_n1138));
  NOR2_X1   g0938(.A1(new_n771), .A2(new_n207), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n756), .A2(new_n202), .B1(new_n816), .B2(new_n811), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n821), .A2(G97), .B1(new_n776), .B2(new_n383), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1141), .B1(new_n219), .B2(new_n764), .C1(new_n779), .C2(new_n203), .ZN(new_n1142));
  NOR4_X1   g0942(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT58), .Z(new_n1144));
  OAI21_X1  g0944(.A(new_n201), .B1(new_n260), .B2(G41), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n767), .A2(new_n832), .B1(new_n764), .B2(new_n1068), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n771), .A2(new_n1073), .B1(new_n775), .B2(new_n1074), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n780), .C2(G150), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n773), .B2(new_n1067), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT59), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n811), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(KEYINPUT122), .A2(G124), .ZN(new_n1153));
  AOI21_X1  g0953(.A(G33), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1149), .A2(KEYINPUT59), .ZN(new_n1155));
  AOI21_X1  g0955(.A(G41), .B1(new_n757), .B2(G159), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .A4(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1144), .A2(new_n1145), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n734), .B1(new_n1158), .B2(new_n741), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1135), .A2(new_n1136), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1129), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1161), .B1(new_n1162), .B2(new_n971), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1134), .A2(new_n1163), .ZN(G375));
  NOR2_X1   g0964(.A1(new_n1100), .A2(new_n1085), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1089), .B2(new_n1100), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n905), .A2(new_n878), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1168), .A2(new_n1104), .A3(new_n988), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n898), .A2(new_n738), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n811), .A2(new_n465), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1171), .B(new_n932), .C1(G107), .C2(new_n787), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n767), .A2(new_n219), .B1(new_n764), .B2(new_n526), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n262), .B1(new_n773), .B2(new_n206), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n780), .C2(new_n383), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(new_n816), .C2(new_n771), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n756), .A2(new_n202), .B1(new_n1073), .B2(new_n811), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n832), .A2(new_n764), .B1(new_n767), .B2(new_n1067), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n255), .B1(new_n771), .B2(new_n1074), .C1(new_n824), .C2(new_n773), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n201), .B2(new_n779), .C1(new_n288), .C2(new_n775), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1176), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1182), .A2(new_n741), .B1(new_n203), .B2(new_n835), .ZN(new_n1183));
  AND3_X1   g0983(.A1(new_n1170), .A2(new_n735), .A3(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n970), .B(KEYINPUT124), .Z(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1184), .B1(new_n1102), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1169), .A2(new_n1187), .ZN(G381));
  NAND3_X1  g0988(.A1(new_n1134), .A2(new_n1107), .A3(new_n1163), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(G384), .A3(G381), .ZN(new_n1190));
  OR2_X1    g0990(.A1(G393), .A2(G396), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(G387), .A2(G390), .A3(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(KEYINPUT125), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT125), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1193), .A2(new_n1194), .ZN(G407));
  OAI221_X1 g0995(.A(G213), .B1(G343), .B2(new_n1189), .C1(new_n1193), .C2(new_n1194), .ZN(G409));
  XNOR2_X1  g0996(.A(G390), .B(new_n990), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(G393), .A2(G396), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1191), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n968), .A2(new_n989), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT117), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1201), .A2(new_n1202), .A3(new_n946), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G390), .B1(new_n1203), .B2(new_n991), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT126), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1199), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(G390), .A2(new_n1201), .A3(new_n946), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1200), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT61), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n670), .A2(G213), .A3(G2897), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT60), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1032), .B1(new_n1168), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1166), .A2(new_n1167), .A3(KEYINPUT60), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1104), .A3(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1218), .A2(G384), .A3(new_n1187), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G384), .B1(new_n1218), .B2(new_n1187), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1214), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1221), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n1219), .A3(new_n1213), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1107), .B1(new_n1134), .B2(new_n1163), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n670), .A2(G213), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1186), .B1(new_n1109), .B2(new_n988), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1160), .B1(new_n1228), .B2(new_n1129), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1227), .B1(new_n1229), .B2(G378), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1225), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1226), .A2(new_n1230), .A3(new_n1233), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1212), .B(new_n1231), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(G375), .A2(G378), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1230), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1237), .A2(new_n1238), .A3(new_n1232), .ZN(new_n1239));
  OR2_X1    g1039(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1211), .B1(new_n1236), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT63), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1239), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G390), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n992), .B2(new_n993), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1208), .B1(new_n1248), .B2(KEYINPUT126), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n1249), .A2(new_n1206), .B1(new_n1199), .B2(new_n1197), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT61), .B1(new_n1234), .B2(KEYINPUT63), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1246), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1242), .A2(new_n1252), .ZN(G405));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1189), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1211), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1250), .A2(new_n1189), .A3(new_n1237), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n1233), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1256), .A3(new_n1232), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(G402));
endmodule


