//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT5), .ZN(new_n203));
  XNOR2_X1  g002(.A(G141gat), .B(G148gat), .ZN(new_n204));
  AND2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT78), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT78), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT2), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n204), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n212), .B1(G155gat), .B2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(KEYINPUT77), .ZN(new_n214));
  OAI22_X1  g013(.A1(new_n213), .A2(new_n214), .B1(G155gat), .B2(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT79), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n206), .B1(new_n220), .B2(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G141gat), .ZN(new_n222));
  INV_X1    g021(.A(G148gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n224), .B(new_n225), .C1(new_n205), .C2(new_n226), .ZN(new_n227));
  OAI22_X1  g026(.A1(new_n211), .A2(new_n215), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  INV_X1    g028(.A(G120gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT1), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n229), .B2(new_n230), .ZN(new_n232));
  XNOR2_X1  g031(.A(G127gat), .B(G134gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT71), .B(G120gat), .ZN(new_n236));
  OAI211_X1 g035(.A(new_n231), .B(new_n233), .C1(new_n236), .C2(new_n229), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n228), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n203), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT2), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n209), .B1(new_n208), .B2(KEYINPUT2), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n224), .B(new_n225), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n214), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n208), .A2(KEYINPUT77), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n226), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT79), .B(G162gat), .ZN(new_n250));
  INV_X1    g049(.A(G155gat), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT2), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n205), .A2(new_n226), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(new_n204), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n246), .A2(new_n249), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n243), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n228), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n228), .B2(KEYINPUT3), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n255), .A2(KEYINPUT81), .A3(new_n256), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n259), .A2(new_n263), .A3(new_n238), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT82), .ZN(new_n265));
  INV_X1    g064(.A(new_n238), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n255), .A3(KEYINPUT4), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n228), .B2(new_n238), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n267), .A2(new_n269), .A3(new_n240), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n264), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n265), .B1(new_n264), .B2(new_n270), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n242), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274));
  XNOR2_X1  g073(.A(G1gat), .B(G29gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT0), .ZN(new_n276));
  XNOR2_X1  g075(.A(G57gat), .B(G85gat), .ZN(new_n277));
  XOR2_X1   g076(.A(new_n276), .B(new_n277), .Z(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n264), .A2(new_n270), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n279), .B1(new_n280), .B2(new_n203), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n273), .A2(new_n274), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n274), .B1(new_n273), .B2(new_n281), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n202), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n242), .ZN(new_n287));
  INV_X1    g086(.A(new_n272), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n264), .A2(new_n265), .A3(new_n270), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n264), .A2(new_n270), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n291), .A2(KEYINPUT5), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n279), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n273), .A2(new_n281), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT83), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n295), .A2(KEYINPUT84), .A3(new_n283), .A4(new_n282), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n286), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT6), .B(new_n279), .C1(new_n290), .C2(new_n292), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n292), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n278), .B1(new_n273), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(KEYINPUT85), .A3(KEYINPUT6), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n297), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT26), .ZN(new_n309));
  INV_X1    g108(.A(G183gat), .ZN(new_n310));
  INV_X1    g109(.A(G190gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n308), .A2(KEYINPUT26), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n309), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT27), .B(G183gat), .Z(new_n316));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n317));
  NOR3_X1   g116(.A1(new_n316), .A2(new_n317), .A3(G190gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n310), .A2(KEYINPUT69), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G183gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n319), .B1(new_n323), .B2(KEYINPUT27), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n317), .B1(new_n324), .B2(G190gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n318), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n319), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT69), .B(G183gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT27), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT28), .B1(new_n331), .B2(new_n311), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(KEYINPUT70), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n315), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(G169gat), .B2(G176gat), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n306), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT66), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n343));
  NAND3_X1  g142(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n310), .A2(new_n311), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n342), .A2(new_n343), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n344), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT65), .B1(new_n347), .B2(new_n341), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n335), .A2(KEYINPUT66), .A3(new_n337), .A4(new_n306), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n340), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  XOR2_X1   g149(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n351));
  XNOR2_X1  g150(.A(new_n341), .B(KEYINPUT68), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n352), .B(new_n344), .C1(G190gat), .C2(new_n323), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT67), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n335), .A2(new_n354), .A3(new_n306), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n335), .B2(new_n306), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n337), .A2(KEYINPUT25), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n350), .A2(new_n351), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(KEYINPUT75), .B1(new_n334), .B2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n318), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n332), .B2(KEYINPUT70), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n325), .A2(new_n326), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n314), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n351), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n353), .A2(new_n358), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n365), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n360), .A2(new_n361), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n365), .A2(new_n368), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n361), .A2(KEYINPUT29), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT73), .B(G197gat), .ZN(new_n378));
  INV_X1    g177(.A(G204gat), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n378), .A2(new_n379), .ZN(new_n381));
  INV_X1    g180(.A(G211gat), .ZN(new_n382));
  INV_X1    g181(.A(G218gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n380), .A2(new_n381), .B1(KEYINPUT22), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(KEYINPUT74), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n377), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n388), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n376), .A3(new_n386), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n334), .A2(KEYINPUT75), .A3(new_n359), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n369), .B1(new_n365), .B2(new_n368), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n373), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n392), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n365), .A2(new_n368), .A3(new_n361), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(G64gat), .B(G92gat), .ZN(new_n401));
  XOR2_X1   g200(.A(new_n400), .B(new_n401), .Z(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n393), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n373), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n360), .B2(new_n370), .ZN(new_n406));
  INV_X1    g205(.A(new_n398), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n406), .A2(new_n392), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n397), .B1(new_n371), .B2(new_n374), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n402), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n403), .B1(new_n393), .B2(new_n399), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT76), .B1(new_n413), .B2(KEYINPUT30), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT76), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n415), .A3(new_n411), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n305), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(G22gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT31), .B(G50gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n256), .B1(new_n392), .B2(KEYINPUT29), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n228), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n261), .A2(new_n262), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n392), .B1(KEYINPUT29), .B2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G78gat), .B(G106gat), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n425), .B2(new_n427), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n423), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n425), .A2(new_n427), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n428), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n425), .A2(new_n427), .A3(new_n429), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n422), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n365), .A2(new_n368), .A3(new_n266), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT72), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT72), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n365), .A2(new_n368), .A3(new_n440), .A4(new_n266), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n372), .A2(new_n238), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT34), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n266), .B1(new_n365), .B2(new_n368), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(KEYINPUT72), .B2(new_n438), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT34), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n444), .A4(new_n441), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(G71gat), .B(G99gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n443), .A2(new_n445), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT33), .B1(new_n443), .B2(new_n445), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n446), .B(new_n450), .C1(new_n459), .C2(new_n454), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(KEYINPUT32), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n462), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n458), .A2(new_n464), .A3(new_n460), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(KEYINPUT36), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT36), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n458), .A2(new_n464), .A3(new_n460), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n464), .B1(new_n458), .B2(new_n460), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n418), .A2(new_n437), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n408), .A2(new_n409), .A3(new_n402), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(KEYINPUT30), .B2(new_n413), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n413), .A2(KEYINPUT76), .A3(KEYINPUT30), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n415), .B1(new_n410), .B2(new_n411), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT86), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n417), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n267), .A2(new_n269), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n264), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n241), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT87), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n484), .A3(new_n241), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n279), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n239), .A2(new_n241), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n483), .A2(KEYINPUT39), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n488), .A2(KEYINPUT40), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT40), .B1(new_n488), .B2(new_n490), .ZN(new_n492));
  NOR3_X1   g291(.A1(new_n491), .A2(new_n492), .A3(new_n302), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n479), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n437), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n403), .A2(KEYINPUT37), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n404), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n392), .B1(new_n406), .B2(new_n407), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n371), .A2(new_n374), .A3(new_n397), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(KEYINPUT37), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT88), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT38), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT88), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT37), .A4(new_n499), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n497), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n505), .A2(new_n410), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n295), .A2(new_n293), .A3(new_n283), .A4(new_n282), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n393), .A2(new_n399), .A3(KEYINPUT37), .ZN(new_n508));
  INV_X1    g307(.A(new_n496), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n472), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT38), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n506), .A2(new_n304), .A3(new_n507), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n471), .A2(new_n513), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n468), .A2(new_n469), .A3(new_n437), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n305), .A2(new_n515), .A3(new_n417), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n477), .A2(new_n479), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT35), .B1(new_n304), .B2(new_n507), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n514), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT90), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n524), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OR2_X1    g329(.A1(new_n529), .A2(new_n525), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n530), .A2(new_n531), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  XOR2_X1   g331(.A(G43gat), .B(G50gat), .Z(new_n533));
  INV_X1    g332(.A(KEYINPUT15), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n533), .A2(new_n534), .B1(new_n529), .B2(new_n523), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n535), .B(new_n537), .C1(new_n527), .C2(new_n528), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G15gat), .B(G22gat), .ZN(new_n540));
  INV_X1    g339(.A(G1gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT16), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  OAI221_X1 g343(.A(new_n543), .B1(KEYINPUT91), .B2(new_n544), .C1(G1gat), .C2(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT91), .ZN(new_n546));
  XOR2_X1   g345(.A(new_n545), .B(new_n546), .Z(new_n547));
  NOR2_X1   g346(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n547), .B(KEYINPUT92), .Z(new_n549));
  OR2_X1    g348(.A1(new_n539), .A2(KEYINPUT17), .ZN(new_n550));
  AND2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n539), .A2(KEYINPUT17), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT93), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n548), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(KEYINPUT18), .A3(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n539), .B(new_n547), .Z(new_n557));
  XOR2_X1   g356(.A(new_n555), .B(KEYINPUT13), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  INV_X1    g365(.A(G197gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT11), .B(G169gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT89), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT94), .B1(new_n562), .B2(new_n563), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n575), .B(KEYINPUT18), .C1(new_n554), .C2(new_n555), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n556), .A2(new_n560), .A3(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(G85gat), .A2(G92gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT7), .ZN(new_n582));
  NAND2_X1  g381(.A1(G99gat), .A2(G106gat), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(KEYINPUT8), .A2(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G99gat), .B(G106gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  NAND3_X1  g388(.A1(new_n553), .A2(new_n550), .A3(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n539), .A2(new_n589), .ZN(new_n591));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT41), .ZN(new_n594));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  OAI22_X1  g394(.A1(new_n593), .A2(KEYINPUT97), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(KEYINPUT97), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n599), .B(KEYINPUT98), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n598), .B(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n594), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT96), .ZN(new_n603));
  XOR2_X1   g402(.A(G134gat), .B(G162gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(new_n605), .ZN(new_n606));
  AND2_X1   g405(.A1(G71gat), .A2(G78gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G57gat), .B(G64gat), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT9), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G64gat), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n613), .A2(G57gat), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT95), .B(G57gat), .Z(new_n615));
  AOI21_X1  g414(.A(new_n614), .B1(new_n615), .B2(G64gat), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n607), .B1(KEYINPUT9), .B2(new_n608), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(G127gat), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n547), .B1(new_n619), .B2(new_n618), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G155gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(G183gat), .B(G211gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n625), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n606), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G120gat), .B(G148gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n582), .A2(new_n588), .A3(new_n586), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n618), .B1(KEYINPUT99), .B2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n589), .ZN(new_n638));
  INV_X1    g437(.A(G230gat), .ZN(new_n639));
  INV_X1    g438(.A(G233gat), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(new_n643), .B(KEYINPUT100), .Z(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n638), .A2(new_n645), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n589), .A2(new_n645), .A3(new_n618), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n642), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n635), .B1(new_n644), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n644), .A2(new_n650), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n634), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(KEYINPUT101), .A3(new_n634), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n653), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n522), .A2(new_n580), .A3(new_n631), .A4(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n305), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n541), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n518), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n544), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(KEYINPUT103), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT16), .B(G8gat), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT42), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(G1325gat));
  NAND2_X1  g470(.A1(new_n470), .A2(new_n466), .ZN(new_n672));
  OAI21_X1  g471(.A(G15gat), .B1(new_n662), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n468), .A2(new_n469), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(G15gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n673), .B1(new_n662), .B2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n662), .A2(new_n495), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n606), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n681), .B1(new_n514), .B2(new_n521), .ZN(new_n682));
  INV_X1    g481(.A(new_n580), .ZN(new_n683));
  INV_X1    g482(.A(new_n630), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n683), .A2(new_n684), .A3(new_n660), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n305), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n527), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT104), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT45), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n511), .A2(new_n410), .A3(new_n505), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n507), .A2(new_n303), .A3(new_n300), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n495), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n414), .A2(new_n416), .ZN(new_n696));
  AND3_X1   g495(.A1(new_n696), .A2(new_n478), .A3(new_n473), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n478), .B1(new_n696), .B2(new_n473), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n695), .B1(new_n699), .B2(new_n493), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n476), .B1(new_n297), .B2(new_n304), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n672), .B1(new_n701), .B2(new_n495), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n692), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n471), .A2(KEYINPUT105), .A3(new_n513), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT35), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n674), .A2(new_n705), .A3(new_n495), .A4(new_n694), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n699), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n701), .B2(new_n515), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT106), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n710), .B1(new_n517), .B2(new_n520), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n703), .B(new_n704), .C1(new_n709), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n712), .B2(new_n606), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n685), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n305), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n691), .A2(new_n717), .ZN(G1328gat));
  OAI21_X1  g517(.A(G36gat), .B1(new_n716), .B2(new_n518), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n686), .A2(G36gat), .A3(new_n518), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1329gat));
  INV_X1    g521(.A(G43gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n682), .A2(new_n723), .A3(new_n674), .A4(new_n685), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT107), .ZN(new_n725));
  INV_X1    g524(.A(new_n672), .ZN(new_n726));
  AND3_X1   g525(.A1(new_n715), .A2(new_n726), .A3(new_n685), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n729), .A2(KEYINPUT108), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G43gat), .B1(new_n716), .B2(new_n672), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n733), .A2(KEYINPUT108), .A3(new_n729), .A4(new_n725), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n732), .A2(new_n734), .ZN(G1330gat));
  NAND2_X1  g534(.A1(new_n437), .A2(G50gat), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n686), .A2(new_n495), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n716), .A2(new_n736), .B1(G50gat), .B2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT48), .ZN(G1331gat));
  AND4_X1   g538(.A1(new_n683), .A2(new_n712), .A3(new_n631), .A4(new_n660), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n687), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(new_n615), .Z(G1332gat));
  AOI21_X1  g541(.A(new_n518), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT109), .Z(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT110), .ZN(new_n746));
  NOR2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1333gat));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n726), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n675), .A2(G71gat), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n749), .A2(G71gat), .B1(new_n740), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n437), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g553(.A1(new_n660), .A2(new_n584), .A3(new_n687), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n712), .A2(KEYINPUT111), .A3(new_n606), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n580), .A2(new_n684), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(KEYINPUT111), .B1(new_n712), .B2(new_n606), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(new_n760), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(KEYINPUT51), .A3(new_n758), .A4(new_n757), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n755), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n758), .A2(new_n660), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n713), .A2(new_n714), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n584), .B1(new_n766), .B2(new_n687), .ZN(new_n767));
  OR3_X1    g566(.A1(new_n764), .A2(KEYINPUT112), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT112), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(G1336gat));
  NOR3_X1   g569(.A1(new_n661), .A2(G92gat), .A3(new_n518), .ZN(new_n771));
  INV_X1    g570(.A(new_n758), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n700), .A2(new_n692), .A3(new_n702), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT105), .B1(new_n471), .B2(new_n513), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n521), .A2(KEYINPUT106), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n517), .A2(new_n710), .A3(new_n520), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n681), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n772), .B1(new_n779), .B2(KEYINPUT111), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n780), .B2(new_n762), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n759), .A2(new_n756), .A3(new_n760), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n771), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g582(.A1(new_n713), .A2(new_n714), .A3(new_n518), .A4(new_n765), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n585), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n783), .B(new_n786), .C1(new_n787), .C2(KEYINPUT52), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n784), .B2(new_n585), .ZN(new_n790));
  INV_X1    g589(.A(new_n771), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n761), .B2(new_n763), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n789), .B(new_n790), .C1(new_n792), .C2(new_n785), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n788), .A2(new_n793), .ZN(G1337gat));
  INV_X1    g593(.A(G99gat), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n766), .A2(new_n726), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(KEYINPUT114), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(KEYINPUT114), .B2(new_n796), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n660), .A2(new_n795), .A3(new_n674), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT115), .Z(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n781), .B2(new_n782), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(G1338gat));
  INV_X1    g601(.A(G106gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n660), .A2(new_n803), .A3(new_n437), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT116), .Z(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n761), .B2(new_n763), .ZN(new_n807));
  NOR4_X1   g606(.A1(new_n713), .A2(new_n714), .A3(new_n495), .A4(new_n765), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n808), .A2(new_n803), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n808), .B2(new_n803), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(KEYINPUT53), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT53), .B(new_n812), .C1(new_n807), .C2(new_n809), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(G1339gat));
  NAND3_X1  g615(.A1(new_n683), .A2(new_n631), .A3(new_n661), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n635), .B1(new_n649), .B2(KEYINPUT54), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n649), .A2(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n646), .A2(new_n641), .A3(new_n647), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(KEYINPUT55), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n606), .A2(new_n659), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n557), .A2(new_n559), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT118), .Z(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n555), .B2(new_n554), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n570), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n579), .A2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(KEYINPUT119), .B1(new_n825), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n659), .A2(new_n823), .A3(new_n824), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n577), .A2(new_n578), .B1(new_n570), .B2(new_n828), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n606), .ZN(new_n835));
  AOI22_X1  g634(.A1(new_n580), .A2(new_n832), .B1(new_n660), .B2(new_n834), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n831), .B(new_n835), .C1(new_n836), .C2(new_n606), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n818), .B1(new_n837), .B2(new_n630), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n305), .A3(new_n437), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n699), .A2(new_n675), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g640(.A1(new_n841), .A2(new_n683), .B1(KEYINPUT120), .B2(G113gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(KEYINPUT120), .A2(G113gat), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT121), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n842), .B(new_n844), .ZN(G1340gat));
  OR3_X1    g644(.A1(new_n841), .A2(new_n236), .A3(new_n661), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n230), .B1(new_n841), .B2(new_n661), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n847), .B1(new_n846), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1341gat));
  NOR2_X1   g650(.A1(new_n841), .A2(new_n630), .ZN(new_n852));
  XOR2_X1   g651(.A(new_n852), .B(G127gat), .Z(G1342gat));
  NOR2_X1   g652(.A1(new_n681), .A2(new_n699), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n675), .A2(G134gat), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n839), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XOR2_X1   g655(.A(new_n856), .B(KEYINPUT56), .Z(new_n857));
  OAI21_X1  g656(.A(G134gat), .B1(new_n841), .B2(new_n681), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1343gat));
  NOR2_X1   g658(.A1(new_n726), .A2(new_n305), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n518), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n831), .A2(new_n835), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n580), .A2(new_n832), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n660), .A2(new_n834), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n606), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n630), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n817), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT57), .B1(new_n868), .B2(new_n437), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n838), .A2(new_n870), .A3(new_n495), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n580), .B(new_n862), .C1(new_n869), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT123), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(KEYINPUT57), .A3(new_n437), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n838), .B2(new_n495), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n861), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(new_n580), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n873), .A2(G141gat), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n838), .A2(new_n495), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n862), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n881), .A2(G141gat), .A3(new_n683), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(KEYINPUT58), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n879), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n222), .B1(new_n876), .B2(new_n580), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT58), .B1(new_n885), .B2(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1344gat));
  INV_X1    g686(.A(new_n881), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n888), .A2(new_n223), .A3(new_n660), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n661), .B1(new_n861), .B2(new_n891), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n836), .A2(new_n606), .B1(new_n830), .B2(new_n825), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n818), .B1(new_n893), .B2(new_n630), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n870), .B1(new_n894), .B2(new_n495), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OAI221_X1 g695(.A(new_n892), .B1(new_n891), .B2(new_n861), .C1(new_n896), .C2(new_n871), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n890), .B1(new_n897), .B2(G148gat), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT59), .B(new_n223), .C1(new_n876), .C2(new_n660), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n889), .B1(new_n898), .B2(new_n899), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n888), .A2(new_n251), .A3(new_n684), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n876), .A2(new_n684), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n901), .B1(new_n902), .B2(new_n251), .ZN(G1346gat));
  NAND4_X1  g702(.A1(new_n880), .A2(new_n250), .A3(new_n854), .A4(new_n860), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n876), .A2(new_n606), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n250), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n518), .A2(new_n687), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n838), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n515), .ZN(new_n910));
  INV_X1    g709(.A(G169gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n910), .A2(new_n911), .A3(new_n683), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n909), .A2(new_n515), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT125), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n580), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n912), .B1(new_n915), .B2(new_n911), .ZN(G1348gat));
  INV_X1    g715(.A(G176gat), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n914), .A2(new_n917), .A3(new_n660), .ZN(new_n918));
  OAI21_X1  g717(.A(G176gat), .B1(new_n910), .B2(new_n661), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(G1349gat));
  AOI21_X1  g719(.A(new_n329), .B1(new_n913), .B2(new_n684), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT60), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n913), .A2(new_n684), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n922), .B(new_n923), .C1(new_n316), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n316), .ZN(new_n926));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n926), .B2(new_n921), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n914), .A2(new_n311), .A3(new_n606), .ZN(new_n929));
  OAI21_X1  g728(.A(G190gat), .B1(new_n910), .B2(new_n681), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT61), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1351gat));
  NOR4_X1   g732(.A1(new_n838), .A2(new_n495), .A3(new_n726), .A4(new_n908), .ZN(new_n934));
  AOI21_X1  g733(.A(G197gat), .B1(new_n934), .B2(new_n580), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n908), .A2(new_n726), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n874), .B2(new_n895), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n683), .A2(new_n567), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n935), .B1(new_n938), .B2(new_n939), .ZN(G1352gat));
  XNOR2_X1  g739(.A(KEYINPUT126), .B(G204gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n934), .A2(new_n660), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n938), .A2(new_n660), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n943), .B(new_n944), .C1(new_n945), .C2(new_n941), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n934), .A2(new_n382), .A3(new_n684), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n938), .A2(new_n684), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n948), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n949));
  AOI21_X1  g748(.A(KEYINPUT63), .B1(new_n948), .B2(G211gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(G1354gat));
  AOI21_X1  g750(.A(new_n383), .B1(new_n938), .B2(new_n606), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n934), .A2(new_n383), .A3(new_n606), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT127), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT127), .B1(new_n952), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1355gat));
endmodule


