

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U562 ( .A(n745), .ZN(n725) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n658) );
  XOR2_X1 U564 ( .A(KEYINPUT27), .B(n716), .Z(n528) );
  AND2_X1 U565 ( .A1(n823), .A2(n822), .ZN(n529) );
  OR2_X1 U566 ( .A1(n744), .A2(n743), .ZN(n774) );
  NOR2_X1 U567 ( .A1(n785), .A2(n784), .ZN(n786) );
  AND2_X1 U568 ( .A1(n821), .A2(n830), .ZN(n822) );
  INV_X1 U569 ( .A(G651), .ZN(n547) );
  NOR2_X1 U570 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X2 U571 ( .A1(n644), .A2(n547), .ZN(n662) );
  XNOR2_X1 U572 ( .A(KEYINPUT1), .B(n549), .ZN(n654) );
  NAND2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n530) );
  XNOR2_X1 U574 ( .A(n530), .B(KEYINPUT65), .ZN(n892) );
  NAND2_X1 U575 ( .A1(n892), .A2(G114), .ZN(n533) );
  INV_X1 U576 ( .A(G2105), .ZN(n535) );
  NOR2_X1 U577 ( .A1(n535), .A2(G2104), .ZN(n531) );
  XNOR2_X1 U578 ( .A(n531), .B(KEYINPUT64), .ZN(n893) );
  NAND2_X1 U579 ( .A1(G126), .A2(n893), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n540) );
  OR2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XNOR2_X2 U582 ( .A(KEYINPUT17), .B(n534), .ZN(n887) );
  NAND2_X1 U583 ( .A1(G138), .A2(n887), .ZN(n537) );
  AND2_X1 U584 ( .A1(n535), .A2(G2104), .ZN(n888) );
  NAND2_X1 U585 ( .A1(G102), .A2(n888), .ZN(n536) );
  NAND2_X1 U586 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U587 ( .A(KEYINPUT93), .B(n538), .Z(n539) );
  NOR2_X1 U588 ( .A1(n540), .A2(n539), .ZN(G164) );
  AND2_X1 U589 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U590 ( .A(G132), .ZN(G219) );
  INV_X1 U591 ( .A(G82), .ZN(G220) );
  INV_X1 U592 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U593 ( .A(KEYINPUT82), .B(KEYINPUT7), .ZN(n557) );
  NAND2_X1 U594 ( .A1(n658), .A2(G89), .ZN(n541) );
  XNOR2_X1 U595 ( .A(n541), .B(KEYINPUT4), .ZN(n544) );
  XNOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .ZN(n542) );
  XNOR2_X1 U597 ( .A(n542), .B(KEYINPUT67), .ZN(n644) );
  NAND2_X1 U598 ( .A1(G76), .A2(n662), .ZN(n543) );
  NAND2_X1 U599 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U600 ( .A(n545), .B(KEYINPUT5), .ZN(n555) );
  XNOR2_X1 U601 ( .A(KEYINPUT6), .B(KEYINPUT81), .ZN(n553) );
  NOR2_X1 U602 ( .A1(G651), .A2(n644), .ZN(n653) );
  NAND2_X1 U603 ( .A1(n653), .A2(G51), .ZN(n546) );
  XNOR2_X1 U604 ( .A(n546), .B(KEYINPUT80), .ZN(n551) );
  NOR2_X1 U605 ( .A1(G543), .A2(n547), .ZN(n548) );
  XOR2_X1 U606 ( .A(KEYINPUT68), .B(n548), .Z(n549) );
  NAND2_X1 U607 ( .A1(G63), .A2(n654), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U609 ( .A(n553), .B(n552), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n557), .B(n556), .ZN(G168) );
  XOR2_X1 U612 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  XOR2_X1 U613 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n559) );
  NAND2_X1 U614 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n559), .B(n558), .ZN(G223) );
  INV_X1 U616 ( .A(G223), .ZN(n840) );
  NAND2_X1 U617 ( .A1(n840), .A2(G567), .ZN(n560) );
  XOR2_X1 U618 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  XOR2_X1 U619 ( .A(G860), .B(KEYINPUT77), .Z(n604) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n562) );
  NAND2_X1 U621 ( .A1(G56), .A2(n654), .ZN(n561) );
  XNOR2_X1 U622 ( .A(n562), .B(n561), .ZN(n571) );
  NAND2_X1 U623 ( .A1(n658), .A2(G81), .ZN(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT12), .B(n563), .ZN(n566) );
  NAND2_X1 U625 ( .A1(n662), .A2(G68), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT75), .B(n564), .Z(n565) );
  NAND2_X1 U627 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U628 ( .A(n567), .B(KEYINPUT13), .ZN(n569) );
  NAND2_X1 U629 ( .A1(G43), .A2(n653), .ZN(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT76), .B(n572), .Z(n982) );
  INV_X1 U632 ( .A(n982), .ZN(n573) );
  NAND2_X1 U633 ( .A1(n604), .A2(n573), .ZN(G153) );
  NAND2_X1 U634 ( .A1(G52), .A2(n653), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT70), .B(n574), .Z(n579) );
  NAND2_X1 U636 ( .A1(G90), .A2(n658), .ZN(n576) );
  NAND2_X1 U637 ( .A1(G77), .A2(n662), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U640 ( .A1(n579), .A2(n578), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G64), .A2(n654), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G301), .A2(G868), .ZN(n582) );
  XNOR2_X1 U644 ( .A(n582), .B(KEYINPUT78), .ZN(n592) );
  INV_X1 U645 ( .A(G868), .ZN(n674) );
  NAND2_X1 U646 ( .A1(n653), .A2(G54), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G92), .A2(n658), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G79), .A2(n662), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G66), .A2(n654), .ZN(n585) );
  XNOR2_X1 U651 ( .A(KEYINPUT79), .B(n585), .ZN(n586) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n590), .Z(n987) );
  NAND2_X1 U655 ( .A1(n674), .A2(n987), .ZN(n591) );
  NAND2_X1 U656 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G53), .A2(n653), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G65), .A2(n654), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(KEYINPUT72), .B(n595), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G78), .A2(n662), .ZN(n596) );
  XNOR2_X1 U662 ( .A(KEYINPUT71), .B(n596), .ZN(n597) );
  NOR2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U664 ( .A1(n658), .A2(G91), .ZN(n599) );
  NAND2_X1 U665 ( .A1(n600), .A2(n599), .ZN(G299) );
  NAND2_X1 U666 ( .A1(G868), .A2(G286), .ZN(n602) );
  NAND2_X1 U667 ( .A1(G299), .A2(n674), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(G297) );
  INV_X1 U669 ( .A(G559), .ZN(n603) );
  NOR2_X1 U670 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U671 ( .A1(n987), .A2(n605), .ZN(n606) );
  XOR2_X1 U672 ( .A(KEYINPUT16), .B(n606), .Z(G148) );
  NOR2_X1 U673 ( .A1(n982), .A2(G868), .ZN(n607) );
  XOR2_X1 U674 ( .A(KEYINPUT83), .B(n607), .Z(n610) );
  INV_X1 U675 ( .A(n987), .ZN(n908) );
  NAND2_X1 U676 ( .A1(G868), .A2(n908), .ZN(n608) );
  NOR2_X1 U677 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U678 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U679 ( .A1(n893), .A2(G123), .ZN(n611) );
  XNOR2_X1 U680 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n888), .A2(G99), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U683 ( .A1(G135), .A2(n887), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G111), .A2(n892), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n932) );
  XNOR2_X1 U687 ( .A(n932), .B(G2096), .ZN(n619) );
  INV_X1 U688 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U690 ( .A1(G559), .A2(n908), .ZN(n620) );
  XNOR2_X1 U691 ( .A(n620), .B(n982), .ZN(n671) );
  NOR2_X1 U692 ( .A1(G860), .A2(n671), .ZN(n630) );
  NAND2_X1 U693 ( .A1(G67), .A2(n654), .ZN(n621) );
  XOR2_X1 U694 ( .A(KEYINPUT85), .B(n621), .Z(n623) );
  NAND2_X1 U695 ( .A1(n653), .A2(G55), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U697 ( .A(KEYINPUT86), .B(n624), .ZN(n629) );
  NAND2_X1 U698 ( .A1(G80), .A2(n662), .ZN(n625) );
  XNOR2_X1 U699 ( .A(n625), .B(KEYINPUT84), .ZN(n627) );
  NAND2_X1 U700 ( .A1(n658), .A2(G93), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n628) );
  OR2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n673) );
  XOR2_X1 U703 ( .A(n630), .B(n673), .Z(G145) );
  NAND2_X1 U704 ( .A1(G61), .A2(n654), .ZN(n637) );
  NAND2_X1 U705 ( .A1(G48), .A2(n653), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G86), .A2(n658), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n662), .A2(G73), .ZN(n633) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U710 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  XOR2_X1 U712 ( .A(KEYINPUT89), .B(n638), .Z(G305) );
  NAND2_X1 U713 ( .A1(G74), .A2(G651), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n639), .B(KEYINPUT88), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G49), .A2(n653), .ZN(n640) );
  XOR2_X1 U716 ( .A(KEYINPUT87), .B(n640), .Z(n641) );
  NAND2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n654), .A2(n643), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n644), .A2(G87), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U721 ( .A1(G88), .A2(n658), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G75), .A2(n662), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G50), .A2(n653), .ZN(n650) );
  NAND2_X1 U725 ( .A1(G62), .A2(n654), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U727 ( .A1(n652), .A2(n651), .ZN(G166) );
  NAND2_X1 U728 ( .A1(G47), .A2(n653), .ZN(n656) );
  NAND2_X1 U729 ( .A1(G60), .A2(n654), .ZN(n655) );
  NAND2_X1 U730 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U731 ( .A(KEYINPUT69), .B(n657), .Z(n661) );
  NAND2_X1 U732 ( .A1(G85), .A2(n658), .ZN(n659) );
  XOR2_X1 U733 ( .A(KEYINPUT66), .B(n659), .Z(n660) );
  NOR2_X1 U734 ( .A1(n661), .A2(n660), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n662), .A2(G72), .ZN(n663) );
  NAND2_X1 U736 ( .A1(n664), .A2(n663), .ZN(G290) );
  XOR2_X1 U737 ( .A(n673), .B(G305), .Z(n670) );
  XNOR2_X1 U738 ( .A(KEYINPUT90), .B(KEYINPUT19), .ZN(n666) );
  XNOR2_X1 U739 ( .A(G288), .B(G166), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U741 ( .A(n667), .B(G290), .Z(n668) );
  XNOR2_X1 U742 ( .A(G299), .B(n668), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n670), .B(n669), .ZN(n907) );
  XNOR2_X1 U744 ( .A(n671), .B(n907), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n672), .A2(G868), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U747 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT91), .ZN(n678) );
  XNOR2_X1 U750 ( .A(KEYINPUT20), .B(n678), .ZN(n679) );
  NAND2_X1 U751 ( .A1(n679), .A2(G2090), .ZN(n680) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U753 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n682) );
  NOR2_X1 U756 ( .A1(G237), .A2(n682), .ZN(n683) );
  XNOR2_X1 U757 ( .A(KEYINPUT92), .B(n683), .ZN(n684) );
  NAND2_X1 U758 ( .A1(n684), .A2(G108), .ZN(n929) );
  NAND2_X1 U759 ( .A1(n929), .A2(G567), .ZN(n689) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n685) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n685), .Z(n686) );
  NOR2_X1 U762 ( .A1(G218), .A2(n686), .ZN(n687) );
  NAND2_X1 U763 ( .A1(G96), .A2(n687), .ZN(n930) );
  NAND2_X1 U764 ( .A1(n930), .A2(G2106), .ZN(n688) );
  NAND2_X1 U765 ( .A1(n689), .A2(n688), .ZN(n845) );
  NAND2_X1 U766 ( .A1(G483), .A2(G661), .ZN(n690) );
  NOR2_X1 U767 ( .A1(n845), .A2(n690), .ZN(n842) );
  NAND2_X1 U768 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(n887), .A2(G137), .ZN(n693) );
  NAND2_X1 U770 ( .A1(G101), .A2(n888), .ZN(n691) );
  XOR2_X1 U771 ( .A(KEYINPUT23), .B(n691), .Z(n692) );
  NAND2_X1 U772 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U773 ( .A1(n892), .A2(G113), .ZN(n695) );
  NAND2_X1 U774 ( .A1(G125), .A2(n893), .ZN(n694) );
  NAND2_X1 U775 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U776 ( .A1(n697), .A2(n696), .ZN(G160) );
  INV_X1 U777 ( .A(G166), .ZN(G303) );
  INV_X1 U778 ( .A(G301), .ZN(G171) );
  INV_X1 U779 ( .A(G1996), .ZN(n699) );
  NOR2_X2 U780 ( .A1(G164), .A2(G1384), .ZN(n809) );
  NAND2_X1 U781 ( .A1(G160), .A2(G40), .ZN(n808) );
  INV_X1 U782 ( .A(n808), .ZN(n698) );
  NAND2_X2 U783 ( .A1(n809), .A2(n698), .ZN(n745) );
  OR2_X1 U784 ( .A1(n699), .A2(n745), .ZN(n700) );
  XNOR2_X1 U785 ( .A(n700), .B(KEYINPUT26), .ZN(n702) );
  NAND2_X1 U786 ( .A1(KEYINPUT26), .A2(G1341), .ZN(n701) );
  OR2_X1 U787 ( .A1(n725), .A2(n701), .ZN(n705) );
  NAND2_X1 U788 ( .A1(n702), .A2(n705), .ZN(n704) );
  INV_X1 U789 ( .A(KEYINPUT99), .ZN(n703) );
  NAND2_X1 U790 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U791 ( .A1(n705), .A2(KEYINPUT99), .ZN(n706) );
  NAND2_X1 U792 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U793 ( .A1(n982), .A2(n708), .ZN(n712) );
  NAND2_X1 U794 ( .A1(G1348), .A2(n745), .ZN(n710) );
  NAND2_X1 U795 ( .A1(G2067), .A2(n725), .ZN(n709) );
  NAND2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n713) );
  NOR2_X1 U797 ( .A1(n987), .A2(n713), .ZN(n711) );
  NOR2_X1 U798 ( .A1(n712), .A2(n711), .ZN(n715) );
  AND2_X1 U799 ( .A1(n987), .A2(n713), .ZN(n714) );
  NOR2_X1 U800 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U801 ( .A1(n725), .A2(G2072), .ZN(n716) );
  NAND2_X1 U802 ( .A1(G1956), .A2(n745), .ZN(n717) );
  NAND2_X1 U803 ( .A1(n528), .A2(n717), .ZN(n720) );
  NOR2_X1 U804 ( .A1(G299), .A2(n720), .ZN(n718) );
  NOR2_X1 U805 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U806 ( .A1(G299), .A2(n720), .ZN(n721) );
  XOR2_X1 U807 ( .A(KEYINPUT28), .B(n721), .Z(n722) );
  NOR2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U809 ( .A(n724), .B(KEYINPUT29), .ZN(n729) );
  XOR2_X1 U810 ( .A(G1961), .B(KEYINPUT98), .Z(n1025) );
  NAND2_X1 U811 ( .A1(n1025), .A2(n745), .ZN(n727) );
  XNOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .ZN(n959) );
  NAND2_X1 U813 ( .A1(n725), .A2(n959), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n727), .A2(n726), .ZN(n735) );
  NAND2_X1 U815 ( .A1(G171), .A2(n735), .ZN(n728) );
  NAND2_X1 U816 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U817 ( .A(n730), .B(KEYINPUT100), .ZN(n753) );
  NAND2_X1 U818 ( .A1(G8), .A2(n745), .ZN(n784) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n784), .ZN(n741) );
  NOR2_X1 U820 ( .A1(n745), .A2(G2084), .ZN(n731) );
  XNOR2_X1 U821 ( .A(n731), .B(KEYINPUT97), .ZN(n739) );
  NAND2_X1 U822 ( .A1(G8), .A2(n739), .ZN(n732) );
  NOR2_X1 U823 ( .A1(n741), .A2(n732), .ZN(n733) );
  XOR2_X1 U824 ( .A(KEYINPUT30), .B(n733), .Z(n734) );
  NOR2_X1 U825 ( .A1(G168), .A2(n734), .ZN(n737) );
  NOR2_X1 U826 ( .A1(G171), .A2(n735), .ZN(n736) );
  NOR2_X1 U827 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U828 ( .A(KEYINPUT31), .B(n738), .Z(n751) );
  AND2_X1 U829 ( .A1(n753), .A2(n751), .ZN(n744) );
  INV_X1 U830 ( .A(n739), .ZN(n740) );
  AND2_X1 U831 ( .A1(G8), .A2(n740), .ZN(n742) );
  OR2_X1 U832 ( .A1(n742), .A2(n741), .ZN(n743) );
  INV_X1 U833 ( .A(G8), .ZN(n750) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n784), .ZN(n747) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n745), .ZN(n746) );
  NOR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n748), .A2(G303), .ZN(n749) );
  OR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n754) );
  AND2_X1 U839 ( .A1(n751), .A2(n754), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n757) );
  INV_X1 U841 ( .A(n754), .ZN(n755) );
  OR2_X1 U842 ( .A1(n755), .A2(G286), .ZN(n756) );
  NAND2_X1 U843 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U844 ( .A(n758), .B(KEYINPUT32), .ZN(n776) );
  NAND2_X1 U845 ( .A1(n774), .A2(n776), .ZN(n761) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U847 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  XNOR2_X1 U849 ( .A(n762), .B(KEYINPUT104), .ZN(n763) );
  NAND2_X1 U850 ( .A1(n763), .A2(n784), .ZN(n764) );
  XNOR2_X1 U851 ( .A(n764), .B(KEYINPUT105), .ZN(n768) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n765) );
  XOR2_X1 U853 ( .A(n765), .B(KEYINPUT24), .Z(n766) );
  NOR2_X1 U854 ( .A1(n784), .A2(n766), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n791) );
  INV_X1 U856 ( .A(KEYINPUT103), .ZN(n770) );
  NOR2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NAND2_X1 U858 ( .A1(n993), .A2(KEYINPUT33), .ZN(n769) );
  NAND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n772) );
  NAND2_X1 U860 ( .A1(n993), .A2(KEYINPUT103), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n784), .A2(n773), .ZN(n788) );
  AND2_X1 U863 ( .A1(n774), .A2(n770), .ZN(n775) );
  NAND2_X1 U864 ( .A1(n776), .A2(n775), .ZN(n781) );
  NOR2_X1 U865 ( .A1(G1971), .A2(G303), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT101), .B(n777), .Z(n778) );
  NOR2_X1 U867 ( .A1(n778), .A2(n993), .ZN(n779) );
  OR2_X1 U868 ( .A1(KEYINPUT103), .A2(n779), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G288), .A2(G1976), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT102), .ZN(n994) );
  NAND2_X1 U872 ( .A1(n783), .A2(n994), .ZN(n785) );
  NOR2_X1 U873 ( .A1(KEYINPUT33), .A2(n786), .ZN(n787) );
  NOR2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U875 ( .A(G1981), .B(G305), .Z(n984) );
  NAND2_X1 U876 ( .A1(n789), .A2(n984), .ZN(n790) );
  NAND2_X1 U877 ( .A1(n791), .A2(n790), .ZN(n823) );
  NAND2_X1 U878 ( .A1(G131), .A2(n887), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G95), .A2(n888), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U881 ( .A1(n892), .A2(G107), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G119), .A2(n893), .ZN(n794) );
  NAND2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n901) );
  INV_X1 U885 ( .A(G1991), .ZN(n957) );
  NOR2_X1 U886 ( .A1(n901), .A2(n957), .ZN(n807) );
  NAND2_X1 U887 ( .A1(n892), .A2(G117), .ZN(n804) );
  NAND2_X1 U888 ( .A1(G141), .A2(n887), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G129), .A2(n893), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n888), .A2(G105), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT38), .B(n800), .Z(n801) );
  NOR2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U895 ( .A(KEYINPUT95), .B(n805), .Z(n872) );
  AND2_X1 U896 ( .A1(n872), .A2(G1996), .ZN(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n939) );
  NOR2_X1 U898 ( .A1(n809), .A2(n808), .ZN(n835) );
  XOR2_X1 U899 ( .A(n835), .B(KEYINPUT96), .Z(n810) );
  NOR2_X1 U900 ( .A1(n939), .A2(n810), .ZN(n827) );
  INV_X1 U901 ( .A(n827), .ZN(n821) );
  NAND2_X1 U902 ( .A1(G140), .A2(n887), .ZN(n812) );
  NAND2_X1 U903 ( .A1(G104), .A2(n888), .ZN(n811) );
  NAND2_X1 U904 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT34), .B(n813), .ZN(n819) );
  NAND2_X1 U906 ( .A1(n892), .A2(G116), .ZN(n815) );
  NAND2_X1 U907 ( .A1(G128), .A2(n893), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U909 ( .A(KEYINPUT35), .B(n816), .Z(n817) );
  XNOR2_X1 U910 ( .A(KEYINPUT94), .B(n817), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U912 ( .A(KEYINPUT36), .B(n820), .ZN(n904) );
  XNOR2_X1 U913 ( .A(G2067), .B(KEYINPUT37), .ZN(n832) );
  NOR2_X1 U914 ( .A1(n904), .A2(n832), .ZN(n937) );
  NAND2_X1 U915 ( .A1(n835), .A2(n937), .ZN(n830) );
  XNOR2_X1 U916 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U917 ( .A1(n998), .A2(n835), .ZN(n824) );
  NAND2_X1 U918 ( .A1(n529), .A2(n824), .ZN(n838) );
  NOR2_X1 U919 ( .A1(G1996), .A2(n872), .ZN(n950) );
  AND2_X1 U920 ( .A1(n957), .A2(n901), .ZN(n933) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n933), .A2(n825), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n950), .A2(n828), .ZN(n829) );
  XNOR2_X1 U925 ( .A(KEYINPUT39), .B(n829), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n831), .A2(n830), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n832), .A2(n904), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n833), .B(KEYINPUT106), .ZN(n948) );
  NAND2_X1 U929 ( .A1(n834), .A2(n948), .ZN(n836) );
  NAND2_X1 U930 ( .A1(n836), .A2(n835), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U932 ( .A(KEYINPUT40), .B(n839), .ZN(G329) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U935 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G1), .A2(G3), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U938 ( .A(n844), .B(KEYINPUT108), .ZN(G188) );
  INV_X1 U939 ( .A(n845), .ZN(G319) );
  XOR2_X1 U940 ( .A(KEYINPUT109), .B(G2078), .Z(n847) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2084), .ZN(n846) );
  XNOR2_X1 U942 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U943 ( .A(n848), .B(G2100), .Z(n850) );
  XNOR2_X1 U944 ( .A(G2072), .B(G2090), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n852) );
  XNOR2_X1 U947 ( .A(G2678), .B(KEYINPUT42), .ZN(n851) );
  XNOR2_X1 U948 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U949 ( .A(n854), .B(n853), .Z(G227) );
  XNOR2_X1 U950 ( .A(G1966), .B(KEYINPUT41), .ZN(n864) );
  XOR2_X1 U951 ( .A(G1961), .B(G1976), .Z(n856) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1981), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U954 ( .A(G1971), .B(G1956), .Z(n858) );
  XNOR2_X1 U955 ( .A(G1996), .B(G1991), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U957 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U958 ( .A(G2474), .B(KEYINPUT110), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n863) );
  XNOR2_X1 U960 ( .A(n864), .B(n863), .ZN(G229) );
  NAND2_X1 U961 ( .A1(n893), .A2(G124), .ZN(n865) );
  XNOR2_X1 U962 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U963 ( .A1(n888), .A2(G100), .ZN(n866) );
  NAND2_X1 U964 ( .A1(n867), .A2(n866), .ZN(n871) );
  NAND2_X1 U965 ( .A1(G136), .A2(n887), .ZN(n869) );
  NAND2_X1 U966 ( .A1(G112), .A2(n892), .ZN(n868) );
  NAND2_X1 U967 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U968 ( .A1(n871), .A2(n870), .ZN(G162) );
  XOR2_X1 U969 ( .A(n932), .B(G162), .Z(n874) );
  XOR2_X1 U970 ( .A(G160), .B(n872), .Z(n873) );
  XNOR2_X1 U971 ( .A(n874), .B(n873), .ZN(n886) );
  XOR2_X1 U972 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n884) );
  NAND2_X1 U973 ( .A1(n892), .A2(G115), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G127), .A2(n893), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n877), .B(KEYINPUT47), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G139), .A2(n887), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n882) );
  NAND2_X1 U979 ( .A1(n888), .A2(G103), .ZN(n880) );
  XOR2_X1 U980 ( .A(KEYINPUT112), .B(n880), .Z(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n940) );
  XNOR2_X1 U982 ( .A(n940), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U983 ( .A(n884), .B(n883), .ZN(n885) );
  XOR2_X1 U984 ( .A(n886), .B(n885), .Z(n903) );
  NAND2_X1 U985 ( .A1(G142), .A2(n887), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G106), .A2(n888), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n891), .B(KEYINPUT45), .ZN(n898) );
  NAND2_X1 U989 ( .A1(n892), .A2(G118), .ZN(n895) );
  NAND2_X1 U990 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(KEYINPUT111), .B(n896), .ZN(n897) );
  NAND2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(G164), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U997 ( .A(n905), .B(n904), .Z(n906) );
  NOR2_X1 U998 ( .A1(G37), .A2(n906), .ZN(G395) );
  XNOR2_X1 U999 ( .A(G286), .B(n907), .ZN(n910) );
  XNOR2_X1 U1000 ( .A(G171), .B(n908), .ZN(n909) );
  XNOR2_X1 U1001 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1002 ( .A(n982), .B(n911), .Z(n912) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n912), .ZN(n913) );
  XNOR2_X1 U1004 ( .A(KEYINPUT114), .B(n913), .ZN(G397) );
  XOR2_X1 U1005 ( .A(KEYINPUT107), .B(G2446), .Z(n915) );
  XNOR2_X1 U1006 ( .A(G2435), .B(G2438), .ZN(n914) );
  XNOR2_X1 U1007 ( .A(n915), .B(n914), .ZN(n922) );
  XOR2_X1 U1008 ( .A(G2451), .B(G2430), .Z(n917) );
  XNOR2_X1 U1009 ( .A(G2454), .B(G2427), .ZN(n916) );
  XNOR2_X1 U1010 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1011 ( .A(n918), .B(G2443), .Z(n920) );
  XNOR2_X1 U1012 ( .A(G1341), .B(G1348), .ZN(n919) );
  XNOR2_X1 U1013 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(n922), .B(n921), .ZN(n923) );
  NAND2_X1 U1015 ( .A1(n923), .A2(G14), .ZN(n931) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n931), .ZN(n926) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n924) );
  XNOR2_X1 U1018 ( .A(KEYINPUT49), .B(n924), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n928) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n927) );
  NAND2_X1 U1021 ( .A1(n928), .A2(n927), .ZN(G225) );
  XNOR2_X1 U1022 ( .A(KEYINPUT115), .B(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G120), .ZN(G236) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(G96), .ZN(G221) );
  INV_X1 U1027 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(G325) );
  INV_X1 U1029 ( .A(G325), .ZN(G261) );
  INV_X1 U1030 ( .A(n931), .ZN(G401) );
  XNOR2_X1 U1031 ( .A(G160), .B(G2084), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n946) );
  XOR2_X1 U1036 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1038 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n943), .Z(n944) );
  XNOR2_X1 U1040 ( .A(KEYINPUT116), .B(n944), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n953) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(KEYINPUT51), .B(n951), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  INV_X1 U1048 ( .A(KEYINPUT55), .ZN(n978) );
  NAND2_X1 U1049 ( .A1(n955), .A2(n978), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n956), .A2(G29), .ZN(n1041) );
  XNOR2_X1 U1051 ( .A(G2090), .B(G35), .ZN(n971) );
  XNOR2_X1 U1052 ( .A(G25), .B(n957), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G28), .ZN(n968) );
  XNOR2_X1 U1054 ( .A(G27), .B(n959), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(G1996), .B(G32), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(G2067), .B(G26), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G2072), .B(G33), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(KEYINPUT117), .B(n962), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n969), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT118), .B(n972), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(G34), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G2084), .B(n974), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n978), .B(n977), .ZN(n980) );
  INV_X1 U1071 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n981), .ZN(n1039) );
  XNOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XNOR2_X1 U1075 ( .A(G1341), .B(n982), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(n983), .B(KEYINPUT123), .ZN(n1007) );
  XNOR2_X1 U1077 ( .A(G1966), .B(G168), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1079 ( .A(KEYINPUT57), .B(n986), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT120), .ZN(n988) );
  XNOR2_X1 U1081 ( .A(n988), .B(n987), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G1961), .B(G301), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n1005) );
  INV_X1 U1085 ( .A(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1087 ( .A(KEYINPUT121), .B(n996), .Z(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(G299), .B(G1956), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G303), .B(G1971), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(KEYINPUT122), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1037) );
  INV_X1 U1097 ( .A(G16), .ZN(n1035) );
  XOR2_X1 U1098 ( .A(G1976), .B(G23), .Z(n1011) );
  XOR2_X1 U1099 ( .A(G1971), .B(G22), .Z(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G24), .B(G1986), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(KEYINPUT58), .B(n1014), .Z(n1032) );
  XOR2_X1 U1104 ( .A(KEYINPUT124), .B(G4), .Z(n1016) );
  XNOR2_X1 U1105 ( .A(G1348), .B(KEYINPUT59), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(n1016), .B(n1015), .ZN(n1023) );
  INV_X1 U1107 ( .A(G1341), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(G19), .B(n1017), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(G1981), .B(G6), .ZN(n1019) );
  XNOR2_X1 U1110 ( .A(G1956), .B(G20), .ZN(n1018) );
  NOR2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1112 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(KEYINPUT60), .B(n1024), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(n1025), .B(G5), .ZN(n1026) );
  NAND2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(G21), .B(G1966), .ZN(n1028) );
  NOR2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT125), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1126 ( .A(n1042), .B(KEYINPUT62), .ZN(n1043) );
  XNOR2_X1 U1127 ( .A(KEYINPUT126), .B(n1043), .ZN(G150) );
  INV_X1 U1128 ( .A(G150), .ZN(G311) );
endmodule

