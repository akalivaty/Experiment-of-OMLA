

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XNOR2_X1 U323 ( .A(n298), .B(n329), .ZN(n299) );
  XNOR2_X1 U324 ( .A(n396), .B(n395), .ZN(n570) );
  INV_X1 U325 ( .A(KEYINPUT11), .ZN(n308) );
  XNOR2_X1 U326 ( .A(n307), .B(n306), .ZN(n578) );
  XNOR2_X1 U327 ( .A(n305), .B(n304), .ZN(n306) );
  OR2_X1 U328 ( .A1(n570), .A2(n436), .ZN(n437) );
  XNOR2_X1 U329 ( .A(n322), .B(n321), .ZN(n563) );
  XOR2_X1 U330 ( .A(n368), .B(KEYINPUT113), .Z(n291) );
  XNOR2_X1 U331 ( .A(n369), .B(KEYINPUT47), .ZN(n370) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G106GAT), .ZN(n292) );
  INV_X1 U333 ( .A(KEYINPUT124), .ZN(n394) );
  XNOR2_X1 U334 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U335 ( .A(n292), .B(G85GAT), .ZN(n311) );
  XNOR2_X1 U336 ( .A(n394), .B(KEYINPUT54), .ZN(n395) );
  XNOR2_X1 U337 ( .A(n311), .B(n310), .ZN(n314) );
  XNOR2_X1 U338 ( .A(KEYINPUT101), .B(KEYINPUT36), .ZN(n323) );
  XNOR2_X1 U339 ( .A(n320), .B(n350), .ZN(n321) );
  XNOR2_X1 U340 ( .A(n549), .B(n323), .ZN(n586) );
  NOR2_X1 U341 ( .A1(n533), .A2(n532), .ZN(n553) );
  NOR2_X1 U342 ( .A1(n537), .A2(n536), .ZN(n550) );
  XOR2_X1 U343 ( .A(n472), .B(KEYINPUT28), .Z(n537) );
  XNOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n457) );
  XNOR2_X1 U345 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  INV_X1 U346 ( .A(KEYINPUT32), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n311), .B(n293), .ZN(n295) );
  NAND2_X1 U348 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n300) );
  XOR2_X1 U350 ( .A(G120GAT), .B(G71GAT), .Z(n438) );
  XOR2_X1 U351 ( .A(G148GAT), .B(G78GAT), .Z(n426) );
  XOR2_X1 U352 ( .A(n438), .B(n426), .Z(n298) );
  XOR2_X1 U353 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n297) );
  XNOR2_X1 U354 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n329) );
  XNOR2_X1 U356 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U357 ( .A(G176GAT), .B(G64GAT), .Z(n384) );
  XNOR2_X1 U358 ( .A(n301), .B(n384), .ZN(n307) );
  XOR2_X1 U359 ( .A(KEYINPUT73), .B(KEYINPUT31), .Z(n303) );
  XNOR2_X1 U360 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n302) );
  XOR2_X1 U361 ( .A(n303), .B(n302), .Z(n305) );
  XOR2_X1 U362 ( .A(G204GAT), .B(G92GAT), .Z(n304) );
  INV_X1 U363 ( .A(n578), .ZN(n344) );
  NAND2_X1 U364 ( .A1(G232GAT), .A2(G233GAT), .ZN(n309) );
  XOR2_X1 U365 ( .A(G134GAT), .B(KEYINPUT75), .Z(n397) );
  XNOR2_X1 U366 ( .A(n397), .B(KEYINPUT9), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n312), .B(KEYINPUT10), .ZN(n313) );
  XOR2_X1 U368 ( .A(n314), .B(n313), .Z(n322) );
  XNOR2_X1 U369 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n315), .B(G162GAT), .ZN(n425) );
  XOR2_X1 U371 ( .A(G92GAT), .B(G218GAT), .Z(n317) );
  XNOR2_X1 U372 ( .A(G36GAT), .B(G190GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n381) );
  XNOR2_X1 U374 ( .A(n425), .B(n381), .ZN(n320) );
  XOR2_X1 U375 ( .A(G29GAT), .B(G43GAT), .Z(n319) );
  XNOR2_X1 U376 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n350) );
  XNOR2_X1 U378 ( .A(KEYINPUT76), .B(n563), .ZN(n549) );
  XOR2_X1 U379 ( .A(G78GAT), .B(G183GAT), .Z(n325) );
  XNOR2_X1 U380 ( .A(G127GAT), .B(G71GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U382 ( .A(n326), .B(G211GAT), .Z(n328) );
  XOR2_X1 U383 ( .A(G15GAT), .B(G1GAT), .Z(n348) );
  XNOR2_X1 U384 ( .A(G8GAT), .B(n348), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U386 ( .A(G22GAT), .B(G155GAT), .Z(n422) );
  XOR2_X1 U387 ( .A(n329), .B(n422), .Z(n331) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n333), .B(n332), .Z(n341) );
  XOR2_X1 U391 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n335) );
  XNOR2_X1 U392 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n334) );
  XNOR2_X1 U393 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(KEYINPUT15), .Z(n337) );
  XNOR2_X1 U395 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n582) );
  NOR2_X1 U399 ( .A1(n586), .A2(n582), .ZN(n342) );
  XOR2_X1 U400 ( .A(KEYINPUT45), .B(n342), .Z(n343) );
  NOR2_X1 U401 ( .A1(n344), .A2(n343), .ZN(n345) );
  XNOR2_X1 U402 ( .A(KEYINPUT116), .B(n345), .ZN(n364) );
  XOR2_X1 U403 ( .A(G197GAT), .B(G113GAT), .Z(n347) );
  XNOR2_X1 U404 ( .A(G50GAT), .B(G36GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n349) );
  XOR2_X1 U406 ( .A(n349), .B(n348), .Z(n355) );
  XOR2_X1 U407 ( .A(n350), .B(KEYINPUT30), .Z(n352) );
  NAND2_X1 U408 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n390) );
  XNOR2_X1 U411 ( .A(n353), .B(n390), .ZN(n354) );
  XNOR2_X1 U412 ( .A(n355), .B(n354), .ZN(n363) );
  XOR2_X1 U413 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n357) );
  XNOR2_X1 U414 ( .A(G141GAT), .B(G22GAT), .ZN(n356) );
  XNOR2_X1 U415 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U416 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n359) );
  XNOR2_X1 U417 ( .A(KEYINPUT66), .B(KEYINPUT69), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U419 ( .A(n361), .B(n360), .Z(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n574) );
  NAND2_X1 U421 ( .A1(n364), .A2(n574), .ZN(n373) );
  INV_X1 U422 ( .A(n574), .ZN(n538) );
  XNOR2_X1 U423 ( .A(n578), .B(KEYINPUT64), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT41), .ZN(n541) );
  NAND2_X1 U425 ( .A1(n538), .A2(n541), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n366), .B(KEYINPUT46), .ZN(n367) );
  NAND2_X1 U427 ( .A1(n367), .A2(n582), .ZN(n368) );
  NOR2_X1 U428 ( .A1(n563), .A2(n291), .ZN(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT115), .B(KEYINPUT114), .Z(n369) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  NAND2_X1 U431 ( .A1(n373), .A2(n372), .ZN(n375) );
  INV_X1 U432 ( .A(KEYINPUT48), .ZN(n374) );
  XNOR2_X1 U433 ( .A(n375), .B(n374), .ZN(n533) );
  XOR2_X1 U434 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n377) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U437 ( .A(n378), .B(KEYINPUT90), .Z(n383) );
  XOR2_X1 U438 ( .A(G183GAT), .B(KEYINPUT17), .Z(n380) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n439) );
  XNOR2_X1 U441 ( .A(n439), .B(n381), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U443 ( .A(n385), .B(n384), .Z(n392) );
  XNOR2_X1 U444 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n386), .B(KEYINPUT21), .ZN(n387) );
  XOR2_X1 U446 ( .A(n387), .B(KEYINPUT84), .Z(n389) );
  XNOR2_X1 U447 ( .A(G197GAT), .B(G204GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n432) );
  XNOR2_X1 U449 ( .A(n390), .B(n432), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n526) );
  XNOR2_X1 U451 ( .A(n526), .B(KEYINPUT123), .ZN(n393) );
  NOR2_X1 U452 ( .A1(n533), .A2(n393), .ZN(n396) );
  XOR2_X1 U453 ( .A(n397), .B(G85GAT), .Z(n400) );
  XNOR2_X1 U454 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n398), .B(G127GAT), .ZN(n442) );
  XNOR2_X1 U456 ( .A(n442), .B(G162GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n413) );
  XOR2_X1 U458 ( .A(G155GAT), .B(G148GAT), .Z(n402) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(G120GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U461 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n404) );
  XNOR2_X1 U462 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n403) );
  XNOR2_X1 U463 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U464 ( .A(n406), .B(n405), .Z(n411) );
  XOR2_X1 U465 ( .A(KEYINPUT5), .B(G57GAT), .Z(n408) );
  NAND2_X1 U466 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U468 ( .A(G1GAT), .B(n409), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U470 ( .A(n413), .B(n412), .ZN(n418) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n415) );
  XNOR2_X1 U472 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n414) );
  XNOR2_X1 U473 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U474 ( .A(G141GAT), .B(n416), .Z(n431) );
  INV_X1 U475 ( .A(n431), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n571) );
  INV_X1 U477 ( .A(n571), .ZN(n435) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n420) );
  XNOR2_X1 U479 ( .A(KEYINPUT88), .B(KEYINPUT22), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U481 ( .A(n421), .B(G106GAT), .Z(n424) );
  XNOR2_X1 U482 ( .A(n422), .B(G218GAT), .ZN(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n430) );
  XOR2_X1 U484 ( .A(n426), .B(n425), .Z(n428) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U487 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n472) );
  NAND2_X1 U490 ( .A1(n435), .A2(n472), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(KEYINPUT55), .ZN(n455) );
  XOR2_X1 U492 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U493 ( .A(G99GAT), .B(G134GAT), .ZN(n440) );
  XNOR2_X1 U494 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U495 ( .A(n442), .B(KEYINPUT20), .Z(n444) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U497 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U498 ( .A(n446), .B(n445), .Z(n454) );
  XOR2_X1 U499 ( .A(KEYINPUT81), .B(KEYINPUT82), .Z(n448) );
  XNOR2_X1 U500 ( .A(G43GAT), .B(G190GAT), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT83), .B(G176GAT), .Z(n450) );
  XNOR2_X1 U503 ( .A(G169GAT), .B(G15GAT), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U506 ( .A(n454), .B(n453), .ZN(n534) );
  NAND2_X1 U507 ( .A1(n455), .A2(n534), .ZN(n568) );
  INV_X1 U508 ( .A(n568), .ZN(n456) );
  NAND2_X1 U509 ( .A1(n456), .A2(n549), .ZN(n458) );
  INV_X1 U510 ( .A(n541), .ZN(n555) );
  NOR2_X1 U511 ( .A1(n555), .A2(n568), .ZN(n461) );
  XNOR2_X1 U512 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n459), .B(G176GAT), .ZN(n460) );
  XNOR2_X1 U514 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U515 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n482) );
  NAND2_X1 U516 ( .A1(n538), .A2(n578), .ZN(n496) );
  NOR2_X1 U517 ( .A1(n549), .A2(n582), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT16), .ZN(n480) );
  NAND2_X1 U519 ( .A1(n534), .A2(n526), .ZN(n463) );
  NAND2_X1 U520 ( .A1(n472), .A2(n463), .ZN(n464) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n464), .Z(n469) );
  XOR2_X1 U522 ( .A(n526), .B(KEYINPUT93), .Z(n465) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n465), .ZN(n473) );
  NOR2_X1 U524 ( .A1(n534), .A2(n472), .ZN(n466) );
  XOR2_X1 U525 ( .A(KEYINPUT26), .B(n466), .Z(n467) );
  XNOR2_X1 U526 ( .A(KEYINPUT95), .B(n467), .ZN(n572) );
  NAND2_X1 U527 ( .A1(n473), .A2(n572), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U529 ( .A(KEYINPUT96), .B(n470), .Z(n471) );
  NOR2_X1 U530 ( .A1(n571), .A2(n471), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n571), .A2(n473), .ZN(n532) );
  NOR2_X1 U532 ( .A1(n537), .A2(n532), .ZN(n475) );
  INV_X1 U533 ( .A(n534), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n476) );
  XOR2_X1 U535 ( .A(KEYINPUT94), .B(n476), .Z(n477) );
  NOR2_X1 U536 ( .A1(n478), .A2(n477), .ZN(n492) );
  INV_X1 U537 ( .A(n492), .ZN(n479) );
  NAND2_X1 U538 ( .A1(n480), .A2(n479), .ZN(n509) );
  NOR2_X1 U539 ( .A1(n496), .A2(n509), .ZN(n487) );
  NAND2_X1 U540 ( .A1(n487), .A2(n571), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n483), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n487), .A2(n526), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U546 ( .A1(n487), .A2(n534), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n489) );
  NAND2_X1 U549 ( .A1(n487), .A2(n537), .ZN(n488) );
  XNOR2_X1 U550 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  XNOR2_X1 U553 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n491), .B(KEYINPUT37), .ZN(n495) );
  NOR2_X1 U555 ( .A1(n586), .A2(n492), .ZN(n493) );
  NAND2_X1 U556 ( .A1(n582), .A2(n493), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n522) );
  NOR2_X1 U558 ( .A1(n496), .A2(n522), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT38), .ZN(n507) );
  NAND2_X1 U560 ( .A1(n507), .A2(n571), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U562 ( .A(n500), .B(KEYINPUT104), .Z(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT100), .B(KEYINPUT105), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  NAND2_X1 U565 ( .A1(n507), .A2(n526), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n503), .B(KEYINPUT106), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(n504), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n507), .A2(n534), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  NAND2_X1 U571 ( .A1(n507), .A2(n537), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT107), .Z(n512) );
  NAND2_X1 U574 ( .A1(n541), .A2(n574), .ZN(n523) );
  NOR2_X1 U575 ( .A1(n523), .A2(n509), .ZN(n510) );
  XNOR2_X1 U576 ( .A(KEYINPUT108), .B(n510), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n519), .A2(n571), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n512), .B(n511), .ZN(n514) );
  XOR2_X1 U579 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U581 ( .A1(n519), .A2(n526), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n517) );
  NAND2_X1 U584 ( .A1(n534), .A2(n519), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U586 ( .A(G71GAT), .B(n518), .ZN(G1334GAT) );
  XOR2_X1 U587 ( .A(G78GAT), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U588 ( .A1(n537), .A2(n519), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(G1335GAT) );
  NOR2_X1 U590 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT112), .ZN(n529) );
  NAND2_X1 U592 ( .A1(n571), .A2(n529), .ZN(n525) );
  XNOR2_X1 U593 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n526), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n529), .A2(n534), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n529), .A2(n537), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U600 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n553), .ZN(n535) );
  XOR2_X1 U602 ( .A(KEYINPUT117), .B(n535), .Z(n536) );
  NAND2_X1 U603 ( .A1(n538), .A2(n550), .ZN(n539) );
  XNOR2_X1 U604 ( .A(KEYINPUT118), .B(n539), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .Z(n543) );
  NAND2_X1 U607 ( .A1(n550), .A2(n541), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  INV_X1 U609 ( .A(n582), .ZN(n544) );
  NAND2_X1 U610 ( .A1(n544), .A2(n550), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n546) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(KEYINPUT120), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U615 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NAND2_X1 U618 ( .A1(n553), .A2(n572), .ZN(n561) );
  NOR2_X1 U619 ( .A1(n574), .A2(n561), .ZN(n554) );
  XOR2_X1 U620 ( .A(G141GAT), .B(n554), .Z(G1344GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n561), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U625 ( .A1(n582), .A2(n561), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1346GAT) );
  INV_X1 U628 ( .A(n561), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT122), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G162GAT), .B(n565), .ZN(G1347GAT) );
  NOR2_X1 U632 ( .A1(n574), .A2(n568), .ZN(n567) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(KEYINPUT125), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  NOR2_X1 U635 ( .A1(n582), .A2(n568), .ZN(n569) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n569), .Z(G1350GAT) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n585) );
  NOR2_X1 U639 ( .A1(n574), .A2(n585), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n585), .ZN(n580) );
  XNOR2_X1 U644 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

