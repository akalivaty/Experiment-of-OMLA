//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT2), .B(G113), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G116), .B(G119), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n191), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT30), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT11), .A2(G134), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G131), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G137), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n200), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n203), .A2(G134), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n206), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(G137), .B1(new_n202), .B2(new_n204), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n215), .A2(KEYINPUT65), .A3(KEYINPUT11), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n199), .B(new_n208), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n196), .A2(new_n201), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n200), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  INV_X1    g035(.A(G143), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n225), .A3(G128), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n221), .B(new_n223), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n219), .A2(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n217), .A2(KEYINPUT67), .A3(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT67), .B1(new_n217), .B2(new_n230), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n221), .A2(new_n223), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT0), .A3(G128), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT0), .B(G128), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT65), .B1(new_n215), .B2(KEYINPUT11), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(G134), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n209), .B(new_n213), .C1(new_n240), .C2(G137), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n198), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n205), .A2(new_n206), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n200), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  AOI211_X1 g059(.A(new_n198), .B(new_n207), .C1(new_n239), .C2(new_n241), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n238), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n195), .B1(new_n233), .B2(new_n247), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n199), .B(new_n244), .C1(new_n214), .C2(new_n216), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n237), .B1(new_n250), .B2(new_n217), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n219), .A2(new_n229), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n251), .A2(KEYINPUT30), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n194), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g069(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n256));
  NOR2_X1   g070(.A1(G237), .A2(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n256), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n194), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n264), .B1(new_n246), .B2(new_n252), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n217), .A2(KEYINPUT67), .A3(new_n230), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n247), .A2(new_n263), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n255), .A2(new_n262), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n267), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n266), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT30), .B1(new_n272), .B2(new_n251), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n247), .B(new_n195), .C1(new_n246), .C2(new_n252), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n275), .B2(new_n194), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(KEYINPUT31), .A3(new_n262), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n194), .B1(new_n251), .B2(new_n253), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n267), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT28), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT69), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n251), .A2(new_n253), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n285), .B2(new_n263), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n261), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n188), .B1(new_n278), .B2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT70), .B1(new_n290), .B2(KEYINPUT32), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT32), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n270), .A2(new_n277), .B1(new_n288), .B2(new_n261), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n188), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n194), .B1(new_n272), .B2(new_n251), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n267), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n286), .B1(new_n297), .B2(KEYINPUT28), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n262), .A2(KEYINPUT29), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n255), .A2(new_n267), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n301), .B2(new_n261), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n286), .A2(new_n261), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n284), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT69), .B1(new_n280), .B2(KEYINPUT28), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT28), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n282), .B(new_n307), .C1(new_n279), .C2(new_n267), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT71), .B1(new_n309), .B2(new_n303), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n300), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n290), .A2(KEYINPUT32), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n291), .A2(new_n295), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(G210), .B1(G237), .B2(G902), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n315), .B(KEYINPUT84), .Z(new_n316));
  MUX2_X1   g130(.A(new_n229), .B(new_n237), .S(G125), .Z(new_n317));
  INV_X1    g131(.A(G224), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G953), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n317), .B(new_n319), .Z(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G122), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n321), .B(KEYINPUT82), .Z(new_n322));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n323));
  INV_X1    g137(.A(G107), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(G104), .ZN(new_n325));
  INV_X1    g139(.A(G104), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT77), .A3(G107), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n324), .A2(KEYINPUT3), .A3(G104), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT3), .B1(new_n324), .B2(G104), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n325), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G101), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n194), .B1(new_n331), .B2(KEYINPUT4), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(new_n333), .A3(G101), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n326), .B2(G107), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n324), .A2(KEYINPUT3), .A3(G104), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G101), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n338), .A2(new_n339), .A3(new_n325), .A4(new_n327), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n334), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n333), .B1(new_n330), .B2(G101), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT79), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(new_n342), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n340), .A2(KEYINPUT4), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .A4(new_n334), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n332), .B1(new_n343), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n191), .A2(KEYINPUT5), .ZN(new_n349));
  INV_X1    g163(.A(G116), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n350), .A2(KEYINPUT5), .A3(G119), .ZN(new_n351));
  INV_X1    g165(.A(G113), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n326), .A2(G107), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n324), .A2(G104), .ZN(new_n356));
  OAI21_X1  g170(.A(G101), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n354), .A2(new_n340), .A3(new_n193), .A4(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n322), .B1(new_n348), .B2(new_n360), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n348), .A2(new_n322), .A3(new_n360), .ZN(new_n362));
  NAND2_X1  g176(.A1(KEYINPUT83), .A2(KEYINPUT6), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n363), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n322), .B(new_n365), .C1(new_n348), .C2(new_n360), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n320), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT7), .B1(new_n318), .B2(G953), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n317), .B(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n322), .B(KEYINPUT8), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n354), .A2(new_n193), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n340), .A2(new_n357), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n358), .B2(new_n373), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n343), .A2(new_n347), .ZN(new_n376));
  INV_X1    g190(.A(new_n332), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n322), .ZN(new_n379));
  INV_X1    g193(.A(new_n360), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G902), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n316), .B1(new_n367), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n316), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n375), .B2(new_n381), .ZN(new_n387));
  INV_X1    g201(.A(new_n366), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n381), .A2(new_n365), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n388), .B1(new_n389), .B2(new_n361), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n386), .B(new_n387), .C1(new_n390), .C2(new_n320), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT20), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n394), .A2(new_n395), .A3(G125), .ZN(new_n396));
  XNOR2_X1  g210(.A(G125), .B(G140), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G146), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n220), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n222), .A2(KEYINPUT85), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(G214), .A3(new_n257), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT85), .B(G143), .ZN(new_n404));
  INV_X1    g218(.A(G237), .ZN(new_n405));
  INV_X1    g219(.A(G953), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n405), .A2(new_n406), .A3(G214), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n403), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n200), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G143), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n412), .A2(new_n402), .B1(new_n257), .B2(G214), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n406), .A3(G214), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n411), .A2(G143), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(G131), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  OAI221_X1 g231(.A(new_n401), .B1(new_n408), .B2(new_n410), .C1(new_n409), .C2(new_n417), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n403), .B(new_n200), .C1(new_n404), .C2(new_n407), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(KEYINPUT86), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n412), .A2(new_n402), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n414), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n200), .A4(new_n403), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(KEYINPUT87), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT16), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n395), .A3(G125), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT74), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n428), .B(G146), .C1(new_n398), .C2(new_n426), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n397), .A2(KEYINPUT19), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT19), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n430), .B1(new_n398), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n220), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n425), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(KEYINPUT87), .B1(new_n420), .B2(new_n424), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n418), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G113), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(new_n326), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n428), .B1(new_n398), .B2(new_n426), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n220), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n200), .B1(new_n422), .B2(new_n403), .ZN(new_n443));
  AOI21_X1  g257(.A(KEYINPUT88), .B1(new_n443), .B2(KEYINPUT17), .ZN(new_n444));
  AND4_X1   g258(.A1(KEYINPUT88), .A2(new_n408), .A3(KEYINPUT17), .A4(G131), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n442), .B(new_n429), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT17), .B1(new_n420), .B2(new_n424), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n438), .B(new_n418), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(G475), .A2(G902), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT89), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n393), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AOI211_X1 g267(.A(KEYINPUT20), .B(new_n451), .C1(new_n440), .C2(new_n448), .ZN(new_n454));
  INV_X1    g268(.A(G475), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n418), .B1(new_n446), .B2(new_n447), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n439), .ZN(new_n457));
  AOI21_X1  g271(.A(G902), .B1(new_n457), .B2(new_n448), .ZN(new_n458));
  OAI22_X1  g272(.A1(new_n453), .A2(new_n454), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT92), .ZN(new_n460));
  INV_X1    g274(.A(G122), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G116), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n350), .A2(G122), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G107), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(new_n324), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n227), .A2(G143), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n222), .A2(G128), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n240), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT13), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n473), .B1(new_n227), .B2(G143), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT90), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n222), .A2(G128), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT90), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n227), .A2(G143), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n476), .B2(new_n473), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n201), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT91), .B1(new_n472), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n465), .A2(new_n466), .B1(new_n470), .B2(new_n240), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT91), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n481), .B1(new_n478), .B2(new_n475), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n486), .C1(new_n201), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n350), .A2(KEYINPUT14), .A3(G122), .ZN(new_n489));
  OAI211_X1 g303(.A(G107), .B(new_n489), .C1(new_n464), .C2(KEYINPUT14), .ZN(new_n490));
  INV_X1    g304(.A(new_n471), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n470), .A2(new_n240), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n466), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n484), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT9), .B(G234), .ZN(new_n495));
  INV_X1    g309(.A(G217), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(G953), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n484), .A2(new_n488), .A3(new_n493), .A4(new_n497), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n460), .B(G902), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G478), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(G902), .B1(new_n499), .B2(new_n500), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(KEYINPUT92), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n503), .B1(new_n507), .B2(new_n501), .ZN(new_n508));
  INV_X1    g322(.A(G952), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G953), .ZN(new_n510));
  INV_X1    g324(.A(G234), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n405), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n383), .B(new_n406), .C1(G234), .C2(G237), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n508), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n459), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G214), .B1(G237), .B2(G902), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n392), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G137), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n406), .A2(G221), .A3(G234), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT75), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n227), .A2(G119), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n227), .A2(G119), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n528), .B1(KEYINPUT72), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(KEYINPUT72), .B(KEYINPUT23), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n527), .C1(new_n534), .C2(new_n528), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n531), .B1(new_n535), .B2(G110), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n537), .B1(new_n442), .B2(new_n429), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n529), .A2(new_n530), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n535), .B2(G110), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n429), .A2(new_n540), .A3(new_n400), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n526), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n442), .A2(new_n429), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n536), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n541), .A3(new_n524), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT25), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n383), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n496), .B1(G234), .B2(new_n383), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n546), .A3(new_n383), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(KEYINPUT25), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n550), .A2(G902), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n543), .A2(new_n546), .A3(new_n555), .ZN(new_n556));
  OR2_X1    g370(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(G221), .B1(new_n495), .B2(G902), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G469), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n383), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n340), .A2(new_n228), .A3(new_n226), .A4(new_n357), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT10), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n331), .A2(KEYINPUT4), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n237), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n376), .B2(new_n568), .ZN(new_n569));
  AOI211_X1 g383(.A(new_n243), .B(new_n198), .C1(new_n239), .C2(new_n241), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n217), .B1(new_n570), .B2(new_n200), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT80), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT80), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n250), .A2(new_n573), .A3(new_n217), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n576));
  INV_X1    g390(.A(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n372), .A2(new_n229), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n564), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n576), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(KEYINPUT12), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G140), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n406), .A2(G227), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n585), .B(new_n586), .Z(new_n587));
  AND2_X1   g401(.A1(new_n572), .A2(new_n574), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(new_n569), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n569), .A2(new_n577), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n584), .A2(new_n587), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n563), .B1(new_n591), .B2(G469), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n589), .A2(new_n583), .ZN(new_n593));
  INV_X1    g407(.A(new_n587), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n590), .B2(new_n575), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n562), .B(new_n383), .C1(new_n593), .C2(new_n595), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n559), .B(new_n561), .C1(new_n592), .C2(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n521), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n314), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(KEYINPUT93), .B(G101), .Z(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G3));
  OAI21_X1  g415(.A(G472), .B1(new_n294), .B2(G902), .ZN(new_n602));
  NOR3_X1   g416(.A1(new_n306), .A2(new_n308), .A3(new_n286), .ZN(new_n603));
  AOI21_X1  g417(.A(KEYINPUT31), .B1(new_n276), .B2(new_n262), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n263), .B1(new_n273), .B2(new_n274), .ZN(new_n605));
  NOR4_X1   g419(.A1(new_n605), .A2(new_n271), .A3(new_n269), .A4(new_n261), .ZN(new_n606));
  OAI22_X1  g420(.A1(new_n603), .A2(new_n262), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n187), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n602), .A2(new_n597), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT94), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n385), .A2(new_n391), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n367), .A2(new_n384), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(KEYINPUT94), .A3(new_n386), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n612), .A2(new_n614), .A3(new_n520), .ZN(new_n615));
  NAND2_X1  g429(.A1(G478), .A2(G902), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n499), .A2(new_n500), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n383), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n618), .B2(G478), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n494), .B2(KEYINPUT95), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n617), .B(new_n621), .Z(new_n622));
  AOI21_X1  g436(.A(new_n619), .B1(new_n622), .B2(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n459), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n615), .A2(new_n516), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n610), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  AND2_X1   g442(.A1(new_n614), .A2(new_n520), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n420), .A2(new_n424), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n632), .A2(new_n429), .A3(new_n425), .A4(new_n433), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n438), .B1(new_n633), .B2(new_n418), .ZN(new_n634));
  INV_X1    g448(.A(new_n448), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n452), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT20), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n449), .A2(new_n393), .A3(new_n452), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n457), .A2(new_n448), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n455), .B1(new_n640), .B2(new_n383), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n505), .A2(new_n508), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n639), .A2(new_n643), .A3(new_n644), .A4(new_n517), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n629), .A2(new_n645), .A3(new_n612), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n610), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n647), .B(KEYINPUT97), .Z(new_n648));
  XNOR2_X1  g462(.A(KEYINPUT35), .B(G107), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT36), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n525), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT98), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n538), .A2(new_n542), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(new_n555), .B1(new_n549), .B2(new_n553), .ZN(new_n656));
  AOI211_X1 g470(.A(new_n561), .B(new_n656), .C1(new_n592), .C2(new_n596), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n602), .A2(new_n521), .A3(new_n657), .A4(new_n608), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  NAND2_X1  g474(.A1(new_n592), .A2(new_n596), .ZN(new_n661));
  INV_X1    g475(.A(new_n656), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n560), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n513), .B1(new_n514), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n643), .A2(new_n639), .A3(new_n644), .A4(new_n666), .ZN(new_n667));
  NOR3_X1   g481(.A1(new_n663), .A2(new_n615), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n314), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT99), .B(G128), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G30));
  XOR2_X1   g485(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n392), .B(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n618), .A2(new_n460), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n506), .A2(KEYINPUT92), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n504), .B1(new_n677), .B2(new_n503), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n661), .A2(new_n560), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n665), .B(new_n681), .Z(new_n682));
  NOR2_X1   g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n520), .B(new_n679), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n673), .B(new_n685), .C1(new_n684), .C2(new_n683), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n297), .A2(new_n261), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n268), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n383), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n290), .A2(KEYINPUT32), .B1(G472), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n291), .A3(new_n295), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n686), .A2(new_n656), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT102), .B(G143), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G45));
  NAND3_X1  g508(.A1(new_n459), .A2(new_n623), .A3(new_n666), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n663), .A2(new_n615), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n314), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G146), .ZN(G48));
  INV_X1    g512(.A(new_n559), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n590), .A2(new_n575), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n700), .A2(new_n587), .B1(new_n589), .B2(new_n583), .ZN(new_n701));
  OAI21_X1  g515(.A(G469), .B1(new_n701), .B2(G902), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n560), .A3(new_n596), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n314), .A2(new_n699), .A3(new_n625), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND4_X1  g521(.A1(new_n314), .A2(new_n699), .A3(new_n646), .A4(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NAND2_X1  g523(.A1(new_n519), .A2(new_n662), .ZN(new_n710));
  NOR3_X1   g524(.A1(new_n615), .A2(new_n703), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n314), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  XNOR2_X1  g527(.A(KEYINPUT103), .B(G472), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n607), .B2(new_n383), .ZN(new_n716));
  OR2_X1    g530(.A1(new_n298), .A2(new_n262), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n188), .B1(new_n278), .B2(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n559), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT104), .B1(new_n674), .B2(new_n678), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n459), .A2(new_n721), .A3(new_n644), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n720), .A2(new_n722), .A3(new_n517), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n615), .A2(new_n723), .A3(new_n703), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR3_X1   g540(.A1(new_n716), .A2(new_n656), .A3(new_n718), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n615), .A2(new_n695), .A3(new_n703), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND3_X1  g544(.A1(new_n385), .A2(new_n391), .A3(new_n520), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n680), .A2(new_n695), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n314), .A2(new_n699), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT42), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT105), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n294), .A2(new_n293), .A3(new_n188), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT32), .B1(new_n607), .B2(new_n187), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n293), .B1(new_n294), .B2(new_n188), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n313), .A2(new_n740), .A3(KEYINPUT105), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n312), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n732), .A2(KEYINPUT42), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n699), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G131), .ZN(G33));
  NOR3_X1   g560(.A1(new_n680), .A2(new_n667), .A3(new_n731), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n314), .A2(new_n699), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  AOI21_X1  g563(.A(new_n656), .B1(new_n602), .B2(new_n608), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n674), .A2(new_n623), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT43), .Z(new_n753));
  AND2_X1   g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT107), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT44), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n584), .A2(new_n587), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n589), .A2(new_n590), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n562), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(new_n764), .B2(new_n763), .ZN(new_n766));
  INV_X1    g580(.A(new_n563), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(KEYINPUT46), .A3(new_n767), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n596), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n560), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n682), .ZN(new_n774));
  INV_X1    g588(.A(new_n731), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n760), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n759), .A2(new_n777), .ZN(new_n778));
  XOR2_X1   g592(.A(KEYINPUT108), .B(G137), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT109), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n778), .B(new_n780), .ZN(G39));
  XOR2_X1   g595(.A(new_n773), .B(KEYINPUT47), .Z(new_n782));
  NOR4_X1   g596(.A1(new_n314), .A2(new_n699), .A3(new_n695), .A4(new_n731), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  INV_X1    g599(.A(new_n691), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n702), .A2(new_n596), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n787), .A2(KEYINPUT49), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n699), .A2(new_n560), .A3(new_n520), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n788), .A2(new_n789), .A3(new_n752), .A4(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n786), .A2(new_n791), .A3(new_n673), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT114), .ZN(new_n793));
  AOI22_X1  g607(.A1(new_n314), .A2(new_n711), .B1(new_n719), .B2(new_n724), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n794), .A2(new_n705), .A3(new_n708), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n680), .A2(new_n731), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n643), .A2(new_n639), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n797), .A2(new_n644), .A3(new_n656), .A4(new_n665), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n314), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n727), .A2(new_n732), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n748), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n745), .A3(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n624), .B(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n392), .A2(new_n520), .A3(new_n517), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n610), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n599), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n459), .A2(new_n678), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n520), .A2(new_n392), .A3(new_n811), .A4(new_n517), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n608), .A3(new_n602), .A4(new_n597), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT112), .B1(new_n813), .B2(new_n658), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(new_n658), .A3(KEYINPUT112), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n599), .A2(new_n807), .A3(KEYINPUT111), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n810), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n802), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n314), .A2(new_n668), .B1(new_n727), .B2(new_n728), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n720), .A2(new_n722), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n615), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n680), .A2(new_n665), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n691), .A2(new_n656), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n825), .A3(new_n697), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n821), .A2(new_n825), .A3(new_n828), .A4(new_n697), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n820), .A2(KEYINPUT53), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT53), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n827), .A2(KEYINPUT113), .A3(new_n829), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT113), .B1(new_n827), .B2(new_n829), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n820), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n832), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n793), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n820), .B(KEYINPUT53), .C1(new_n834), .C2(new_n835), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n748), .A2(new_n799), .A3(new_n800), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n841), .B1(new_n735), .B2(new_n744), .ZN(new_n842));
  INV_X1    g656(.A(new_n818), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT111), .B1(new_n599), .B2(new_n807), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n842), .A2(new_n845), .A3(new_n817), .A4(new_n795), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n827), .A2(new_n829), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n833), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g662(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n840), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n836), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n831), .B1(new_n851), .B2(KEYINPUT53), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n742), .A2(new_n699), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n753), .A2(new_n513), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n703), .A2(new_n731), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT48), .Z(new_n859));
  NAND2_X1  g673(.A1(new_n855), .A2(new_n719), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n615), .A2(new_n703), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n786), .A2(new_n699), .A3(new_n513), .A4(new_n856), .ZN(new_n863));
  OAI221_X1 g677(.A(new_n510), .B1(new_n860), .B2(new_n862), .C1(new_n863), .C2(new_n624), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n855), .A2(new_n719), .A3(new_n775), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT117), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n787), .A2(new_n560), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n867), .B(new_n868), .C1(new_n782), .C2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n520), .B1(KEYINPUT118), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n673), .A2(new_n704), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n459), .A2(new_n623), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n874), .A2(new_n876), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n860), .A2(new_n875), .A3(new_n873), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n857), .A2(new_n727), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(KEYINPUT116), .B1(new_n870), .B2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT51), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n865), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n883), .B2(new_n882), .ZN(new_n885));
  AND4_X1   g699(.A1(new_n839), .A2(new_n850), .A3(new_n853), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(G952), .A2(G953), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT119), .Z(new_n888));
  OAI21_X1  g702(.A(new_n792), .B1(new_n886), .B2(new_n888), .ZN(G75));
  NAND2_X1  g703(.A1(new_n509), .A2(G953), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT121), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n813), .A2(KEYINPUT112), .A3(new_n658), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n814), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n843), .A2(new_n893), .A3(new_n844), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n894), .A2(KEYINPUT53), .A3(new_n795), .A4(new_n842), .ZN(new_n895));
  INV_X1    g709(.A(new_n834), .ZN(new_n896));
  INV_X1    g710(.A(new_n835), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT53), .B1(new_n820), .B2(new_n830), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n383), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT56), .B1(new_n901), .B2(new_n316), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n390), .B(new_n320), .Z(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT55), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n891), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n840), .A2(new_n848), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n906), .A2(new_n907), .A3(G902), .A4(new_n316), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n909), .A3(new_n904), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n901), .A2(new_n316), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(KEYINPUT120), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n905), .A2(new_n912), .ZN(G51));
  AOI211_X1 g727(.A(new_n383), .B(new_n766), .C1(new_n840), .C2(new_n848), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n563), .B(KEYINPUT57), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n840), .A2(new_n848), .A3(new_n849), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n849), .B1(new_n840), .B2(new_n848), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n701), .B(KEYINPUT122), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n891), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT123), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  INV_X1    g737(.A(new_n919), .ZN(new_n924));
  INV_X1    g738(.A(new_n849), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n898), .B2(new_n899), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n850), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n927), .B2(new_n915), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n923), .B(new_n891), .C1(new_n928), .C2(new_n914), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n922), .A2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n449), .ZN(new_n932));
  INV_X1    g746(.A(new_n449), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .A4(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n921), .B1(new_n932), .B2(new_n934), .ZN(G60));
  INV_X1    g749(.A(new_n927), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n616), .B(KEYINPUT59), .Z(new_n937));
  OR2_X1    g751(.A1(new_n622), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n891), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n937), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n853), .A2(new_n850), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT114), .B1(new_n852), .B2(KEYINPUT54), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n939), .B1(new_n943), .B2(new_n622), .ZN(G63));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  XNOR2_X1  g759(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n900), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n655), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n891), .B1(new_n949), .B2(new_n547), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n949), .A2(new_n547), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT61), .A3(new_n891), .A4(new_n950), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(new_n515), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n406), .B1(new_n957), .B2(G224), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n894), .A2(new_n795), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n958), .B1(new_n959), .B2(new_n406), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n390), .B1(G898), .B2(new_n406), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n960), .B(new_n961), .Z(G69));
  AND2_X1   g776(.A1(new_n821), .A2(new_n697), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n692), .A2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(KEYINPUT62), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n804), .B1(new_n459), .B2(new_n678), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n680), .A2(new_n682), .A3(new_n731), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n314), .A2(new_n699), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n965), .A2(new_n784), .A3(new_n966), .A4(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n778), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n406), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n275), .B(new_n432), .Z(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT125), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n973), .B1(G900), .B2(G953), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n774), .A2(new_n854), .A3(new_n823), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n748), .A2(new_n784), .A3(new_n963), .A4(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n778), .A3(new_n745), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n976), .B1(new_n979), .B2(G953), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n975), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n406), .B1(G227), .B2(G900), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(new_n980), .B2(KEYINPUT126), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n975), .B(new_n980), .C1(KEYINPUT126), .C2(new_n982), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  XNOR2_X1  g800(.A(new_n276), .B(KEYINPUT127), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n970), .A2(new_n971), .A3(new_n959), .ZN(new_n988));
  NAND2_X1  g802(.A1(G472), .A2(G902), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n989), .B(KEYINPUT63), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n262), .B(new_n987), .C1(new_n988), .C2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n979), .B2(new_n959), .ZN(new_n993));
  INV_X1    g807(.A(new_n987), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n993), .A2(new_n261), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n992), .A2(new_n891), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n301), .A2(new_n261), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n991), .B(new_n837), .C1(new_n268), .C2(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(G57));
endmodule


