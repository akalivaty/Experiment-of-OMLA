

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784;

  NOR2_X1 U378 ( .A1(n451), .A2(n618), .ZN(n667) );
  XNOR2_X1 U379 ( .A(n566), .B(n457), .ZN(n766) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n508) );
  BUF_X1 U381 ( .A(n739), .Z(n746) );
  NAND2_X1 U382 ( .A1(n413), .A2(n411), .ZN(n378) );
  INV_X1 U383 ( .A(G953), .ZN(n758) );
  XNOR2_X2 U384 ( .A(n384), .B(n375), .ZN(n694) );
  XNOR2_X2 U385 ( .A(KEYINPUT3), .B(KEYINPUT88), .ZN(n374) );
  NAND2_X1 U386 ( .A1(n694), .A2(n693), .ZN(n419) );
  XNOR2_X2 U387 ( .A(n477), .B(n476), .ZN(n709) );
  AND2_X2 U388 ( .A1(n438), .A2(n502), .ZN(n771) );
  AND2_X1 U389 ( .A1(n697), .A2(n360), .ZN(n693) );
  INV_X2 U390 ( .A(G143), .ZN(n394) );
  INV_X4 U391 ( .A(KEYINPUT4), .ZN(n452) );
  AND2_X2 U392 ( .A1(n495), .A2(n492), .ZN(n739) );
  NAND2_X1 U393 ( .A1(n465), .A2(n371), .ZN(n495) );
  OR2_X1 U394 ( .A1(n750), .A2(n493), .ZN(n492) );
  NOR2_X1 U395 ( .A1(n422), .A2(n420), .ZN(n461) );
  NOR2_X1 U396 ( .A1(n783), .A2(KEYINPUT46), .ZN(n426) );
  XNOR2_X1 U397 ( .A(n597), .B(n598), .ZN(n780) );
  NAND2_X1 U398 ( .A1(n403), .A2(n401), .ZN(n407) );
  XNOR2_X1 U399 ( .A(n382), .B(n381), .ZN(n678) );
  XNOR2_X1 U400 ( .A(n538), .B(n449), .ZN(n697) );
  XNOR2_X1 U401 ( .A(n523), .B(n468), .ZN(n592) );
  XNOR2_X1 U402 ( .A(n560), .B(n480), .ZN(n736) );
  OR2_X1 U403 ( .A1(n661), .A2(G902), .ZN(n443) );
  XNOR2_X1 U404 ( .A(n473), .B(n472), .ZN(n755) );
  XNOR2_X1 U405 ( .A(G110), .B(G104), .ZN(n473) );
  NOR2_X2 U406 ( .A1(n635), .A2(n636), .ZN(n637) );
  XNOR2_X2 U407 ( .A(n768), .B(G146), .ZN(n560) );
  XNOR2_X2 U408 ( .A(n548), .B(n547), .ZN(n768) );
  NOR2_X1 U409 ( .A1(n678), .A2(n715), .ZN(n576) );
  NAND2_X1 U410 ( .A1(n421), .A2(n688), .ZN(n420) );
  NAND2_X1 U411 ( .A1(n424), .A2(n423), .ZN(n422) );
  OR2_X1 U412 ( .A1(n779), .A2(KEYINPUT83), .ZN(n643) );
  AND2_X1 U413 ( .A1(n779), .A2(n389), .ZN(n388) );
  INV_X1 U414 ( .A(KEYINPUT38), .ZN(n474) );
  OR2_X1 U415 ( .A1(G237), .A2(G902), .ZN(n574) );
  AND2_X1 U416 ( .A1(n447), .A2(n446), .ZN(n445) );
  NOR2_X1 U417 ( .A1(n361), .A2(n355), .ZN(n446) );
  NOR2_X1 U418 ( .A1(n436), .A2(n434), .ZN(n431) );
  XNOR2_X1 U419 ( .A(n637), .B(KEYINPUT33), .ZN(n719) );
  XNOR2_X1 U420 ( .A(n703), .B(KEYINPUT106), .ZN(n379) );
  XNOR2_X1 U421 ( .A(n614), .B(n613), .ZN(n619) );
  XNOR2_X1 U422 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n613) );
  NAND2_X1 U423 ( .A1(n445), .A2(n444), .ZN(n614) );
  OR2_X1 U424 ( .A1(n603), .A2(KEYINPUT19), .ZN(n444) );
  INV_X1 U425 ( .A(KEYINPUT1), .ZN(n375) );
  XNOR2_X1 U426 ( .A(n537), .B(KEYINPUT25), .ZN(n449) );
  NAND2_X1 U427 ( .A1(n426), .A2(n425), .ZN(n424) );
  NAND2_X1 U428 ( .A1(n377), .A2(n782), .ZN(n633) );
  INV_X1 U429 ( .A(n690), .ZN(n604) );
  XNOR2_X1 U430 ( .A(n549), .B(n463), .ZN(n462) );
  INV_X1 U431 ( .A(KEYINPUT94), .ZN(n463) );
  XNOR2_X1 U432 ( .A(G137), .B(KEYINPUT71), .ZN(n549) );
  XNOR2_X1 U433 ( .A(G137), .B(G140), .ZN(n561) );
  INV_X1 U434 ( .A(KEYINPUT74), .ZN(n460) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n571) );
  XNOR2_X1 U436 ( .A(G116), .B(G113), .ZN(n372) );
  XNOR2_X1 U437 ( .A(n374), .B(n552), .ZN(n373) );
  INV_X1 U438 ( .A(G119), .ZN(n552) );
  XNOR2_X1 U439 ( .A(n484), .B(n483), .ZN(n438) );
  INV_X1 U440 ( .A(KEYINPUT48), .ZN(n483) );
  AND2_X1 U441 ( .A1(n467), .A2(n466), .ZN(n479) );
  INV_X1 U442 ( .A(KEYINPUT89), .ZN(n572) );
  XNOR2_X1 U443 ( .A(n524), .B(n469), .ZN(n468) );
  NOR2_X1 U444 ( .A1(G902), .A2(n744), .ZN(n523) );
  INV_X1 U445 ( .A(G478), .ZN(n469) );
  INV_X1 U446 ( .A(G107), .ZN(n472) );
  XNOR2_X1 U447 ( .A(n518), .B(n471), .ZN(n470) );
  INV_X1 U448 ( .A(KEYINPUT100), .ZN(n471) );
  XNOR2_X1 U449 ( .A(G116), .B(G122), .ZN(n518) );
  INV_X1 U450 ( .A(G134), .ZN(n514) );
  XNOR2_X1 U451 ( .A(n511), .B(n512), .ZN(n661) );
  XNOR2_X1 U452 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U453 ( .A(n547), .B(n440), .ZN(n510) );
  BUF_X1 U454 ( .A(n648), .Z(n750) );
  INV_X1 U455 ( .A(KEYINPUT41), .ZN(n476) );
  NAND2_X1 U456 ( .A1(n615), .A2(n455), .ZN(n477) );
  INV_X1 U457 ( .A(n716), .ZN(n455) );
  NOR2_X1 U458 ( .A1(n431), .A2(n430), .ZN(n429) );
  NOR2_X1 U459 ( .A1(n433), .A2(n435), .ZN(n428) );
  INV_X1 U460 ( .A(n719), .ZN(n402) );
  AND2_X1 U461 ( .A1(n405), .A2(n404), .ZN(n403) );
  NOR2_X2 U462 ( .A1(n398), .A2(n395), .ZN(n384) );
  NAND2_X1 U463 ( .A1(n400), .A2(n399), .ZN(n398) );
  NAND2_X1 U464 ( .A1(n564), .A2(n397), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n557), .B(n487), .ZN(n486) );
  XNOR2_X1 U466 ( .A(n558), .B(KEYINPUT111), .ZN(n487) );
  NAND2_X1 U467 ( .A1(n366), .A2(n379), .ZN(n557) );
  OR2_X1 U468 ( .A1(n619), .A2(n412), .ZN(n411) );
  AND2_X1 U469 ( .A1(n415), .A2(n414), .ZN(n413) );
  BUF_X1 U470 ( .A(n694), .Z(n451) );
  XNOR2_X1 U471 ( .A(n359), .B(n535), .ZN(n385) );
  NOR2_X1 U472 ( .A1(G952), .A2(n758), .ZN(n749) );
  NAND2_X1 U473 ( .A1(n780), .A2(KEYINPUT46), .ZN(n423) );
  AND2_X1 U474 ( .A1(n710), .A2(KEYINPUT19), .ZN(n448) );
  XOR2_X1 U475 ( .A(KEYINPUT97), .B(G140), .Z(n504) );
  XNOR2_X1 U476 ( .A(n441), .B(G131), .ZN(n547) );
  INV_X1 U477 ( .A(KEYINPUT66), .ZN(n441) );
  XNOR2_X1 U478 ( .A(n507), .B(KEYINPUT12), .ZN(n440) );
  INV_X1 U479 ( .A(KEYINPUT11), .ZN(n507) );
  XNOR2_X1 U480 ( .A(n505), .B(n501), .ZN(n506) );
  XOR2_X1 U481 ( .A(G113), .B(G143), .Z(n501) );
  XNOR2_X1 U482 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U483 ( .A(G104), .B(G122), .ZN(n503) );
  INV_X1 U484 ( .A(KEYINPUT79), .ZN(n497) );
  XNOR2_X1 U485 ( .A(n771), .B(KEYINPUT72), .ZN(n498) );
  XOR2_X1 U486 ( .A(G902), .B(KEYINPUT15), .Z(n647) );
  NAND2_X1 U487 ( .A1(G234), .A2(G237), .ZN(n541) );
  XNOR2_X1 U488 ( .A(n594), .B(n478), .ZN(n716) );
  INV_X1 U489 ( .A(KEYINPUT113), .ZN(n478) );
  NOR2_X1 U490 ( .A1(n432), .A2(n434), .ZN(n430) );
  AND2_X1 U491 ( .A1(n711), .A2(n356), .ZN(n432) );
  INV_X1 U492 ( .A(G902), .ZN(n397) );
  NAND2_X1 U493 ( .A1(G469), .A2(G902), .ZN(n399) );
  INV_X1 U494 ( .A(KEYINPUT22), .ZN(n417) );
  XNOR2_X1 U495 ( .A(n462), .B(n453), .ZN(n551) );
  XNOR2_X1 U496 ( .A(n571), .B(n362), .ZN(n554) );
  XNOR2_X1 U497 ( .A(G119), .B(G128), .ZN(n526) );
  XNOR2_X1 U498 ( .A(n380), .B(G110), .ZN(n527) );
  INV_X1 U499 ( .A(KEYINPUT92), .ZN(n380) );
  XOR2_X1 U500 ( .A(KEYINPUT23), .B(KEYINPUT91), .Z(n528) );
  XNOR2_X1 U501 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n457) );
  XNOR2_X1 U502 ( .A(n767), .B(n459), .ZN(n563) );
  XNOR2_X1 U503 ( .A(n562), .B(n460), .ZN(n459) );
  XNOR2_X1 U504 ( .A(n559), .B(n755), .ZN(n565) );
  XNOR2_X1 U505 ( .A(n393), .B(KEYINPUT67), .ZN(n559) );
  XNOR2_X1 U506 ( .A(n409), .B(n408), .ZN(n456) );
  INV_X1 U507 ( .A(KEYINPUT17), .ZN(n408) );
  NAND2_X1 U508 ( .A1(n410), .A2(G224), .ZN(n409) );
  INV_X1 U509 ( .A(G953), .ZN(n410) );
  XNOR2_X1 U510 ( .A(KEYINPUT18), .B(KEYINPUT75), .ZN(n490) );
  XNOR2_X1 U511 ( .A(G122), .B(KEYINPUT16), .ZN(n570) );
  XNOR2_X1 U512 ( .A(n439), .B(n494), .ZN(n493) );
  INV_X1 U513 ( .A(KEYINPUT81), .ZN(n494) );
  BUF_X1 U514 ( .A(n719), .Z(n418) );
  XNOR2_X1 U515 ( .A(n577), .B(n437), .ZN(n436) );
  INV_X1 U516 ( .A(KEYINPUT30), .ZN(n437) );
  BUF_X2 U517 ( .A(n603), .Z(n458) );
  XNOR2_X1 U518 ( .A(n513), .B(G475), .ZN(n442) );
  XNOR2_X1 U519 ( .A(n655), .B(KEYINPUT62), .ZN(n657) );
  XNOR2_X1 U520 ( .A(n517), .B(n470), .ZN(n519) );
  XOR2_X1 U521 ( .A(n661), .B(KEYINPUT59), .Z(n663) );
  INV_X1 U522 ( .A(n771), .ZN(n729) );
  XNOR2_X1 U523 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n454) );
  NAND2_X1 U524 ( .A1(n486), .A2(n376), .ZN(n595) );
  INV_X1 U525 ( .A(KEYINPUT35), .ZN(n406) );
  NAND2_X1 U526 ( .A1(n402), .A2(n357), .ZN(n401) );
  XNOR2_X1 U527 ( .A(n631), .B(KEYINPUT105), .ZN(n387) );
  XNOR2_X1 U528 ( .A(n482), .B(n481), .ZN(n685) );
  XNOR2_X1 U529 ( .A(KEYINPUT96), .B(KEYINPUT31), .ZN(n481) );
  INV_X1 U530 ( .A(KEYINPUT77), .ZN(n381) );
  NAND2_X1 U531 ( .A1(n486), .A2(n383), .ZN(n382) );
  XNOR2_X1 U532 ( .A(n628), .B(KEYINPUT107), .ZN(n782) );
  NAND2_X1 U533 ( .A1(n605), .A2(n500), .ZN(n499) );
  XNOR2_X1 U534 ( .A(n747), .B(n385), .ZN(n748) );
  NOR2_X1 U535 ( .A1(n710), .A2(KEYINPUT19), .ZN(n355) );
  AND2_X1 U536 ( .A1(n367), .A2(n583), .ZN(n356) );
  NOR2_X1 U537 ( .A1(n638), .A2(n369), .ZN(n357) );
  AND2_X1 U538 ( .A1(n638), .A2(n369), .ZN(n358) );
  XOR2_X1 U539 ( .A(n534), .B(n533), .Z(n359) );
  XOR2_X1 U540 ( .A(KEYINPUT93), .B(n696), .Z(n360) );
  OR2_X1 U541 ( .A1(n612), .A2(n611), .ZN(n361) );
  AND2_X1 U542 ( .A1(G210), .A2(n553), .ZN(n362) );
  AND2_X1 U543 ( .A1(n436), .A2(n356), .ZN(n363) );
  XOR2_X1 U544 ( .A(n573), .B(n572), .Z(n364) );
  INV_X1 U545 ( .A(n697), .ZN(n630) );
  AND2_X1 U546 ( .A1(n502), .A2(KEYINPUT2), .ZN(n365) );
  AND2_X1 U547 ( .A1(n556), .A2(n583), .ZN(n366) );
  AND2_X1 U548 ( .A1(n693), .A2(n376), .ZN(n367) );
  AND2_X1 U549 ( .A1(n360), .A2(n417), .ZN(n368) );
  XNOR2_X1 U550 ( .A(KEYINPUT68), .B(KEYINPUT34), .ZN(n369) );
  INV_X1 U551 ( .A(KEYINPUT39), .ZN(n434) );
  XOR2_X1 U552 ( .A(KEYINPUT45), .B(KEYINPUT80), .Z(n370) );
  NAND2_X1 U553 ( .A1(n647), .A2(KEYINPUT2), .ZN(n371) );
  INV_X1 U554 ( .A(n384), .ZN(n376) );
  XNOR2_X1 U555 ( .A(n377), .B(G119), .ZN(G21) );
  XNOR2_X2 U556 ( .A(n386), .B(KEYINPUT32), .ZN(n377) );
  NOR2_X2 U557 ( .A1(n378), .A2(n616), .ZN(n632) );
  NOR2_X1 U558 ( .A1(n378), .A2(n499), .ZN(n628) );
  NAND2_X1 U559 ( .A1(n379), .A2(n710), .ZN(n577) );
  NOR2_X1 U560 ( .A1(n379), .A2(n697), .ZN(n500) );
  NOR2_X1 U561 ( .A1(n575), .A2(n384), .ZN(n383) );
  NOR2_X1 U562 ( .A1(n385), .A2(G902), .ZN(n538) );
  NAND2_X1 U563 ( .A1(n632), .A2(n387), .ZN(n386) );
  NAND2_X1 U564 ( .A1(n390), .A2(n388), .ZN(n450) );
  NAND2_X1 U565 ( .A1(KEYINPUT44), .A2(n634), .ZN(n389) );
  NAND2_X1 U566 ( .A1(n391), .A2(n634), .ZN(n390) );
  INV_X1 U567 ( .A(n392), .ZN(n391) );
  XNOR2_X1 U568 ( .A(n641), .B(KEYINPUT84), .ZN(n392) );
  XNOR2_X1 U569 ( .A(n550), .B(n393), .ZN(n453) );
  XNOR2_X2 U570 ( .A(n452), .B(G101), .ZN(n393) );
  NAND2_X1 U571 ( .A1(n619), .A2(KEYINPUT22), .ZN(n415) );
  NOR2_X2 U572 ( .A1(n658), .A2(n749), .ZN(n660) );
  XNOR2_X2 U573 ( .A(n394), .B(G128), .ZN(n567) );
  NOR2_X1 U574 ( .A1(n736), .A2(n396), .ZN(n395) );
  NAND2_X1 U575 ( .A1(n736), .A2(G469), .ZN(n400) );
  NAND2_X1 U576 ( .A1(n719), .A2(n369), .ZN(n404) );
  NOR2_X1 U577 ( .A1(n358), .A2(n640), .ZN(n405) );
  XNOR2_X2 U578 ( .A(n407), .B(n406), .ZN(n779) );
  NAND2_X1 U579 ( .A1(n615), .A2(n368), .ZN(n412) );
  NAND2_X1 U580 ( .A1(n416), .A2(KEYINPUT22), .ZN(n414) );
  NAND2_X1 U581 ( .A1(n615), .A2(n360), .ZN(n416) );
  XNOR2_X2 U582 ( .A(n419), .B(KEYINPUT70), .ZN(n635) );
  NAND2_X1 U583 ( .A1(n783), .A2(KEYINPUT46), .ZN(n421) );
  INV_X1 U584 ( .A(n780), .ZN(n425) );
  XNOR2_X2 U585 ( .A(n596), .B(n454), .ZN(n783) );
  NAND2_X1 U586 ( .A1(n356), .A2(n434), .ZN(n433) );
  NAND2_X1 U587 ( .A1(n429), .A2(n427), .ZN(n599) );
  NAND2_X1 U588 ( .A1(n436), .A2(n428), .ZN(n427) );
  INV_X1 U589 ( .A(n711), .ZN(n435) );
  NAND2_X1 U590 ( .A1(n438), .A2(n365), .ZN(n439) );
  XNOR2_X2 U591 ( .A(n443), .B(n442), .ZN(n591) );
  NAND2_X1 U592 ( .A1(n458), .A2(n710), .ZN(n606) );
  NAND2_X1 U593 ( .A1(n603), .A2(n448), .ZN(n447) );
  XNOR2_X2 U594 ( .A(n475), .B(n364), .ZN(n603) );
  XNOR2_X1 U595 ( .A(n656), .B(n657), .ZN(n658) );
  XNOR2_X1 U596 ( .A(n662), .B(n663), .ZN(n664) );
  XNOR2_X1 U597 ( .A(n530), .B(n766), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n625), .B(KEYINPUT104), .ZN(n627) );
  XNOR2_X1 U599 ( .A(n554), .B(n551), .ZN(n485) );
  NOR2_X1 U600 ( .A1(n655), .A2(G902), .ZN(n555) );
  XNOR2_X1 U601 ( .A(n555), .B(G472), .ZN(n621) );
  XNOR2_X1 U602 ( .A(n485), .B(n560), .ZN(n655) );
  NAND2_X1 U603 ( .A1(n450), .A2(n479), .ZN(n491) );
  XNOR2_X1 U604 ( .A(n491), .B(n370), .ZN(n648) );
  XNOR2_X1 U605 ( .A(n456), .B(n490), .ZN(n569) );
  XNOR2_X1 U606 ( .A(n632), .B(KEYINPUT82), .ZN(n617) );
  AND2_X1 U607 ( .A1(n627), .A2(n626), .ZN(n466) );
  OR2_X2 U608 ( .A1(n650), .A2(n647), .ZN(n475) );
  XNOR2_X1 U609 ( .A(n569), .B(n568), .ZN(n489) );
  XNOR2_X1 U610 ( .A(n565), .B(n489), .ZN(n488) );
  NOR2_X2 U611 ( .A1(n648), .A2(n645), .ZN(n646) );
  XNOR2_X1 U612 ( .A(n488), .B(n756), .ZN(n650) );
  NAND2_X1 U613 ( .A1(n739), .A2(G210), .ZN(n652) );
  NOR2_X2 U614 ( .A1(n653), .A2(n749), .ZN(n654) );
  NAND2_X1 U615 ( .A1(n644), .A2(KEYINPUT44), .ZN(n467) );
  NAND2_X1 U616 ( .A1(n739), .A2(G475), .ZN(n662) );
  NAND2_X1 U617 ( .A1(n461), .A2(n590), .ZN(n484) );
  BUF_X2 U618 ( .A(n621), .Z(n464) );
  NAND2_X1 U619 ( .A1(n496), .A2(n498), .ZN(n465) );
  XNOR2_X2 U620 ( .A(n458), .B(n474), .ZN(n711) );
  INV_X1 U621 ( .A(n615), .ZN(n713) );
  NOR2_X2 U622 ( .A1(n709), .A2(n595), .ZN(n596) );
  INV_X1 U623 ( .A(n694), .ZN(n605) );
  XNOR2_X1 U624 ( .A(n565), .B(n563), .ZN(n480) );
  NAND2_X1 U625 ( .A1(n705), .A2(n620), .ZN(n482) );
  NOR2_X2 U626 ( .A1(n635), .A2(n464), .ZN(n705) );
  NOR2_X2 U627 ( .A1(n664), .A2(n749), .ZN(n666) );
  INV_X1 U628 ( .A(n492), .ZN(n732) );
  XNOR2_X1 U629 ( .A(n646), .B(n497), .ZN(n496) );
  XNOR2_X1 U630 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X1 U631 ( .A1(n604), .A2(n691), .ZN(n502) );
  BUF_X1 U632 ( .A(n641), .Z(n642) );
  INV_X1 U633 ( .A(G469), .ZN(n564) );
  XNOR2_X1 U634 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U635 ( .A(KEYINPUT63), .ZN(n659) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT64), .ZN(n665) );
  XNOR2_X1 U637 ( .A(KEYINPUT98), .B(KEYINPUT13), .ZN(n513) );
  XOR2_X2 U638 ( .A(G146), .B(G125), .Z(n566) );
  XNOR2_X1 U639 ( .A(n766), .B(n506), .ZN(n512) );
  XOR2_X1 U640 ( .A(KEYINPUT73), .B(n508), .Z(n553) );
  NAND2_X1 U641 ( .A1(G214), .A2(n553), .ZN(n509) );
  XNOR2_X1 U642 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n524) );
  XNOR2_X2 U643 ( .A(n567), .B(n514), .ZN(n548) );
  XOR2_X1 U644 ( .A(KEYINPUT7), .B(KEYINPUT99), .Z(n516) );
  XNOR2_X1 U645 ( .A(G107), .B(KEYINPUT9), .ZN(n515) );
  XNOR2_X1 U646 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U647 ( .A(n519), .B(n548), .Z(n522) );
  NAND2_X1 U648 ( .A1(G234), .A2(n758), .ZN(n520) );
  XOR2_X1 U649 ( .A(KEYINPUT8), .B(n520), .Z(n532) );
  NAND2_X1 U650 ( .A1(G217), .A2(n532), .ZN(n521) );
  XNOR2_X1 U651 ( .A(n522), .B(n521), .ZN(n744) );
  INV_X1 U652 ( .A(n592), .ZN(n525) );
  NOR2_X1 U653 ( .A1(n591), .A2(n525), .ZN(n682) );
  NAND2_X1 U654 ( .A1(n525), .A2(n591), .ZN(n674) );
  INV_X1 U655 ( .A(n674), .ZN(n684) );
  NOR2_X1 U656 ( .A1(n682), .A2(n684), .ZN(n715) );
  XNOR2_X1 U657 ( .A(n527), .B(n526), .ZN(n529) );
  INV_X1 U658 ( .A(n561), .ZN(n531) );
  XOR2_X1 U659 ( .A(n531), .B(KEYINPUT24), .Z(n534) );
  NAND2_X1 U660 ( .A1(G221), .A2(n532), .ZN(n533) );
  INV_X1 U661 ( .A(n647), .ZN(n645) );
  NAND2_X1 U662 ( .A1(n645), .A2(G234), .ZN(n536) );
  XNOR2_X1 U663 ( .A(n536), .B(KEYINPUT20), .ZN(n539) );
  NAND2_X1 U664 ( .A1(n539), .A2(G217), .ZN(n537) );
  NAND2_X1 U665 ( .A1(G221), .A2(n539), .ZN(n540) );
  XOR2_X1 U666 ( .A(KEYINPUT21), .B(n540), .Z(n696) );
  NAND2_X1 U667 ( .A1(n630), .A2(n696), .ZN(n585) );
  INV_X1 U668 ( .A(n585), .ZN(n556) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n541), .Z(n612) );
  INV_X1 U670 ( .A(n612), .ZN(n724) );
  NAND2_X1 U671 ( .A1(G953), .A2(G902), .ZN(n608) );
  NOR2_X1 U672 ( .A1(G900), .A2(n608), .ZN(n542) );
  NAND2_X1 U673 ( .A1(n724), .A2(n542), .ZN(n543) );
  XNOR2_X1 U674 ( .A(n543), .B(KEYINPUT109), .ZN(n545) );
  NAND2_X1 U675 ( .A1(n758), .A2(G952), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n612), .A2(n607), .ZN(n544) );
  NOR2_X1 U677 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U678 ( .A(KEYINPUT78), .B(n546), .Z(n583) );
  XOR2_X1 U679 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n550) );
  INV_X1 U680 ( .A(n621), .ZN(n703) );
  XNOR2_X1 U681 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n558) );
  XNOR2_X1 U682 ( .A(KEYINPUT90), .B(n561), .ZN(n767) );
  NAND2_X1 U683 ( .A1(G227), .A2(n758), .ZN(n562) );
  XNOR2_X1 U684 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U685 ( .A(n571), .B(n570), .ZN(n756) );
  NAND2_X1 U686 ( .A1(G210), .A2(n574), .ZN(n573) );
  NAND2_X1 U687 ( .A1(G214), .A2(n574), .ZN(n710) );
  XOR2_X1 U688 ( .A(n606), .B(KEYINPUT19), .Z(n575) );
  XNOR2_X1 U689 ( .A(n576), .B(KEYINPUT47), .ZN(n581) );
  OR2_X1 U690 ( .A1(n592), .A2(n591), .ZN(n578) );
  XNOR2_X1 U691 ( .A(n578), .B(KEYINPUT108), .ZN(n639) );
  INV_X1 U692 ( .A(n458), .ZN(n579) );
  NOR2_X1 U693 ( .A1(n639), .A2(n579), .ZN(n580) );
  NAND2_X1 U694 ( .A1(n363), .A2(n580), .ZN(n677) );
  NAND2_X1 U695 ( .A1(n581), .A2(n677), .ZN(n582) );
  XNOR2_X1 U696 ( .A(n582), .B(KEYINPUT69), .ZN(n590) );
  XOR2_X1 U697 ( .A(KEYINPUT6), .B(n464), .Z(n636) );
  NAND2_X1 U698 ( .A1(n583), .A2(n710), .ZN(n584) );
  NOR2_X1 U699 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U700 ( .A1(n682), .A2(n586), .ZN(n587) );
  NOR2_X1 U701 ( .A1(n636), .A2(n587), .ZN(n600) );
  AND2_X1 U702 ( .A1(n458), .A2(n600), .ZN(n588) );
  XNOR2_X1 U703 ( .A(n588), .B(KEYINPUT36), .ZN(n589) );
  XNOR2_X1 U704 ( .A(n605), .B(KEYINPUT87), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n589), .A2(n629), .ZN(n688) );
  NAND2_X1 U706 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X2 U707 ( .A(n593), .B(KEYINPUT103), .ZN(n615) );
  NAND2_X1 U708 ( .A1(n711), .A2(n710), .ZN(n594) );
  XOR2_X1 U709 ( .A(KEYINPUT40), .B(KEYINPUT112), .Z(n598) );
  NAND2_X1 U710 ( .A1(n599), .A2(n682), .ZN(n597) );
  NAND2_X1 U711 ( .A1(n684), .A2(n599), .ZN(n690) );
  NAND2_X1 U712 ( .A1(n605), .A2(n600), .ZN(n601) );
  XOR2_X1 U713 ( .A(KEYINPUT43), .B(n601), .Z(n602) );
  NOR2_X1 U714 ( .A1(n458), .A2(n602), .ZN(n691) );
  INV_X1 U715 ( .A(n607), .ZN(n610) );
  NOR2_X1 U716 ( .A1(G898), .A2(n608), .ZN(n609) );
  NOR2_X1 U717 ( .A1(n610), .A2(n609), .ZN(n611) );
  INV_X1 U718 ( .A(n636), .ZN(n616) );
  NAND2_X1 U719 ( .A1(n617), .A2(n697), .ZN(n618) );
  BUF_X1 U720 ( .A(n619), .Z(n638) );
  INV_X1 U721 ( .A(n638), .ZN(n620) );
  NAND2_X1 U722 ( .A1(n367), .A2(n464), .ZN(n622) );
  NOR2_X1 U723 ( .A1(n638), .A2(n622), .ZN(n670) );
  NOR2_X1 U724 ( .A1(n685), .A2(n670), .ZN(n623) );
  NOR2_X1 U725 ( .A1(n715), .A2(n623), .ZN(n624) );
  NOR2_X1 U726 ( .A1(n667), .A2(n624), .ZN(n625) );
  INV_X1 U727 ( .A(KEYINPUT83), .ZN(n634) );
  OR2_X1 U728 ( .A1(KEYINPUT44), .A2(n634), .ZN(n626) );
  NAND2_X1 U729 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X2 U730 ( .A(n633), .B(KEYINPUT85), .ZN(n641) );
  XNOR2_X1 U731 ( .A(KEYINPUT76), .B(n639), .ZN(n640) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U733 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n649) );
  XNOR2_X1 U734 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U735 ( .A(n654), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U736 ( .A1(n739), .A2(G472), .ZN(n656) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(G57) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(G60) );
  XNOR2_X1 U739 ( .A(G101), .B(n667), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT115), .ZN(G3) );
  NAND2_X1 U741 ( .A1(n670), .A2(n682), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(G104), .ZN(G6) );
  XOR2_X1 U743 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n672) );
  NAND2_X1 U744 ( .A1(n670), .A2(n684), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U746 ( .A(G107), .B(n673), .ZN(G9) );
  NOR2_X1 U747 ( .A1(n674), .A2(n678), .ZN(n676) );
  XNOR2_X1 U748 ( .A(G128), .B(KEYINPUT29), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(G30) );
  XNOR2_X1 U750 ( .A(G143), .B(n677), .ZN(G45) );
  INV_X1 U751 ( .A(n682), .ZN(n679) );
  NOR2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U753 ( .A(G146), .B(n680), .Z(n681) );
  XNOR2_X1 U754 ( .A(KEYINPUT116), .B(n681), .ZN(G48) );
  NAND2_X1 U755 ( .A1(n685), .A2(n682), .ZN(n683) );
  XNOR2_X1 U756 ( .A(n683), .B(G113), .ZN(G15) );
  NAND2_X1 U757 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(G116), .ZN(G18) );
  XOR2_X1 U759 ( .A(G125), .B(KEYINPUT37), .Z(n687) );
  XNOR2_X1 U760 ( .A(n688), .B(n687), .ZN(G27) );
  XOR2_X1 U761 ( .A(G134), .B(KEYINPUT117), .Z(n689) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(G36) );
  XOR2_X1 U763 ( .A(G140), .B(n691), .Z(G42) );
  NOR2_X1 U764 ( .A1(n418), .A2(n709), .ZN(n692) );
  NOR2_X1 U765 ( .A1(G953), .A2(n692), .ZN(n728) );
  OR2_X1 U766 ( .A1(n451), .A2(n693), .ZN(n695) );
  XNOR2_X1 U767 ( .A(KEYINPUT50), .B(n695), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n697), .A2(n696), .ZN(n699) );
  XNOR2_X1 U769 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n698) );
  XNOR2_X1 U770 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U772 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U774 ( .A(n706), .B(KEYINPUT51), .ZN(n707) );
  XNOR2_X1 U775 ( .A(KEYINPUT119), .B(n707), .ZN(n708) );
  NOR2_X1 U776 ( .A1(n709), .A2(n708), .ZN(n722) );
  NOR2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U779 ( .A(n714), .B(KEYINPUT120), .ZN(n718) );
  NOR2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n720), .A2(n418), .ZN(n721) );
  NOR2_X1 U783 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U784 ( .A(KEYINPUT52), .B(n723), .Z(n726) );
  AND2_X1 U785 ( .A1(G952), .A2(n724), .ZN(n725) );
  NAND2_X1 U786 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U787 ( .A1(n728), .A2(n727), .ZN(n734) );
  NOR2_X1 U788 ( .A1(n729), .A2(n750), .ZN(n730) );
  NOR2_X1 U789 ( .A1(KEYINPUT2), .A2(n730), .ZN(n731) );
  NOR2_X1 U790 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U791 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U792 ( .A(n735), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U793 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n738) );
  XNOR2_X1 U794 ( .A(n736), .B(KEYINPUT57), .ZN(n737) );
  XNOR2_X1 U795 ( .A(n738), .B(n737), .ZN(n741) );
  NAND2_X1 U796 ( .A1(n746), .A2(G469), .ZN(n740) );
  XNOR2_X1 U797 ( .A(n741), .B(n740), .ZN(n742) );
  NOR2_X1 U798 ( .A1(n749), .A2(n742), .ZN(G54) );
  NAND2_X1 U799 ( .A1(G478), .A2(n746), .ZN(n743) );
  XNOR2_X1 U800 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U801 ( .A1(n749), .A2(n745), .ZN(G63) );
  NAND2_X1 U802 ( .A1(G217), .A2(n746), .ZN(n747) );
  NOR2_X1 U803 ( .A1(n749), .A2(n748), .ZN(G66) );
  OR2_X1 U804 ( .A1(G953), .A2(n750), .ZN(n754) );
  NAND2_X1 U805 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U807 ( .A1(n752), .A2(G898), .ZN(n753) );
  NAND2_X1 U808 ( .A1(n754), .A2(n753), .ZN(n762) );
  XNOR2_X1 U809 ( .A(G101), .B(n755), .ZN(n757) );
  XNOR2_X1 U810 ( .A(n757), .B(n756), .ZN(n760) );
  NOR2_X1 U811 ( .A1(G898), .A2(n758), .ZN(n759) );
  NOR2_X1 U812 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U813 ( .A(n762), .B(n761), .ZN(n763) );
  XNOR2_X1 U814 ( .A(KEYINPUT122), .B(n763), .ZN(G69) );
  XNOR2_X1 U815 ( .A(KEYINPUT4), .B(KEYINPUT123), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n764), .B(KEYINPUT124), .ZN(n765) );
  XNOR2_X1 U817 ( .A(n766), .B(n765), .ZN(n770) );
  XNOR2_X1 U818 ( .A(n768), .B(n767), .ZN(n769) );
  XOR2_X1 U819 ( .A(n770), .B(n769), .Z(n774) );
  XNOR2_X1 U820 ( .A(n774), .B(n771), .ZN(n772) );
  NOR2_X1 U821 ( .A1(G953), .A2(n772), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n773), .B(KEYINPUT125), .ZN(n778) );
  XNOR2_X1 U823 ( .A(G227), .B(n774), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(G900), .ZN(n776) );
  NAND2_X1 U825 ( .A1(G953), .A2(n776), .ZN(n777) );
  NAND2_X1 U826 ( .A1(n778), .A2(n777), .ZN(G72) );
  XNOR2_X1 U827 ( .A(G122), .B(n779), .ZN(G24) );
  XNOR2_X1 U828 ( .A(n780), .B(G131), .ZN(n781) );
  XNOR2_X1 U829 ( .A(n781), .B(KEYINPUT127), .ZN(G33) );
  XNOR2_X1 U830 ( .A(G110), .B(n782), .ZN(G12) );
  XOR2_X1 U831 ( .A(n783), .B(G137), .Z(n784) );
  XNOR2_X1 U832 ( .A(KEYINPUT126), .B(n784), .ZN(G39) );
endmodule

