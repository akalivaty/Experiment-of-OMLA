//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n561, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n621, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1246;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AND2_X1   g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n456), .A2(new_n457), .B1(G567), .B2(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n465), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n470), .B2(G2105), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g052(.A1(new_n477), .A2(KEYINPUT66), .A3(G137), .A4(new_n462), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n471), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n468), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n468), .A2(new_n462), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT67), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g061(.A1(KEYINPUT67), .A2(G100), .A3(G2105), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n462), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  AND3_X1   g063(.A1(new_n482), .A2(new_n484), .A3(new_n488), .ZN(G162));
  INV_X1    g064(.A(G126), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n475), .B2(new_n476), .ZN(new_n491));
  AND2_X1   g066(.A1(G114), .A2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n462), .C1(new_n466), .C2(new_n467), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n477), .A2(new_n498), .B1(G102), .B2(G2104), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n493), .B(new_n496), .C1(G2105), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n502), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT69), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(G62), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G166));
  OAI21_X1  g099(.A(G543), .B1(new_n503), .B2(new_n504), .ZN(new_n525));
  INV_X1    g100(.A(new_n510), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n527), .A2(G89), .A3(new_n505), .A4(new_n518), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT71), .B(G51), .ZN(new_n529));
  INV_X1    g104(.A(new_n517), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT6), .A2(G651), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT70), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n516), .B2(new_n517), .ZN(new_n534));
  OAI211_X1 g109(.A(G543), .B(new_n529), .C1(new_n532), .C2(new_n534), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n505), .B(new_n536), .C1(new_n509), .C2(new_n510), .ZN(new_n537));
  NAND3_X1  g112(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n538), .B(KEYINPUT7), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n528), .A2(new_n535), .A3(new_n537), .A4(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND3_X1  g116(.A1(new_n527), .A2(G64), .A3(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n515), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n527), .A2(G90), .A3(new_n505), .A4(new_n518), .ZN(new_n545));
  OAI211_X1 g120(.A(G52), .B(G543), .C1(new_n532), .C2(new_n534), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  XOR2_X1   g123(.A(KEYINPUT72), .B(G81), .Z(new_n549));
  NAND4_X1  g124(.A1(new_n527), .A2(new_n505), .A3(new_n518), .A4(new_n549), .ZN(new_n550));
  OAI211_X1 g125(.A(G43), .B(G543), .C1(new_n532), .C2(new_n534), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT73), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT73), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n550), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n511), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n553), .A2(new_n555), .B1(G651), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  INV_X1    g141(.A(G78), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n511), .A2(new_n566), .B1(new_n567), .B2(new_n506), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT74), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  OAI221_X1 g145(.A(new_n570), .B1(new_n567), .B2(new_n506), .C1(new_n511), .C2(new_n566), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G651), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n534), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n516), .A2(new_n533), .A3(new_n517), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n506), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n575), .A2(new_n576), .A3(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(G543), .B1(new_n532), .B2(new_n534), .ZN(new_n578));
  INV_X1    g153(.A(G53), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT9), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n527), .A2(new_n505), .A3(new_n518), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n577), .A2(new_n580), .B1(G91), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n572), .A2(new_n583), .ZN(G299));
  INV_X1    g159(.A(G171), .ZN(G301));
  OR2_X1    g160(.A1(new_n520), .A2(new_n523), .ZN(G303));
  OAI21_X1  g161(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n582), .A2(G87), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n575), .A2(G49), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G288));
  OAI211_X1 g165(.A(new_n505), .B(G61), .C1(new_n509), .C2(new_n510), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT75), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n593), .A2(new_n596), .A3(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(G48), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n511), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n518), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n582), .A2(G85), .B1(new_n575), .B2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n511), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(G290));
  NAND4_X1  g183(.A1(new_n527), .A2(G92), .A3(new_n505), .A4(new_n518), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n511), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(G54), .B2(new_n575), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G868), .ZN(new_n617));
  MUX2_X1   g192(.A(G301), .B(new_n616), .S(new_n617), .Z(G284));
  MUX2_X1   g193(.A(G301), .B(new_n616), .S(new_n617), .Z(G321));
  NAND2_X1  g194(.A1(G168), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G299), .B2(G868), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(G297));
  XNOR2_X1  g197(.A(new_n621), .B(KEYINPUT76), .ZN(G280));
  AND2_X1   g198(.A1(new_n611), .A2(new_n615), .ZN(new_n624));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n558), .A2(G651), .ZN(new_n627));
  INV_X1    g202(.A(new_n555), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n554), .B1(new_n550), .B2(new_n551), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n624), .A2(new_n625), .ZN(new_n631));
  MUX2_X1   g206(.A(new_n630), .B(new_n631), .S(G868), .Z(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n481), .A2(G135), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT77), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n483), .A2(G123), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n638));
  AND2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI22_X1  g214(.A1(new_n637), .A2(new_n638), .B1(G111), .B2(new_n462), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n635), .B(new_n636), .C1(new_n639), .C2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT12), .Z(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT13), .Z(new_n646));
  INV_X1    g221(.A(G2100), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n648), .A3(new_n649), .ZN(G156));
  XOR2_X1   g225(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n654), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n657), .A3(new_n651), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n660), .A2(new_n662), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT15), .B(G2435), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT81), .B(G2438), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2427), .B(G2430), .ZN(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  INV_X1    g249(.A(KEYINPUT14), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n668), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n666), .A2(new_n676), .A3(new_n667), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(G14), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  OAI21_X1  g260(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n685), .A2(new_n682), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n686), .B(new_n687), .C1(new_n690), .C2(new_n683), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n685), .A2(new_n683), .A3(new_n682), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT82), .B(KEYINPUT18), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n691), .A2(KEYINPUT83), .A3(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2096), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n642), .A3(new_n698), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(new_n647), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(G2100), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(G227));
  XNOR2_X1  g280(.A(G1971), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1956), .B(G2474), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1961), .B(G1966), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT20), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n709), .A2(new_n710), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n708), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT85), .ZN(new_n716));
  OR3_X1    g291(.A1(new_n708), .A2(new_n714), .A3(new_n711), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n713), .A2(new_n716), .A3(new_n717), .A4(new_n719), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1991), .B(G1996), .ZN(new_n723));
  XNOR2_X1  g298(.A(G1981), .B(G1986), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n721), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n721), .B2(new_n722), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(G229));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  AND2_X1   g305(.A1(KEYINPUT24), .A2(G34), .ZN(new_n731));
  NOR2_X1   g306(.A1(KEYINPUT24), .A2(G34), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n479), .B2(new_n730), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n737));
  AND2_X1   g312(.A1(G115), .A2(G2104), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n477), .B2(G127), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(new_n739), .B2(new_n462), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n481), .A2(G139), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n739), .A2(new_n737), .A3(new_n462), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G29), .B2(G33), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G2072), .ZN(new_n751));
  OR2_X1    g326(.A1(G29), .A2(G32), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n483), .A2(G129), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT98), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT98), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n483), .A2(new_n755), .A3(G129), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AND3_X1   g332(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n758));
  NAND3_X1  g333(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT26), .ZN(new_n760));
  AOI211_X1 g335(.A(new_n758), .B(new_n760), .C1(G141), .C2(new_n481), .ZN(new_n761));
  AOI21_X1  g336(.A(KEYINPUT99), .B1(new_n757), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n757), .A2(new_n761), .A3(KEYINPUT99), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n752), .B1(new_n765), .B2(new_n730), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT100), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n736), .B(new_n751), .C1(new_n767), .C2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT101), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NOR2_X1   g348(.A1(G4), .A2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT93), .ZN(new_n775));
  INV_X1    g350(.A(G16), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n616), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n776), .A2(G5), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G171), .B2(new_n776), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1961), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT102), .Z(new_n783));
  AOI211_X1 g358(.A(new_n779), .B(new_n783), .C1(new_n767), .C2(new_n769), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n772), .A2(new_n773), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G35), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G162), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT103), .B(KEYINPUT29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2090), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n730), .A2(G26), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT96), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT28), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G128), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT95), .ZN(new_n795));
  MUX2_X1   g370(.A(G104), .B(G116), .S(G2105), .Z(new_n796));
  AOI22_X1  g371(.A1(new_n481), .A2(G140), .B1(G2104), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n793), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G2067), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n790), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n781), .A2(G1961), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT31), .B(G11), .Z(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT30), .B(G28), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n803), .B1(new_n730), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G27), .A2(G29), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G164), .B2(G29), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n805), .B1(G2078), .B2(new_n807), .C1(new_n641), .C2(new_n730), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n807), .A2(G2078), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n734), .A2(new_n735), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n801), .A2(new_n802), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G19), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n813), .B1(new_n559), .B2(G16), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT94), .B(G1341), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT104), .B(KEYINPUT23), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n776), .A2(G20), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G299), .B2(G16), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(G1956), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n776), .A2(G21), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G168), .B2(new_n776), .ZN(new_n823));
  INV_X1    g398(.A(G1966), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n812), .A2(new_n816), .A3(new_n821), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n785), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G16), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(G6), .B2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT89), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT32), .B(G1981), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT90), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT89), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n831), .B(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n834), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G16), .A2(G22), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(G166), .B2(G16), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(G1971), .ZN(new_n842));
  NOR2_X1   g417(.A1(G16), .A2(G23), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT91), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n844), .B1(G288), .B2(new_n776), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT33), .B(G1976), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n835), .A2(new_n839), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(KEYINPUT34), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT34), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n835), .A2(new_n839), .A3(new_n851), .A4(new_n848), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n730), .A2(G25), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n481), .A2(G131), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n854), .B(KEYINPUT86), .Z(new_n855));
  MUX2_X1   g430(.A(G95), .B(G107), .S(G2105), .Z(new_n856));
  AOI22_X1  g431(.A1(new_n483), .A2(G119), .B1(G2104), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT87), .Z(new_n859));
  AOI21_X1  g434(.A(new_n853), .B1(new_n859), .B2(G29), .ZN(new_n860));
  XOR2_X1   g435(.A(KEYINPUT35), .B(G1991), .Z(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT88), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n860), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(G16), .A2(G24), .ZN(new_n864));
  INV_X1    g439(.A(G290), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(G16), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(G1986), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n850), .A2(new_n852), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT92), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT36), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n869), .A2(new_n872), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n828), .B1(new_n873), .B2(new_n874), .ZN(G311));
  INV_X1    g450(.A(new_n873), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n869), .A2(new_n872), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n827), .B1(new_n876), .B2(new_n877), .ZN(G150));
  XNOR2_X1  g453(.A(KEYINPUT106), .B(G93), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n582), .A2(new_n879), .B1(new_n575), .B2(G55), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n505), .B(G67), .C1(new_n509), .C2(new_n510), .ZN(new_n882));
  NAND2_X1  g457(.A1(G80), .A2(G543), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n881), .B1(new_n884), .B2(G651), .ZN(new_n885));
  AOI211_X1 g460(.A(KEYINPUT105), .B(new_n515), .C1(new_n882), .C2(new_n883), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G860), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT37), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(G651), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT105), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n884), .A2(new_n881), .A3(G651), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n559), .A2(new_n893), .A3(new_n880), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n887), .A2(new_n630), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT38), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n616), .A2(new_n625), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(KEYINPUT39), .ZN(new_n900));
  INV_X1    g475(.A(G860), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n899), .B2(KEYINPUT39), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n889), .B1(new_n900), .B2(new_n902), .ZN(G145));
  XOR2_X1   g478(.A(new_n479), .B(G162), .Z(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n641), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n763), .A2(G164), .A3(new_n764), .ZN(new_n906));
  INV_X1    g481(.A(new_n764), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n500), .B1(new_n907), .B2(new_n762), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n481), .A2(G142), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n483), .A2(G130), .ZN(new_n911));
  MUX2_X1   g486(.A(G106), .B(G118), .S(G2105), .Z(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G2104), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n914), .A2(new_n645), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n645), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n858), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n855), .A2(new_n915), .A3(new_n857), .A4(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n909), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(new_n798), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n906), .A2(new_n908), .A3(new_n919), .A4(new_n918), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n921), .B2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n905), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  INV_X1    g503(.A(new_n923), .ZN(new_n929));
  INV_X1    g504(.A(new_n924), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n906), .A2(new_n908), .B1(new_n918), .B2(new_n919), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n905), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n921), .A2(new_n923), .A3(new_n924), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n927), .A2(new_n928), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g512(.A1(new_n893), .A2(new_n617), .A3(new_n880), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(G303), .A2(G305), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n829), .A2(G166), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(G290), .B(G288), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n942), .B(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT108), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n631), .B(new_n945), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(new_n896), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n896), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(new_n616), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n572), .A2(new_n583), .A3(new_n611), .A4(new_n615), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n950), .A2(KEYINPUT41), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT41), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n949), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT42), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n950), .A2(new_n951), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n947), .A2(new_n948), .A3(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n956), .B1(new_n955), .B2(new_n959), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n944), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n955), .A2(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT42), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n942), .B(new_n943), .Z(new_n965));
  NAND3_X1  g540(.A1(new_n955), .A2(new_n956), .A3(new_n959), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n939), .B1(new_n968), .B2(G868), .ZN(G295));
  AOI21_X1  g544(.A(new_n939), .B1(new_n968), .B2(G868), .ZN(G331));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT41), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n957), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n950), .A2(KEYINPUT41), .A3(new_n951), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n542), .A2(new_n543), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G651), .ZN(new_n976));
  INV_X1    g551(.A(new_n547), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n976), .A2(new_n977), .B1(new_n978), .B2(new_n528), .ZN(new_n979));
  NOR3_X1   g554(.A1(G286), .A2(new_n544), .A3(new_n547), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  AND3_X1   g556(.A1(new_n894), .A2(new_n981), .A3(new_n895), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n894), .B2(new_n895), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n973), .B(new_n974), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n894), .A2(new_n981), .A3(new_n895), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n896), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n894), .A2(new_n981), .A3(new_n895), .A4(KEYINPUT109), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n987), .A2(new_n958), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n965), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n954), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n982), .A2(new_n983), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n958), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n995), .A2(new_n944), .A3(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n998), .A3(new_n928), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  AOI22_X1  g575(.A1(new_n994), .A2(new_n954), .B1(new_n996), .B2(new_n958), .ZN(new_n1001));
  AOI21_X1  g576(.A(G37), .B1(new_n1001), .B2(new_n944), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n995), .A2(new_n997), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n965), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n971), .B1(new_n1000), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n999), .A2(new_n1005), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1002), .A2(new_n1004), .A3(KEYINPUT43), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT44), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT110), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n998), .A2(new_n928), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n944), .B1(new_n995), .B2(new_n997), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1012), .A2(KEYINPUT43), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1005), .B1(new_n1002), .B2(new_n993), .ZN(new_n1015));
  OAI21_X1  g590(.A(KEYINPUT44), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1012), .A2(new_n1005), .A3(new_n1013), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT43), .B1(new_n1002), .B2(new_n993), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n971), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT110), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1011), .A2(new_n1021), .ZN(G397));
  XNOR2_X1  g597(.A(new_n798), .B(G2067), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n500), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n471), .A2(G40), .A3(new_n474), .A4(new_n478), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT112), .ZN(new_n1031));
  INV_X1    g606(.A(G1996), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1029), .B1(new_n765), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n1032), .B2(new_n765), .ZN(new_n1034));
  OR3_X1    g609(.A1(new_n1031), .A2(KEYINPUT113), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n1031), .B2(new_n1034), .ZN(new_n1036));
  XOR2_X1   g611(.A(new_n858), .B(new_n862), .Z(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n1029), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G290), .A2(G1986), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT111), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1029), .ZN(new_n1042));
  XOR2_X1   g617(.A(new_n1042), .B(KEYINPUT48), .Z(new_n1043));
  OAI21_X1  g618(.A(new_n1029), .B1(new_n1023), .B2(new_n765), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT124), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1046), .B(KEYINPUT46), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1045), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1050));
  OAI22_X1  g625(.A1(new_n1039), .A2(new_n1043), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1052));
  INV_X1    g627(.A(new_n859), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(new_n862), .ZN(new_n1054));
  OAI22_X1  g629(.A1(new_n1052), .A2(new_n1054), .B1(G2067), .B2(new_n798), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1051), .B1(new_n1055), .B2(new_n1029), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G102), .A2(G2104), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n468), .B2(new_n497), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1058), .A2(new_n462), .B1(new_n495), .B2(new_n494), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1384), .B1(new_n1059), .B2(new_n493), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1028), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(KEYINPUT115), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1025), .A2(new_n1064), .A3(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1961), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1028), .B1(new_n1060), .B2(KEYINPUT45), .ZN(new_n1069));
  INV_X1    g644(.A(G2078), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT121), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1069), .A2(new_n1070), .A3(new_n1027), .A4(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n474), .A2(new_n478), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1074), .A2(G40), .A3(new_n471), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1024), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1027), .A2(new_n1070), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1072), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1068), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(G171), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n735), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1060), .A2(KEYINPUT45), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n824), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT116), .B(G8), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G286), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT51), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1092), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1081), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1086), .A2(G8), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1094), .B1(new_n1104), .B2(new_n1089), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1095), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1091), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT62), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1088), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1976), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1110), .B(KEYINPUT117), .C1(new_n1111), .C2(G288), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G288), .A2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1113), .B1(new_n1114), .B2(new_n1109), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1112), .B(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(G1981), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n595), .A2(new_n1117), .A3(new_n597), .A4(new_n601), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n601), .A2(new_n594), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G1981), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1118), .A2(KEYINPUT49), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT118), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT118), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1118), .A2(new_n1120), .A3(new_n1123), .A4(KEYINPUT49), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT49), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1126), .A2(new_n1109), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1125), .A2(KEYINPUT119), .A3(new_n1127), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1116), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(G8), .B1(new_n520), .B2(new_n523), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT55), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n500), .A2(new_n1061), .A3(new_n1024), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1075), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1062), .A2(KEYINPUT120), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(G2090), .ZN(new_n1143));
  INV_X1    g718(.A(G1971), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1069), .A2(new_n1027), .ZN(new_n1145));
  AOI22_X1  g720(.A1(new_n1142), .A2(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1134), .B1(new_n1146), .B2(new_n1087), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1133), .B(KEYINPUT55), .Z(new_n1148));
  INV_X1    g723(.A(KEYINPUT114), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1150), .B2(G1971), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1145), .A2(KEYINPUT114), .A3(new_n1144), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .A4(new_n1143), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1148), .A2(G8), .A3(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1147), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1103), .A2(new_n1108), .A3(new_n1132), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1116), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1086), .A2(G168), .A3(new_n1088), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1154), .A2(G8), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n1134), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1158), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(KEYINPUT63), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1147), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1160), .A2(KEYINPUT63), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1155), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1132), .ZN(new_n1168));
  OR2_X1    g743(.A1(G288), .A2(G1976), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1169), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1118), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1110), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1157), .A2(new_n1164), .A3(new_n1168), .A4(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(G2067), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1066), .A2(new_n778), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1176), .A2(new_n616), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1178));
  INV_X1    g753(.A(G1956), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT56), .B(G2072), .Z(new_n1181));
  INV_X1    g756(.A(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1069), .A2(new_n1027), .A3(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT57), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n572), .A2(new_n1184), .A3(new_n583), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1178), .A2(new_n1180), .A3(new_n1183), .A4(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1177), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1178), .A2(new_n1185), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1186), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1176), .A2(new_n1195), .A3(new_n624), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1083), .A2(new_n1084), .A3(G1996), .ZN(new_n1197));
  XNOR2_X1  g772(.A(KEYINPUT58), .B(G1341), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1175), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n559), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT59), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1202), .B(new_n559), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1190), .A2(KEYINPUT61), .A3(new_n1186), .ZN(new_n1205));
  AND4_X1   g780(.A1(new_n1194), .A2(new_n1196), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  AND2_X1   g781(.A1(new_n1176), .A2(new_n616), .ZN(new_n1207));
  OAI21_X1  g782(.A(KEYINPUT60), .B1(new_n1207), .B2(new_n1177), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1191), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1132), .A2(new_n1156), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1027), .A2(new_n1211), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1077), .A2(new_n1212), .A3(KEYINPUT53), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1077), .B1(KEYINPUT53), .B2(new_n1212), .ZN(new_n1214));
  OAI211_X1 g789(.A(G301), .B(new_n1068), .C1(new_n1213), .C2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1081), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT54), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g793(.A1(new_n1068), .A2(G301), .A3(new_n1079), .A4(new_n1073), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1150), .B(new_n1070), .C1(new_n1211), .C2(new_n1071), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1077), .A2(new_n1212), .A3(KEYINPUT53), .ZN(new_n1221));
  AOI22_X1  g796(.A1(new_n1220), .A2(new_n1221), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1222));
  OAI211_X1 g797(.A(KEYINPUT54), .B(new_n1219), .C1(new_n1222), .C2(G301), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1218), .A2(new_n1107), .A3(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1210), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n1226));
  AOI21_X1  g801(.A(new_n1209), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g802(.A(KEYINPUT123), .B1(new_n1210), .B2(new_n1224), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1173), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1041), .B1(G1986), .B2(G290), .ZN(new_n1230));
  NOR3_X1   g805(.A1(new_n1230), .A2(new_n1028), .A3(new_n1027), .ZN(new_n1231));
  OR2_X1    g806(.A1(new_n1039), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1056), .B1(new_n1229), .B2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  OAI211_X1 g808(.A(new_n680), .B(G319), .C1(new_n726), .C2(new_n727), .ZN(new_n1235));
  OAI21_X1  g809(.A(KEYINPUT126), .B1(new_n1235), .B2(G227), .ZN(new_n1236));
  INV_X1    g810(.A(G227), .ZN(new_n1237));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n1238));
  INV_X1    g812(.A(G14), .ZN(new_n1239));
  AOI21_X1  g813(.A(new_n1239), .B1(new_n668), .B2(new_n677), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n460), .B1(new_n1240), .B2(new_n679), .ZN(new_n1241));
  NAND4_X1  g815(.A1(new_n1237), .A2(new_n728), .A3(new_n1238), .A4(new_n1241), .ZN(new_n1242));
  AND2_X1   g816(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g817(.A1(new_n1008), .A2(new_n1243), .A3(new_n936), .A4(new_n1009), .ZN(new_n1244));
  XNOR2_X1  g818(.A(new_n1244), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1246));
  XNOR2_X1  g820(.A(new_n1244), .B(new_n1246), .ZN(G225));
endmodule


