

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(G2104), .B(KEYINPUT66), .ZN(n526) );
  XNOR2_X2 U550 ( .A(n617), .B(KEYINPUT64), .ZN(n662) );
  NAND2_X1 U551 ( .A1(n663), .A2(G8), .ZN(n709) );
  XNOR2_X1 U552 ( .A(n554), .B(KEYINPUT94), .ZN(G164) );
  INV_X1 U553 ( .A(KEYINPUT102), .ZN(n632) );
  AND2_X1 U554 ( .A1(n526), .A2(n525), .ZN(n549) );
  NOR2_X1 U555 ( .A1(n526), .A2(n525), .ZN(n544) );
  NOR2_X1 U556 ( .A1(n645), .A2(n975), .ZN(n633) );
  XNOR2_X1 U557 ( .A(n651), .B(n650), .ZN(n655) );
  INV_X1 U558 ( .A(KEYINPUT103), .ZN(n650) );
  NOR2_X1 U559 ( .A1(n592), .A2(n536), .ZN(n807) );
  NOR2_X1 U560 ( .A1(G651), .A2(n592), .ZN(n802) );
  XNOR2_X1 U561 ( .A(n524), .B(n523), .ZN(n528) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n523) );
  AND2_X1 U563 ( .A1(n533), .A2(n532), .ZN(n517) );
  XOR2_X1 U564 ( .A(n752), .B(KEYINPUT98), .Z(n518) );
  XOR2_X1 U565 ( .A(n766), .B(KEYINPUT113), .Z(n519) );
  AND2_X1 U566 ( .A1(n518), .A2(n753), .ZN(n520) );
  NOR2_X1 U567 ( .A1(n690), .A2(n689), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n687), .A2(n686), .ZN(n522) );
  XNOR2_X1 U569 ( .A(n618), .B(KEYINPUT65), .ZN(n619) );
  NOR2_X1 U570 ( .A1(n978), .A2(n621), .ZN(n623) );
  BUF_X1 U571 ( .A(n636), .Z(n657) );
  NOR2_X1 U572 ( .A1(n670), .A2(n669), .ZN(n671) );
  BUF_X1 U573 ( .A(n662), .Z(n663) );
  NOR2_X1 U574 ( .A1(G164), .A2(G1384), .ZN(n740) );
  XNOR2_X1 U575 ( .A(KEYINPUT13), .B(KEYINPUT78), .ZN(n610) );
  INV_X1 U576 ( .A(KEYINPUT17), .ZN(n530) );
  XNOR2_X1 U577 ( .A(KEYINPUT15), .B(n631), .ZN(n975) );
  XNOR2_X1 U578 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U579 ( .A1(n903), .A2(G138), .ZN(n550) );
  XOR2_X1 U580 ( .A(KEYINPUT1), .B(n535), .Z(n803) );
  NOR2_X1 U581 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U582 ( .A1(n553), .A2(n552), .ZN(n554) );
  INV_X1 U583 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n549), .A2(G101), .ZN(n524) );
  BUF_X2 U585 ( .A(n544), .Z(n908) );
  NAND2_X1 U586 ( .A1(n908), .A2(G125), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U588 ( .A(n529), .B(KEYINPUT67), .ZN(n534) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n907) );
  NAND2_X1 U590 ( .A1(G113), .A2(n907), .ZN(n533) );
  NOR2_X1 U591 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XNOR2_X2 U592 ( .A(n531), .B(n530), .ZN(n903) );
  NAND2_X1 U593 ( .A1(G137), .A2(n903), .ZN(n532) );
  AND2_X2 U594 ( .A1(n534), .A2(n517), .ZN(G160) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(G651), .Z(n536) );
  NOR2_X1 U596 ( .A1(G543), .A2(n536), .ZN(n535) );
  NAND2_X1 U597 ( .A1(G65), .A2(n803), .ZN(n538) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n592) );
  NAND2_X1 U599 ( .A1(G78), .A2(n807), .ZN(n537) );
  NAND2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n541) );
  NOR2_X1 U601 ( .A1(G651), .A2(G543), .ZN(n806) );
  NAND2_X1 U602 ( .A1(G91), .A2(n806), .ZN(n539) );
  XNOR2_X1 U603 ( .A(KEYINPUT71), .B(n539), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n802), .A2(G53), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(G299) );
  NAND2_X1 U607 ( .A1(G126), .A2(n544), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G114), .A2(n907), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n548) );
  INV_X1 U610 ( .A(KEYINPUT93), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(n553) );
  BUF_X2 U612 ( .A(n549), .Z(n904) );
  NAND2_X1 U613 ( .A1(n904), .A2(G102), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U615 ( .A1(G90), .A2(n806), .ZN(n556) );
  NAND2_X1 U616 ( .A1(G77), .A2(n807), .ZN(n555) );
  NAND2_X1 U617 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U618 ( .A(n557), .B(KEYINPUT9), .ZN(n559) );
  NAND2_X1 U619 ( .A1(G52), .A2(n802), .ZN(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U621 ( .A1(G64), .A2(n803), .ZN(n560) );
  XNOR2_X1 U622 ( .A(KEYINPUT69), .B(n560), .ZN(n561) );
  NOR2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(KEYINPUT70), .B(n563), .ZN(G171) );
  NAND2_X1 U625 ( .A1(G63), .A2(n803), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT84), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G51), .A2(n802), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(KEYINPUT85), .Z(n567) );
  XNOR2_X1 U630 ( .A(n568), .B(n567), .ZN(n577) );
  NAND2_X1 U631 ( .A1(G76), .A2(n807), .ZN(n569) );
  XNOR2_X1 U632 ( .A(KEYINPUT82), .B(n569), .ZN(n573) );
  XOR2_X1 U633 ( .A(KEYINPUT4), .B(KEYINPUT81), .Z(n571) );
  NAND2_X1 U634 ( .A1(G89), .A2(n806), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U637 ( .A(n574), .B(KEYINPUT83), .ZN(n575) );
  XNOR2_X1 U638 ( .A(KEYINPUT5), .B(n575), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT7), .B(n578), .Z(G168) );
  NAND2_X1 U640 ( .A1(G88), .A2(n806), .ZN(n580) );
  NAND2_X1 U641 ( .A1(G75), .A2(n807), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U643 ( .A1(n802), .A2(G50), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G62), .A2(n803), .ZN(n581) );
  NAND2_X1 U645 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U646 ( .A1(n584), .A2(n583), .ZN(G166) );
  INV_X1 U647 ( .A(G166), .ZN(G303) );
  XOR2_X1 U648 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U649 ( .A1(G86), .A2(n806), .ZN(n586) );
  NAND2_X1 U650 ( .A1(G48), .A2(n802), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U652 ( .A1(n807), .A2(G73), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT2), .B(n587), .Z(n588) );
  NOR2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G61), .A2(n803), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(G305) );
  NAND2_X1 U657 ( .A1(G87), .A2(n592), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G74), .A2(G651), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U660 ( .A1(n803), .A2(n595), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n802), .A2(G49), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n597), .A2(n596), .ZN(G288) );
  NAND2_X1 U663 ( .A1(n806), .A2(G85), .ZN(n599) );
  NAND2_X1 U664 ( .A1(G60), .A2(n803), .ZN(n598) );
  NAND2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U666 ( .A1(n802), .A2(G47), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G72), .A2(n807), .ZN(n600) );
  NAND2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U669 ( .A1(n603), .A2(n602), .ZN(G290) );
  XOR2_X1 U670 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n605) );
  NAND2_X1 U671 ( .A1(G56), .A2(n803), .ZN(n604) );
  XNOR2_X1 U672 ( .A(n605), .B(n604), .ZN(n613) );
  NAND2_X1 U673 ( .A1(G68), .A2(n807), .ZN(n606) );
  XNOR2_X1 U674 ( .A(KEYINPUT77), .B(n606), .ZN(n609) );
  NAND2_X1 U675 ( .A1(n806), .A2(G81), .ZN(n607) );
  XOR2_X1 U676 ( .A(n607), .B(KEYINPUT12), .Z(n608) );
  NOR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n611) );
  NOR2_X1 U678 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n802), .A2(G43), .ZN(n614) );
  NAND2_X1 U680 ( .A1(n615), .A2(n614), .ZN(n978) );
  NAND2_X1 U681 ( .A1(G160), .A2(G40), .ZN(n739) );
  INV_X1 U682 ( .A(n739), .ZN(n616) );
  NAND2_X1 U683 ( .A1(n616), .A2(n740), .ZN(n617) );
  INV_X2 U684 ( .A(n662), .ZN(n636) );
  NAND2_X1 U685 ( .A1(G1996), .A2(n636), .ZN(n620) );
  XOR2_X1 U686 ( .A(KEYINPUT26), .B(KEYINPUT101), .Z(n618) );
  XNOR2_X1 U687 ( .A(n620), .B(n619), .ZN(n621) );
  INV_X1 U688 ( .A(n636), .ZN(n674) );
  NAND2_X1 U689 ( .A1(n674), .A2(G1341), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n623), .A2(n622), .ZN(n645) );
  NAND2_X1 U691 ( .A1(n806), .A2(G92), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G66), .A2(n803), .ZN(n624) );
  NAND2_X1 U693 ( .A1(n625), .A2(n624), .ZN(n630) );
  NAND2_X1 U694 ( .A1(n802), .A2(G54), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G79), .A2(n807), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U697 ( .A(KEYINPUT79), .B(n628), .Z(n629) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n633), .B(n632), .ZN(n643) );
  NOR2_X1 U700 ( .A1(G2067), .A2(n674), .ZN(n635) );
  NOR2_X1 U701 ( .A1(G1348), .A2(n657), .ZN(n634) );
  NOR2_X1 U702 ( .A1(n635), .A2(n634), .ZN(n641) );
  NAND2_X1 U703 ( .A1(n636), .A2(G2072), .ZN(n638) );
  XNOR2_X1 U704 ( .A(KEYINPUT100), .B(KEYINPUT27), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n638), .B(n637), .ZN(n640) );
  INV_X1 U706 ( .A(G1956), .ZN(n981) );
  NOR2_X1 U707 ( .A1(n657), .A2(n981), .ZN(n639) );
  OR2_X2 U708 ( .A1(n640), .A2(n639), .ZN(n652) );
  OR2_X2 U709 ( .A1(G299), .A2(n652), .ZN(n644) );
  AND2_X1 U710 ( .A1(n641), .A2(n644), .ZN(n642) );
  NAND2_X1 U711 ( .A1(n643), .A2(n642), .ZN(n649) );
  INV_X1 U712 ( .A(n644), .ZN(n647) );
  NAND2_X1 U713 ( .A1(n975), .A2(n645), .ZN(n646) );
  OR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U715 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U716 ( .A1(G299), .A2(n652), .ZN(n653) );
  XOR2_X1 U717 ( .A(KEYINPUT28), .B(n653), .Z(n654) );
  NOR2_X2 U718 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U719 ( .A(n656), .B(KEYINPUT29), .ZN(n661) );
  XNOR2_X1 U720 ( .A(G1961), .B(KEYINPUT99), .ZN(n1001) );
  NOR2_X1 U721 ( .A1(n657), .A2(n1001), .ZN(n659) );
  XNOR2_X1 U722 ( .A(G2078), .B(KEYINPUT25), .ZN(n961) );
  NOR2_X1 U723 ( .A1(n674), .A2(n961), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n667) );
  NAND2_X1 U725 ( .A1(G171), .A2(n667), .ZN(n660) );
  NAND2_X1 U726 ( .A1(n661), .A2(n660), .ZN(n686) );
  NOR2_X1 U727 ( .A1(G1966), .A2(n709), .ZN(n689) );
  NOR2_X1 U728 ( .A1(n674), .A2(G2084), .ZN(n688) );
  NOR2_X1 U729 ( .A1(n689), .A2(n688), .ZN(n664) );
  NAND2_X1 U730 ( .A1(G8), .A2(n664), .ZN(n665) );
  XNOR2_X1 U731 ( .A(KEYINPUT30), .B(n665), .ZN(n666) );
  NOR2_X1 U732 ( .A1(n666), .A2(G168), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n667), .A2(G171), .ZN(n668) );
  XNOR2_X1 U734 ( .A(n668), .B(KEYINPUT104), .ZN(n669) );
  XNOR2_X1 U735 ( .A(n671), .B(KEYINPUT105), .ZN(n672) );
  XNOR2_X1 U736 ( .A(n672), .B(KEYINPUT31), .ZN(n687) );
  INV_X1 U737 ( .A(G8), .ZN(n679) );
  NOR2_X1 U738 ( .A1(G1971), .A2(n709), .ZN(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT106), .ZN(n676) );
  NOR2_X1 U740 ( .A1(n674), .A2(G2090), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n677), .A2(G303), .ZN(n678) );
  OR2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n681) );
  AND2_X1 U744 ( .A1(n687), .A2(n681), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n686), .A2(n680), .ZN(n684) );
  INV_X1 U746 ( .A(n681), .ZN(n682) );
  OR2_X1 U747 ( .A1(n682), .A2(G286), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U749 ( .A(n685), .B(KEYINPUT32), .ZN(n692) );
  AND2_X1 U750 ( .A1(G8), .A2(n688), .ZN(n690) );
  NAND2_X1 U751 ( .A1(n522), .A2(n521), .ZN(n691) );
  NAND2_X1 U752 ( .A1(n692), .A2(n691), .ZN(n694) );
  INV_X1 U753 ( .A(KEYINPUT107), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n694), .B(n693), .ZN(n705) );
  NOR2_X1 U755 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U756 ( .A1(G8), .A2(n695), .ZN(n696) );
  NAND2_X1 U757 ( .A1(n705), .A2(n696), .ZN(n697) );
  XNOR2_X1 U758 ( .A(n697), .B(KEYINPUT110), .ZN(n698) );
  AND2_X2 U759 ( .A1(n698), .A2(n709), .ZN(n720) );
  NOR2_X1 U760 ( .A1(G1981), .A2(G305), .ZN(n699) );
  XOR2_X1 U761 ( .A(n699), .B(KEYINPUT24), .Z(n700) );
  OR2_X1 U762 ( .A1(n709), .A2(n700), .ZN(n718) );
  NOR2_X1 U763 ( .A1(G1976), .A2(G288), .ZN(n708) );
  NOR2_X1 U764 ( .A1(G1971), .A2(G303), .ZN(n701) );
  NOR2_X1 U765 ( .A1(n708), .A2(n701), .ZN(n985) );
  XNOR2_X1 U766 ( .A(KEYINPUT108), .B(n985), .ZN(n703) );
  INV_X1 U767 ( .A(KEYINPUT33), .ZN(n702) );
  AND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n714) );
  INV_X1 U770 ( .A(n709), .ZN(n706) );
  NAND2_X1 U771 ( .A1(G1976), .A2(G288), .ZN(n984) );
  AND2_X1 U772 ( .A1(n706), .A2(n984), .ZN(n707) );
  NOR2_X1 U773 ( .A1(KEYINPUT33), .A2(n707), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n708), .A2(KEYINPUT33), .ZN(n710) );
  NOR2_X1 U775 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  AND2_X1 U777 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U778 ( .A(G1981), .B(KEYINPUT109), .ZN(n715) );
  XNOR2_X1 U779 ( .A(n715), .B(G305), .ZN(n991) );
  NAND2_X1 U780 ( .A1(n716), .A2(n991), .ZN(n717) );
  NAND2_X1 U781 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X2 U782 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U783 ( .A(n721), .B(KEYINPUT111), .ZN(n754) );
  NAND2_X1 U784 ( .A1(G107), .A2(n907), .ZN(n723) );
  NAND2_X1 U785 ( .A1(G131), .A2(n903), .ZN(n722) );
  NAND2_X1 U786 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U787 ( .A1(G119), .A2(n908), .ZN(n725) );
  NAND2_X1 U788 ( .A1(G95), .A2(n904), .ZN(n724) );
  NAND2_X1 U789 ( .A1(n725), .A2(n724), .ZN(n726) );
  OR2_X1 U790 ( .A1(n727), .A2(n726), .ZN(n895) );
  NAND2_X1 U791 ( .A1(G1991), .A2(n895), .ZN(n728) );
  XNOR2_X1 U792 ( .A(n728), .B(KEYINPUT96), .ZN(n738) );
  NAND2_X1 U793 ( .A1(G105), .A2(n904), .ZN(n729) );
  XNOR2_X1 U794 ( .A(n729), .B(KEYINPUT38), .ZN(n736) );
  NAND2_X1 U795 ( .A1(G117), .A2(n907), .ZN(n731) );
  NAND2_X1 U796 ( .A1(G129), .A2(n908), .ZN(n730) );
  NAND2_X1 U797 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U798 ( .A1(G141), .A2(n903), .ZN(n732) );
  XNOR2_X1 U799 ( .A(KEYINPUT97), .B(n732), .ZN(n733) );
  NOR2_X1 U800 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U801 ( .A1(n736), .A2(n735), .ZN(n915) );
  NAND2_X1 U802 ( .A1(G1996), .A2(n915), .ZN(n737) );
  NAND2_X1 U803 ( .A1(n738), .A2(n737), .ZN(n941) );
  NOR2_X1 U804 ( .A1(n740), .A2(n739), .ZN(n765) );
  NAND2_X1 U805 ( .A1(n941), .A2(n765), .ZN(n751) );
  NAND2_X1 U806 ( .A1(G140), .A2(n903), .ZN(n742) );
  NAND2_X1 U807 ( .A1(G104), .A2(n904), .ZN(n741) );
  NAND2_X1 U808 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U809 ( .A(KEYINPUT34), .B(n743), .ZN(n748) );
  NAND2_X1 U810 ( .A1(G116), .A2(n907), .ZN(n745) );
  NAND2_X1 U811 ( .A1(G128), .A2(n908), .ZN(n744) );
  NAND2_X1 U812 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U813 ( .A(KEYINPUT35), .B(n746), .Z(n747) );
  NOR2_X1 U814 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n749), .ZN(n899) );
  XNOR2_X1 U816 ( .A(G2067), .B(KEYINPUT37), .ZN(n762) );
  NOR2_X1 U817 ( .A1(n899), .A2(n762), .ZN(n936) );
  NAND2_X1 U818 ( .A1(n936), .A2(n765), .ZN(n750) );
  XOR2_X1 U819 ( .A(KEYINPUT95), .B(n750), .Z(n760) );
  NAND2_X1 U820 ( .A1(n751), .A2(n760), .ZN(n752) );
  XNOR2_X1 U821 ( .A(G1986), .B(G290), .ZN(n980) );
  NAND2_X1 U822 ( .A1(n765), .A2(n980), .ZN(n753) );
  NAND2_X1 U823 ( .A1(n754), .A2(n520), .ZN(n767) );
  NOR2_X1 U824 ( .A1(n915), .A2(G1996), .ZN(n755) );
  XNOR2_X1 U825 ( .A(n755), .B(KEYINPUT112), .ZN(n934) );
  NOR2_X1 U826 ( .A1(G1991), .A2(n895), .ZN(n942) );
  NOR2_X1 U827 ( .A1(G1986), .A2(G290), .ZN(n756) );
  NOR2_X1 U828 ( .A1(n942), .A2(n756), .ZN(n757) );
  NOR2_X1 U829 ( .A1(n941), .A2(n757), .ZN(n758) );
  NOR2_X1 U830 ( .A1(n934), .A2(n758), .ZN(n759) );
  XNOR2_X1 U831 ( .A(KEYINPUT39), .B(n759), .ZN(n761) );
  NAND2_X1 U832 ( .A1(n761), .A2(n760), .ZN(n763) );
  NAND2_X1 U833 ( .A1(n899), .A2(n762), .ZN(n937) );
  NAND2_X1 U834 ( .A1(n763), .A2(n937), .ZN(n764) );
  NAND2_X1 U835 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U836 ( .A1(n767), .A2(n519), .ZN(n768) );
  XNOR2_X1 U837 ( .A(n768), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U838 ( .A(G171), .ZN(G301) );
  XOR2_X1 U839 ( .A(G2443), .B(G2446), .Z(n770) );
  XNOR2_X1 U840 ( .A(G2427), .B(G2451), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n770), .B(n769), .ZN(n776) );
  XOR2_X1 U842 ( .A(G2430), .B(G2454), .Z(n772) );
  XNOR2_X1 U843 ( .A(G1348), .B(G1341), .ZN(n771) );
  XNOR2_X1 U844 ( .A(n772), .B(n771), .ZN(n774) );
  XOR2_X1 U845 ( .A(G2435), .B(G2438), .Z(n773) );
  XNOR2_X1 U846 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U847 ( .A(n776), .B(n775), .Z(n777) );
  AND2_X1 U848 ( .A1(G14), .A2(n777), .ZN(G401) );
  AND2_X1 U849 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U850 ( .A(G132), .ZN(G219) );
  INV_X1 U851 ( .A(G82), .ZN(G220) );
  NAND2_X1 U852 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U853 ( .A(n778), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U854 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n780) );
  XNOR2_X1 U855 ( .A(G223), .B(KEYINPUT73), .ZN(n845) );
  NAND2_X1 U856 ( .A1(G567), .A2(n845), .ZN(n779) );
  XNOR2_X1 U857 ( .A(n780), .B(n779), .ZN(n781) );
  XOR2_X1 U858 ( .A(KEYINPUT11), .B(n781), .Z(G234) );
  INV_X1 U859 ( .A(G860), .ZN(n815) );
  OR2_X1 U860 ( .A1(n978), .A2(n815), .ZN(G153) );
  NOR2_X1 U861 ( .A1(G868), .A2(n975), .ZN(n783) );
  INV_X1 U862 ( .A(G868), .ZN(n827) );
  NOR2_X1 U863 ( .A1(G301), .A2(n827), .ZN(n782) );
  NOR2_X1 U864 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U865 ( .A(KEYINPUT80), .B(n784), .ZN(G284) );
  NOR2_X1 U866 ( .A1(G286), .A2(n827), .ZN(n786) );
  NOR2_X1 U867 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U868 ( .A1(n786), .A2(n785), .ZN(G297) );
  NAND2_X1 U869 ( .A1(n815), .A2(G559), .ZN(n787) );
  INV_X1 U870 ( .A(n975), .ZN(n812) );
  NAND2_X1 U871 ( .A1(n787), .A2(n812), .ZN(n788) );
  XNOR2_X1 U872 ( .A(n788), .B(KEYINPUT86), .ZN(n789) );
  XNOR2_X1 U873 ( .A(KEYINPUT16), .B(n789), .ZN(G148) );
  NOR2_X1 U874 ( .A1(G868), .A2(n978), .ZN(n792) );
  NAND2_X1 U875 ( .A1(G868), .A2(n812), .ZN(n790) );
  NOR2_X1 U876 ( .A1(G559), .A2(n790), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G282) );
  NAND2_X1 U878 ( .A1(G111), .A2(n907), .ZN(n794) );
  NAND2_X1 U879 ( .A1(G135), .A2(n903), .ZN(n793) );
  NAND2_X1 U880 ( .A1(n794), .A2(n793), .ZN(n799) );
  NAND2_X1 U881 ( .A1(n908), .A2(G123), .ZN(n795) );
  XNOR2_X1 U882 ( .A(n795), .B(KEYINPUT18), .ZN(n797) );
  NAND2_X1 U883 ( .A1(G99), .A2(n904), .ZN(n796) );
  NAND2_X1 U884 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n940) );
  XNOR2_X1 U886 ( .A(G2096), .B(n940), .ZN(n801) );
  INV_X1 U887 ( .A(G2100), .ZN(n800) );
  NAND2_X1 U888 ( .A1(n801), .A2(n800), .ZN(G156) );
  NAND2_X1 U889 ( .A1(n802), .A2(G55), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G67), .A2(n803), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G93), .A2(n806), .ZN(n809) );
  NAND2_X1 U893 ( .A1(G80), .A2(n807), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n809), .A2(n808), .ZN(n810) );
  OR2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n828) );
  XNOR2_X1 U896 ( .A(n828), .B(KEYINPUT88), .ZN(n817) );
  XNOR2_X1 U897 ( .A(n978), .B(KEYINPUT87), .ZN(n814) );
  NAND2_X1 U898 ( .A1(n812), .A2(G559), .ZN(n813) );
  XNOR2_X1 U899 ( .A(n814), .B(n813), .ZN(n824) );
  NAND2_X1 U900 ( .A1(n824), .A2(n815), .ZN(n816) );
  XNOR2_X1 U901 ( .A(n817), .B(n816), .ZN(G145) );
  XOR2_X1 U902 ( .A(KEYINPUT89), .B(KEYINPUT19), .Z(n818) );
  XNOR2_X1 U903 ( .A(G288), .B(n818), .ZN(n819) );
  XNOR2_X1 U904 ( .A(G166), .B(n819), .ZN(n821) );
  XOR2_X1 U905 ( .A(G290), .B(G299), .Z(n820) );
  XNOR2_X1 U906 ( .A(n821), .B(n820), .ZN(n822) );
  XNOR2_X1 U907 ( .A(n828), .B(n822), .ZN(n823) );
  XNOR2_X1 U908 ( .A(G305), .B(n823), .ZN(n870) );
  XNOR2_X1 U909 ( .A(n870), .B(n824), .ZN(n825) );
  NAND2_X1 U910 ( .A1(n825), .A2(G868), .ZN(n826) );
  XNOR2_X1 U911 ( .A(n826), .B(KEYINPUT90), .ZN(n830) );
  NAND2_X1 U912 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U913 ( .A1(n830), .A2(n829), .ZN(G295) );
  NAND2_X1 U914 ( .A1(G2078), .A2(G2084), .ZN(n831) );
  XOR2_X1 U915 ( .A(KEYINPUT20), .B(n831), .Z(n832) );
  NAND2_X1 U916 ( .A1(G2090), .A2(n832), .ZN(n834) );
  XOR2_X1 U917 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n833) );
  XNOR2_X1 U918 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U919 ( .A1(G2072), .A2(n835), .ZN(G158) );
  XOR2_X1 U920 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U921 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U922 ( .A1(G108), .A2(G120), .ZN(n836) );
  NOR2_X1 U923 ( .A1(G237), .A2(n836), .ZN(n837) );
  NAND2_X1 U924 ( .A1(G69), .A2(n837), .ZN(n850) );
  NAND2_X1 U925 ( .A1(n850), .A2(G567), .ZN(n843) );
  NOR2_X1 U926 ( .A1(G220), .A2(G219), .ZN(n838) );
  XOR2_X1 U927 ( .A(KEYINPUT22), .B(n838), .Z(n839) );
  NOR2_X1 U928 ( .A1(G218), .A2(n839), .ZN(n840) );
  NAND2_X1 U929 ( .A1(G96), .A2(n840), .ZN(n849) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n849), .ZN(n841) );
  XNOR2_X1 U931 ( .A(KEYINPUT92), .B(n841), .ZN(n842) );
  NAND2_X1 U932 ( .A1(n843), .A2(n842), .ZN(n851) );
  NAND2_X1 U933 ( .A1(G483), .A2(G661), .ZN(n844) );
  NOR2_X1 U934 ( .A1(n851), .A2(n844), .ZN(n848) );
  NAND2_X1 U935 ( .A1(n848), .A2(G36), .ZN(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n845), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n846) );
  NAND2_X1 U938 ( .A1(G661), .A2(n846), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n847) );
  NAND2_X1 U940 ( .A1(n848), .A2(n847), .ZN(G188) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G108), .ZN(G238) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  INV_X1 U948 ( .A(n851), .ZN(G319) );
  XOR2_X1 U949 ( .A(G2096), .B(KEYINPUT114), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2067), .B(KEYINPUT43), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n854), .B(KEYINPUT42), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2072), .B(G2090), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G2678), .B(G2100), .Z(n858) );
  XNOR2_X1 U956 ( .A(G2078), .B(G2084), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U959 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1956), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n863), .B(G2474), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U965 ( .A(KEYINPUT41), .B(G1981), .Z(n867) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1961), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(G229) );
  XNOR2_X1 U969 ( .A(n870), .B(KEYINPUT121), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n978), .B(G286), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n874) );
  XOR2_X1 U972 ( .A(n975), .B(G301), .Z(n873) );
  XNOR2_X1 U973 ( .A(n874), .B(n873), .ZN(n875) );
  NOR2_X1 U974 ( .A1(G37), .A2(n875), .ZN(G397) );
  NAND2_X1 U975 ( .A1(G112), .A2(n907), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G136), .A2(n903), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G124), .A2(n908), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT115), .B(n878), .Z(n879) );
  XNOR2_X1 U980 ( .A(n879), .B(KEYINPUT44), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G100), .A2(n904), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U984 ( .A1(G118), .A2(n907), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G130), .A2(n908), .ZN(n884) );
  NAND2_X1 U986 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G142), .A2(n903), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G106), .A2(n904), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n888), .Z(n889) );
  XNOR2_X1 U991 ( .A(KEYINPUT116), .B(n889), .ZN(n890) );
  NOR2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n902) );
  XOR2_X1 U993 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n893) );
  XNOR2_X1 U994 ( .A(KEYINPUT119), .B(KEYINPUT118), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n940), .B(n894), .ZN(n897) );
  XNOR2_X1 U997 ( .A(n895), .B(G162), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U999 ( .A(G164), .B(n898), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n917) );
  NAND2_X1 U1002 ( .A1(G139), .A2(n903), .ZN(n906) );
  NAND2_X1 U1003 ( .A1(G103), .A2(n904), .ZN(n905) );
  NAND2_X1 U1004 ( .A1(n906), .A2(n905), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(G115), .A2(n907), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(G127), .A2(n908), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n911), .Z(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1010 ( .A(KEYINPUT117), .B(n914), .Z(n928) );
  XNOR2_X1 U1011 ( .A(n915), .B(n928), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(G160), .B(n918), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G37), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(KEYINPUT120), .B(n920), .ZN(G395) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n921) );
  XOR2_X1 U1017 ( .A(KEYINPUT49), .B(n921), .Z(n922) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n923), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(KEYINPUT122), .B(n924), .ZN(n926) );
  NOR2_X1 U1021 ( .A1(G397), .A2(G395), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT123), .B(n927), .Z(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1025 ( .A(G164), .B(G2078), .ZN(n931) );
  XNOR2_X1 U1026 ( .A(G2072), .B(n928), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT124), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n932), .B(KEYINPUT50), .ZN(n950) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n935), .Z(n948) );
  INV_X1 U1033 ( .A(n936), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(n937), .ZN(n946) );
  XOR2_X1 U1035 ( .A(G160), .B(G2084), .Z(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  NOR2_X1 U1041 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(n951), .ZN(n952) );
  INV_X1 U1043 ( .A(KEYINPUT55), .ZN(n971) );
  NAND2_X1 U1044 ( .A1(n952), .A2(n971), .ZN(n953) );
  NAND2_X1 U1045 ( .A1(n953), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n966) );
  XNOR2_X1 U1047 ( .A(G2067), .B(G26), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(n955), .A2(n954), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G1991), .B(G25), .Z(n956) );
  NAND2_X1 U1051 ( .A1(n956), .A2(G28), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G32), .B(G1996), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1055 ( .A(G27), .B(n961), .Z(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n964), .ZN(n965) );
  NOR2_X1 U1058 ( .A1(n966), .A2(n965), .ZN(n969) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n967), .ZN(n968) );
  NAND2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n971), .B(n970), .ZN(n973) );
  INV_X1 U1063 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n974), .ZN(n1028) );
  XNOR2_X1 U1066 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1067 ( .A(G1348), .B(n975), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G301), .B(G1961), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n998) );
  XNOR2_X1 U1070 ( .A(G1341), .B(n978), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n990) );
  XNOR2_X1 U1072 ( .A(G299), .B(n981), .ZN(n983) );
  NAND2_X1 U1073 ( .A1(G1971), .A2(G303), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n987) );
  NAND2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(n988), .B(KEYINPUT126), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n996) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n993), .B(KEYINPUT125), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(n994), .B(KEYINPUT57), .ZN(n995) );
  NOR2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  INV_X1 U1086 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1087 ( .A(G5), .B(n1001), .ZN(n1014) );
  XNOR2_X1 U1088 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1089 ( .A(n1002), .B(G4), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(G20), .B(G1956), .ZN(n1003) );
  NOR2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1094 ( .A(KEYINPUT127), .B(G1981), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G6), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1010), .Z(n1012) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(G1986), .B(G24), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(G1971), .B(G22), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(G1976), .B(G23), .Z(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1111 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1112 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

