//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n584, new_n585, new_n586,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n599, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n636, new_n639,
    new_n641, new_n642, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OR3_X1    g037(.A1(new_n462), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n462), .B2(G2104), .ZN(new_n465));
  OAI211_X1 g040(.A(new_n463), .B(G137), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n462), .A2(G2104), .ZN(new_n473));
  AND2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n470), .B1(new_n474), .B2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n473), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n476), .A2(KEYINPUT65), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n469), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n468), .B1(new_n479), .B2(G2105), .ZN(G160));
  OAI21_X1  g055(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(KEYINPUT67), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n463), .B(new_n483), .C1(new_n464), .C2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT68), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT68), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n488), .A3(G2105), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n493), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT69), .Z(new_n495));
  NAND2_X1  g070(.A1(new_n485), .A2(new_n493), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G136), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n491), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G162));
  NOR2_X1   g075(.A1(new_n493), .A2(G114), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT70), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n505), .B1(new_n501), .B2(new_n502), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n493), .A2(KEYINPUT4), .A3(G138), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n463), .B(new_n508), .C1(new_n464), .C2(new_n465), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n472), .A2(new_n473), .A3(G138), .A4(new_n493), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(G126), .A2(G2105), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n463), .B(new_n513), .C1(new_n464), .C2(new_n465), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n507), .A2(new_n509), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(KEYINPUT72), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n517), .B(G543), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(KEYINPUT72), .B1(new_n523), .B2(G543), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT6), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT6), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(G543), .B1(new_n518), .B2(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(new_n527), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n535), .B1(new_n538), .B2(new_n520), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n521), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n539), .A2(G88), .B1(G50), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  AND2_X1   g118(.A1(new_n532), .A2(new_n534), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n528), .A2(G89), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n540), .A2(G51), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n547));
  NAND3_X1  g122(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n545), .A2(new_n546), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n520), .B(new_n552), .C1(new_n526), .C2(new_n527), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n552), .B1(new_n538), .B2(new_n520), .ZN(new_n555));
  OAI211_X1 g130(.A(G63), .B(G651), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(G168));
  OAI21_X1  g133(.A(G64), .B1(new_n554), .B2(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(G77), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(G90), .ZN(new_n562));
  AOI211_X1 g137(.A(new_n535), .B(new_n562), .C1(new_n538), .C2(new_n520), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n540), .A2(G52), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT76), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n562), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n528), .A2(new_n544), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n568), .A2(new_n569), .A3(new_n564), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n561), .A2(G651), .B1(new_n566), .B2(new_n570), .ZN(G171));
  INV_X1    g146(.A(G56), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n528), .A2(KEYINPUT73), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n572), .B1(new_n573), .B2(new_n553), .ZN(new_n574));
  INV_X1    g149(.A(G68), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n521), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n539), .A2(G81), .B1(G43), .B2(new_n540), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G860), .ZN(G153));
  AND3_X1   g156(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G36), .ZN(G176));
  NAND2_X1  g158(.A1(G1), .A2(G3), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT77), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT8), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G188));
  NAND2_X1  g162(.A1(new_n540), .A2(G53), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT9), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n539), .A2(G91), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n589), .B(new_n590), .C1(new_n530), .C2(new_n591), .ZN(G299));
  INV_X1    g167(.A(new_n560), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n573), .A2(new_n553), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(G64), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n568), .A2(new_n569), .A3(new_n564), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n569), .B1(new_n568), .B2(new_n564), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n595), .A2(new_n530), .B1(new_n596), .B2(new_n597), .ZN(G301));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  AND3_X1   g174(.A1(new_n551), .A2(new_n599), .A3(new_n556), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n599), .B1(new_n551), .B2(new_n556), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G286));
  OAI21_X1  g178(.A(G651), .B1(new_n594), .B2(G74), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n539), .A2(G87), .B1(G49), .B2(new_n540), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(G288));
  INV_X1    g181(.A(KEYINPUT79), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n544), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G48), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n540), .A2(KEYINPUT79), .A3(G48), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G86), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n528), .A2(new_n544), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n612), .B1(new_n613), .B2(new_n614), .C1(new_n530), .C2(new_n615), .ZN(G305));
  AOI22_X1  g191(.A1(new_n594), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(new_n530), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n539), .A2(G85), .B1(G47), .B2(new_n540), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(G301), .A2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n539), .A2(G92), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT10), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n528), .A2(G66), .ZN(new_n625));
  INV_X1    g200(.A(G79), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n521), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n540), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n621), .B1(new_n630), .B2(G868), .ZN(G284));
  OAI21_X1  g206(.A(new_n621), .B1(new_n630), .B2(G868), .ZN(G321));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n602), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT80), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n635), .B1(G868), .B2(new_n636), .ZN(G297));
  OAI21_X1  g212(.A(new_n635), .B1(G868), .B2(new_n636), .ZN(G280));
  INV_X1    g213(.A(G559), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n630), .B1(new_n639), .B2(G860), .ZN(G148));
  NAND2_X1  g215(.A1(new_n579), .A2(new_n633), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n629), .A2(G559), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n641), .B1(new_n642), .B2(new_n633), .ZN(G323));
  XNOR2_X1  g218(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g219(.A1(new_n471), .A2(G2105), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n474), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  INV_X1    g223(.A(G2100), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT81), .Z(new_n651));
  NAND2_X1  g226(.A1(new_n490), .A2(G123), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  INV_X1    g228(.A(G111), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n653), .B1(new_n654), .B2(G2105), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n497), .B2(G135), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT83), .B(G2096), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n648), .A2(new_n649), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT82), .Z(new_n661));
  NAND3_X1  g236(.A1(new_n651), .A2(new_n659), .A3(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT15), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n665), .A2(G2435), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(G2435), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(KEYINPUT14), .A3(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2443), .B(G2446), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT85), .B(KEYINPUT16), .Z(new_n672));
  XNOR2_X1  g247(.A(G2451), .B(G2454), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT84), .B(KEYINPUT86), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n671), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1341), .B(G1348), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n677), .A2(new_n679), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(G14), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G401));
  XOR2_X1   g260(.A(G2072), .B(G2078), .Z(new_n686));
  XOR2_X1   g261(.A(G2067), .B(G2678), .Z(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2084), .B(G2090), .Z(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n686), .B1(new_n690), .B2(KEYINPUT18), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G2096), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G2100), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(KEYINPUT17), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n688), .A2(new_n689), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT18), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n693), .B(new_n696), .Z(G227));
  XOR2_X1   g272(.A(G1971), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n704), .A2(new_n705), .B1(new_n700), .B2(new_n706), .ZN(new_n707));
  OR3_X1    g282(.A1(new_n700), .A2(new_n703), .A3(new_n706), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n707), .B(new_n708), .C1(new_n705), .C2(new_n704), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1991), .B(G1996), .ZN(new_n712));
  INV_X1    g287(.A(G1981), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n711), .B(new_n715), .ZN(G229));
  NAND3_X1  g291(.A1(new_n490), .A2(KEYINPUT100), .A3(G129), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n488), .B1(new_n485), .B2(G2105), .ZN(new_n718));
  AOI211_X1 g293(.A(KEYINPUT68), .B(new_n493), .C1(new_n482), .C2(new_n484), .ZN(new_n719));
  OAI21_X1  g294(.A(G129), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT100), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n645), .A2(G105), .ZN(new_n724));
  NAND3_X1  g299(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT26), .Z(new_n726));
  INV_X1    g301(.A(G141), .ZN(new_n727));
  OAI211_X1 g302(.A(new_n724), .B(new_n726), .C1(new_n496), .C2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G32), .B(new_n730), .S(G29), .Z(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n732));
  INV_X1    g307(.A(G1996), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n731), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(G162), .A2(G29), .ZN(new_n736));
  OR2_X1    g311(.A1(G29), .A2(G35), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n738), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g315(.A(G2090), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n736), .A2(new_n737), .ZN(new_n742));
  INV_X1    g317(.A(new_n738), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n736), .A2(new_n737), .A3(new_n738), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n630), .A2(G16), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G4), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1348), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n741), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(KEYINPUT90), .A2(G16), .ZN(new_n753));
  NOR2_X1   g328(.A1(KEYINPUT90), .A2(G16), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n580), .B2(new_n756), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT96), .B(G1341), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G29), .A2(G33), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n497), .A2(G139), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n763), .A2(new_n493), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n645), .A2(G103), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  NAND3_X1  g341(.A1(new_n762), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n761), .B1(new_n768), .B2(G29), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G2072), .ZN(new_n770));
  INV_X1    g345(.A(G29), .ZN(new_n771));
  NOR2_X1   g346(.A1(G164), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G27), .B2(new_n771), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n756), .A2(KEYINPUT23), .A3(G20), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT23), .ZN(new_n778));
  INV_X1    g353(.A(G20), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n778), .B1(new_n755), .B2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G16), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n777), .B(new_n780), .C1(new_n636), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT105), .B(G1956), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n773), .A2(new_n774), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n776), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n782), .A2(new_n783), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n657), .A2(new_n771), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n771), .B1(new_n789), .B2(G28), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT103), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n789), .B2(G28), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n787), .A2(new_n788), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n781), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G168), .B2(new_n781), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT102), .B(G1966), .Z(new_n799));
  XOR2_X1   g374(.A(new_n798), .B(new_n799), .Z(new_n800));
  OR2_X1    g375(.A1(KEYINPUT24), .A2(G34), .ZN(new_n801));
  NAND2_X1  g376(.A1(KEYINPUT24), .A2(G34), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n801), .A2(new_n771), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G160), .B2(new_n771), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G2084), .Z(new_n805));
  INV_X1    g380(.A(G11), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n769), .A2(G2072), .B1(KEYINPUT31), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n796), .A2(new_n800), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(G5), .A2(G16), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G171), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1961), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n786), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AND4_X1   g387(.A1(new_n735), .A2(new_n752), .A3(new_n760), .A4(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(KEYINPUT36), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n781), .A2(G23), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n604), .A2(new_n605), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n781), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT33), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n821), .B(new_n817), .C1(new_n818), .C2(new_n781), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G1976), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n756), .A2(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G166), .B2(new_n756), .ZN(new_n827));
  INV_X1    g402(.A(G1971), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n820), .A2(G1976), .A3(new_n822), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n781), .A2(G6), .ZN(new_n831));
  INV_X1    g406(.A(G305), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n831), .B1(new_n832), .B2(new_n781), .ZN(new_n833));
  XNOR2_X1  g408(.A(KEYINPUT32), .B(G1981), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT92), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n833), .B(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n825), .A2(new_n829), .A3(new_n830), .A4(new_n836), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n756), .A2(G24), .ZN(new_n839));
  INV_X1    g414(.A(G290), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n756), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT91), .B(G1986), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n814), .A2(KEYINPUT36), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n771), .A2(G25), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n490), .A2(G119), .ZN(new_n846));
  OAI21_X1  g421(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n847));
  INV_X1    g422(.A(G107), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(G2105), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n497), .B2(G131), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n845), .B1(new_n851), .B2(new_n771), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT35), .B(G1991), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n838), .A2(new_n843), .A3(new_n844), .A4(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT93), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n837), .A2(new_n857), .A3(KEYINPUT34), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n837), .B2(KEYINPUT34), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n816), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n844), .B(new_n855), .C1(new_n837), .C2(KEYINPUT34), .ZN(new_n862));
  INV_X1    g437(.A(new_n843), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n816), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n864), .B(new_n865), .C1(new_n859), .C2(new_n858), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n771), .A2(G26), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  OAI21_X1  g444(.A(G128), .B1(new_n718), .B2(new_n719), .ZN(new_n870));
  OR2_X1    g445(.A1(G104), .A2(G2105), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G116), .C2(new_n493), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT97), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n497), .A2(G140), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n869), .B1(new_n875), .B2(G29), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT99), .B(G2067), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n813), .A2(new_n861), .A3(new_n866), .A4(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n806), .A2(KEYINPUT31), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n749), .A2(new_n750), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR3_X1   g457(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(G311));
  AND3_X1   g458(.A1(new_n813), .A2(new_n861), .A3(new_n866), .ZN(new_n884));
  INV_X1    g459(.A(new_n880), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n885), .A3(new_n881), .A4(new_n878), .ZN(G150));
  INV_X1    g461(.A(G67), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n573), .B2(new_n553), .ZN(new_n888));
  INV_X1    g463(.A(G80), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n521), .ZN(new_n890));
  OAI21_X1  g465(.A(G651), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n539), .A2(G93), .B1(G55), .B2(new_n540), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G860), .ZN(new_n894));
  XOR2_X1   g469(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n577), .A3(new_n578), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n579), .A2(new_n891), .A3(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n630), .A2(G559), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT38), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n900), .B(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n896), .B1(new_n903), .B2(G860), .ZN(G145));
  XNOR2_X1  g479(.A(new_n657), .B(G160), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n499), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n499), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n851), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  INV_X1    g485(.A(new_n851), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n911), .A3(new_n906), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n730), .A2(G164), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n875), .B(KEYINPUT107), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n723), .A2(new_n515), .A3(new_n729), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT107), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n875), .B(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n515), .B1(new_n723), .B2(new_n729), .ZN(new_n920));
  AOI211_X1 g495(.A(G164), .B(new_n728), .C1(new_n717), .C2(new_n722), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n767), .B(KEYINPUT108), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n768), .A2(KEYINPUT108), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n926), .B1(new_n917), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n490), .A2(G130), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n497), .A2(G142), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n493), .A2(G118), .ZN(new_n930));
  OAI21_X1  g505(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT109), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n928), .B(new_n929), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(new_n647), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n925), .A2(new_n927), .A3(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n917), .A2(new_n922), .ZN(new_n937));
  INV_X1    g512(.A(new_n926), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n939), .B2(new_n924), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n913), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n934), .B1(new_n925), .B2(new_n927), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n909), .A2(new_n912), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n939), .A2(new_n924), .A3(new_n936), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n941), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g523(.A1(new_n629), .A2(new_n636), .ZN(new_n949));
  NAND3_X1  g524(.A1(G299), .A2(new_n624), .A3(new_n628), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n899), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n642), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n899), .B1(G559), .B2(new_n629), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(KEYINPUT111), .B(KEYINPUT41), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n949), .A2(new_n950), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT41), .B1(new_n949), .B2(new_n950), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n955), .A2(new_n956), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(G288), .B(G303), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n840), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n965), .A2(new_n840), .ZN(new_n968));
  OAI21_X1  g543(.A(G305), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n965), .A2(new_n840), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(new_n832), .A3(new_n966), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n969), .B2(new_n972), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n957), .B(new_n964), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n969), .A2(new_n972), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT42), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n964), .A2(new_n957), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n969), .A2(new_n972), .A3(new_n970), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n980), .A3(G868), .ZN(new_n981));
  INV_X1    g556(.A(new_n893), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT112), .B1(new_n982), .B2(G868), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n975), .A2(new_n980), .A3(KEYINPUT112), .A4(G868), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(G331));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  NAND2_X1  g562(.A1(G331), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(KEYINPUT113), .A3(new_n985), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(G295));
  OAI211_X1 g565(.A(G171), .B(KEYINPUT115), .C1(new_n600), .C2(new_n601), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n557), .A2(KEYINPUT78), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n551), .A2(new_n599), .A3(new_n556), .ZN(new_n993));
  AOI21_X1  g568(.A(G301), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G171), .B2(new_n557), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n991), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n954), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT115), .B1(G301), .B2(G168), .ZN(new_n999));
  OAI21_X1  g574(.A(G171), .B1(new_n600), .B2(new_n601), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(new_n899), .A3(new_n991), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(KEYINPUT116), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n899), .B1(new_n1001), .B2(new_n991), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n951), .ZN(new_n1008));
  INV_X1    g583(.A(new_n976), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n961), .B1(new_n998), .B2(new_n1002), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g587(.A1(new_n1003), .A2(new_n1006), .B1(new_n949), .B2(new_n950), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n976), .B1(new_n1013), .B2(new_n1010), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1012), .A2(new_n1014), .A3(new_n942), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT44), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1010), .B1(new_n1007), .B2(new_n951), .ZN(new_n1019));
  AOI21_X1  g594(.A(G37), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n951), .A2(KEYINPUT41), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n951), .A2(new_n958), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1003), .A2(new_n1021), .A3(new_n1022), .A4(new_n1006), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n953), .A2(new_n998), .A3(new_n1002), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n976), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1016), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1017), .A2(new_n1018), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1012), .A2(new_n942), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1009), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT43), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1020), .A2(new_n1014), .A3(new_n1027), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1018), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1029), .A2(new_n1034), .ZN(G397));
  NAND2_X1  g610(.A1(new_n466), .A2(new_n467), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n493), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n474), .A2(new_n470), .A3(G125), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT65), .B1(new_n476), .B2(new_n477), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1038), .A2(new_n1039), .B1(G113), .B2(G2104), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1037), .B(G40), .C1(new_n1040), .C2(new_n493), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(G160), .A2(KEYINPUT117), .A3(G40), .ZN(new_n1044));
  INV_X1    g619(.A(G1384), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n515), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1043), .A2(new_n1044), .B1(KEYINPUT50), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n515), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1956), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1046), .B(KEYINPUT45), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT56), .B(G2072), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(G299), .B(KEYINPUT57), .ZN(new_n1057));
  NOR3_X1   g632(.A1(new_n1052), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  INV_X1    g635(.A(G1956), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1046), .A2(KEYINPUT50), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(G160), .B2(G40), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1049), .B(KEYINPUT120), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1053), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1060), .B1(new_n1069), .B2(new_n1057), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1060), .B(new_n1057), .C1(new_n1052), .C2(new_n1056), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(G1348), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1074));
  AOI211_X1 g649(.A(G2067), .B(new_n1046), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1076), .A2(new_n629), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1059), .B1(new_n1073), .B2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT61), .B(new_n1059), .C1(new_n1070), .C2(new_n1072), .ZN(new_n1079));
  NOR4_X1   g654(.A1(new_n1074), .A2(new_n1075), .A3(KEYINPUT60), .A4(new_n629), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(G1996), .ZN(new_n1082));
  XNOR2_X1  g657(.A(KEYINPUT58), .B(G1341), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1046), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1053), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n580), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(KEYINPUT59), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT59), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(new_n580), .C1(new_n1082), .C2(new_n1085), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1080), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  NOR3_X1   g665(.A1(new_n1074), .A2(new_n630), .A3(new_n1075), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT60), .B1(new_n1077), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1079), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT61), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n1095));
  XNOR2_X1  g670(.A(G299), .B(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1094), .B1(new_n1058), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT122), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(new_n1094), .C1(new_n1058), .C2(new_n1097), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1078), .B1(new_n1093), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT119), .B1(G305), .B2(G1981), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n615), .A2(new_n530), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n614), .A2(new_n613), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n713), .A4(new_n612), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(G305), .A2(G1981), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT49), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(G8), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1053), .B2(new_n1084), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1110), .A2(KEYINPUT49), .A3(new_n1111), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n824), .B2(G288), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT52), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1081), .A2(new_n828), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1047), .A2(new_n745), .A3(new_n1049), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1115), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(G303), .A2(G8), .ZN(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(KEYINPUT55), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1047), .A2(new_n745), .A3(new_n1051), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1122), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1130), .B2(G8), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n818), .A2(G1976), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1119), .A2(KEYINPUT52), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1121), .A2(new_n1128), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT53), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1081), .B2(G2078), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1053), .A2(new_n1062), .A3(new_n1049), .ZN(new_n1138));
  INV_X1    g713(.A(G1961), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n468), .A2(new_n1136), .ZN(new_n1142));
  INV_X1    g717(.A(G40), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1040), .A2(KEYINPUT125), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n493), .B1(new_n1040), .B2(KEYINPUT125), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1054), .A2(new_n774), .A3(new_n1142), .A4(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(G301), .B1(new_n1141), .B2(new_n1147), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT53), .A3(new_n774), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1150), .A2(new_n1137), .A3(new_n1140), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n1151), .B2(G171), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1154));
  NAND3_X1  g729(.A1(new_n1141), .A2(G301), .A3(new_n1147), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1151), .A2(G171), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1135), .A2(new_n1153), .A3(new_n1157), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1149), .A2(new_n799), .B1(new_n1138), .B2(G2084), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(G8), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT51), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(KEYINPUT123), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n557), .A2(G8), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1160), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1161), .A2(KEYINPUT123), .ZN(new_n1166));
  OAI211_X1 g741(.A(G8), .B(new_n1162), .C1(new_n1159), .C2(new_n557), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1160), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n557), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1103), .A2(new_n1158), .A3(new_n1171), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1169), .B(new_n602), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1134), .A2(new_n1120), .A3(new_n1118), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT63), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1118), .A2(new_n824), .A3(new_n818), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1110), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n1116), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT63), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1159), .A2(new_n1179), .A3(G8), .A4(new_n602), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1128), .B1(new_n1131), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1181), .A2(new_n1121), .A3(new_n1134), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1175), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1171), .A2(KEYINPUT62), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1135), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1168), .A2(new_n1186), .A3(new_n1170), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1156), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1184), .A2(new_n1185), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1172), .A2(new_n1183), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n851), .A2(new_n854), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n730), .B(new_n733), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n911), .A2(new_n853), .ZN(new_n1193));
  XOR2_X1   g768(.A(new_n875), .B(G2067), .Z(new_n1194));
  AND4_X1   g769(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(G290), .A2(G1986), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(KEYINPUT118), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(G1986), .B2(G290), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  AOI211_X1 g774(.A(KEYINPUT45), .B(new_n1084), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1190), .A2(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(new_n1191), .B(KEYINPUT126), .Z(new_n1203));
  NAND2_X1  g778(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1203), .B1(new_n1204), .B2(new_n1200), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n875), .A2(G2067), .ZN(new_n1207));
  OR3_X1    g782(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1205), .B2(new_n1207), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1208), .A2(new_n1200), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g785(.A(new_n1194), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1200), .B1(new_n1211), .B2(new_n730), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1200), .A2(new_n733), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1213), .B(KEYINPUT46), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g790(.A(new_n1215), .B(KEYINPUT47), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT48), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1200), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1218), .B1(new_n1219), .B2(new_n1195), .ZN(new_n1220));
  AND3_X1   g795(.A1(new_n1210), .A2(new_n1216), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1202), .A2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g797(.A1(G229), .A2(new_n460), .ZN(new_n1224));
  AND4_X1   g798(.A1(new_n942), .A2(new_n1026), .A3(new_n1012), .A4(new_n1027), .ZN(new_n1225));
  AOI21_X1  g799(.A(new_n1027), .B1(new_n1020), .B2(new_n1014), .ZN(new_n1226));
  OAI211_X1 g800(.A(new_n947), .B(new_n1224), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g801(.A(G227), .B1(new_n681), .B2(new_n683), .ZN(new_n1228));
  INV_X1    g802(.A(new_n1228), .ZN(new_n1229));
  NOR2_X1   g803(.A1(new_n1227), .A2(new_n1229), .ZN(G308));
  NAND2_X1  g804(.A1(new_n1017), .A2(new_n1028), .ZN(new_n1231));
  NAND4_X1  g805(.A1(new_n1231), .A2(new_n1228), .A3(new_n947), .A4(new_n1224), .ZN(G225));
endmodule


