

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U552 ( .A1(n706), .A2(n705), .ZN(n756) );
  XNOR2_X1 U553 ( .A(n764), .B(n763), .ZN(n777) );
  XNOR2_X1 U554 ( .A(n746), .B(KEYINPUT30), .ZN(n748) );
  XNOR2_X1 U555 ( .A(n551), .B(n550), .ZN(n552) );
  INV_X1 U556 ( .A(KEYINPUT23), .ZN(n550) );
  XNOR2_X2 U557 ( .A(n537), .B(n536), .ZN(n581) );
  NOR2_X1 U558 ( .A1(n779), .A2(n783), .ZN(n518) );
  AND2_X1 U559 ( .A1(G138), .A2(n882), .ZN(n519) );
  AND2_X1 U560 ( .A1(n525), .A2(n524), .ZN(n520) );
  XOR2_X1 U561 ( .A(KEYINPUT31), .B(n752), .Z(n521) );
  NOR2_X1 U562 ( .A1(n710), .A2(n709), .ZN(n719) );
  INV_X1 U563 ( .A(G168), .ZN(n747) );
  AND2_X1 U564 ( .A1(n748), .A2(n747), .ZN(n751) );
  INV_X1 U565 ( .A(KEYINPUT29), .ZN(n735) );
  INV_X1 U566 ( .A(KEYINPUT105), .ZN(n754) );
  XNOR2_X1 U567 ( .A(n755), .B(n754), .ZN(n761) );
  NOR2_X1 U568 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U569 ( .A1(G8), .A2(n756), .ZN(n799) );
  XNOR2_X1 U570 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U571 ( .A1(G2105), .A2(n526), .ZN(n549) );
  NOR2_X1 U572 ( .A1(n586), .A2(n585), .ZN(n587) );
  BUF_X1 U573 ( .A(n545), .Z(n882) );
  NOR2_X1 U574 ( .A1(G651), .A2(n644), .ZN(n648) );
  NOR2_X1 U575 ( .A1(n644), .A2(n535), .ZN(n653) );
  NAND2_X1 U576 ( .A1(n520), .A2(n527), .ZN(n528) );
  NOR2_X1 U577 ( .A1(n556), .A2(n555), .ZN(G160) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U579 ( .A(n523), .B(n522), .ZN(n545) );
  INV_X1 U580 ( .A(G2104), .ZN(n526) );
  AND2_X1 U581 ( .A1(n526), .A2(G2105), .ZN(n874) );
  NAND2_X1 U582 ( .A1(G126), .A2(n874), .ZN(n525) );
  AND2_X1 U583 ( .A1(G2104), .A2(G2105), .ZN(n875) );
  NAND2_X1 U584 ( .A1(G114), .A2(n875), .ZN(n524) );
  BUF_X1 U585 ( .A(n549), .Z(n880) );
  NAND2_X1 U586 ( .A1(G102), .A2(n880), .ZN(n527) );
  NOR2_X1 U587 ( .A1(n519), .A2(n528), .ZN(G164) );
  NOR2_X1 U588 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U589 ( .A1(n652), .A2(G89), .ZN(n529) );
  XNOR2_X1 U590 ( .A(KEYINPUT4), .B(n529), .ZN(n532) );
  XOR2_X1 U591 ( .A(KEYINPUT0), .B(G543), .Z(n644) );
  INV_X1 U592 ( .A(G651), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n653), .A2(G76), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT79), .B(n530), .Z(n531) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(KEYINPUT5), .ZN(n543) );
  XNOR2_X1 U597 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT68), .ZN(n537) );
  NOR2_X1 U599 ( .A1(G543), .A2(n535), .ZN(n536) );
  NAND2_X1 U600 ( .A1(G63), .A2(n581), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(KEYINPUT80), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G51), .A2(n648), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U604 ( .A(KEYINPUT6), .B(n541), .Z(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U606 ( .A(n544), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U607 ( .A1(G137), .A2(n545), .ZN(n547) );
  NAND2_X1 U608 ( .A1(G113), .A2(n875), .ZN(n546) );
  NAND2_X1 U609 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U610 ( .A(KEYINPUT66), .B(n548), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n874), .A2(G125), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n549), .A2(G101), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n554), .B(KEYINPUT64), .ZN(n555) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G57), .ZN(G237) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  NAND2_X1 U618 ( .A1(n648), .A2(G52), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G64), .A2(n581), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n652), .A2(G90), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT70), .ZN(n561) );
  NAND2_X1 U623 ( .A1(G77), .A2(n653), .ZN(n560) );
  NAND2_X1 U624 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT71), .B(n565), .Z(G171) );
  XOR2_X1 U628 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n567) );
  NAND2_X1 U629 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n567), .B(n566), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n834) );
  NAND2_X1 U632 ( .A1(n834), .A2(G567), .ZN(n568) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n568), .Z(G234) );
  NAND2_X1 U634 ( .A1(n652), .A2(G81), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT12), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G68), .A2(n653), .ZN(n570) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(KEYINPUT76), .Z(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n576) );
  NAND2_X1 U640 ( .A1(G56), .A2(n581), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n574), .Z(n575) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n648), .A2(G43), .ZN(n577) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n941) );
  INV_X1 U645 ( .A(G860), .ZN(n601) );
  OR2_X1 U646 ( .A1(n941), .A2(n601), .ZN(G153) );
  INV_X1 U647 ( .A(G171), .ZN(G301) );
  NAND2_X1 U648 ( .A1(G79), .A2(n653), .ZN(n580) );
  NAND2_X1 U649 ( .A1(G54), .A2(n648), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n580), .A2(n579), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G92), .A2(n652), .ZN(n583) );
  NAND2_X1 U652 ( .A1(G66), .A2(n581), .ZN(n582) );
  NAND2_X1 U653 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT77), .B(n584), .Z(n585) );
  XOR2_X1 U655 ( .A(KEYINPUT15), .B(n587), .Z(n923) );
  NOR2_X1 U656 ( .A1(n923), .A2(G868), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT78), .B(n588), .Z(n590) );
  NAND2_X1 U658 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(G284) );
  XOR2_X1 U660 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U661 ( .A1(G91), .A2(n652), .ZN(n591) );
  XOR2_X1 U662 ( .A(KEYINPUT72), .B(n591), .Z(n596) );
  NAND2_X1 U663 ( .A1(n648), .A2(G53), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G65), .A2(n581), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U666 ( .A(KEYINPUT73), .B(n594), .Z(n595) );
  NOR2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n653), .A2(G78), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(G299) );
  INV_X1 U670 ( .A(G868), .ZN(n666) );
  NOR2_X1 U671 ( .A1(G286), .A2(n666), .ZN(n600) );
  NOR2_X1 U672 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U674 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n602), .A2(n923), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G868), .A2(n941), .ZN(n606) );
  NAND2_X1 U678 ( .A1(G868), .A2(n923), .ZN(n604) );
  NOR2_X1 U679 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G123), .A2(n874), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT18), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n880), .A2(G99), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G135), .A2(n882), .ZN(n611) );
  NAND2_X1 U686 ( .A1(G111), .A2(n875), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(n1004) );
  XNOR2_X1 U689 ( .A(G2096), .B(n1004), .ZN(n615) );
  INV_X1 U690 ( .A(G2100), .ZN(n614) );
  NAND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(G156) );
  NAND2_X1 U692 ( .A1(n923), .A2(G559), .ZN(n664) );
  XNOR2_X1 U693 ( .A(n941), .B(n664), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n616), .A2(G860), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G93), .A2(n652), .ZN(n618) );
  NAND2_X1 U696 ( .A1(G80), .A2(n653), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n648), .A2(G55), .ZN(n620) );
  NAND2_X1 U699 ( .A1(G67), .A2(n581), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(n621) );
  OR2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n667) );
  XOR2_X1 U702 ( .A(n623), .B(n667), .Z(G145) );
  NAND2_X1 U703 ( .A1(G73), .A2(n653), .ZN(n624) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n624), .Z(n631) );
  NAND2_X1 U705 ( .A1(n652), .A2(G86), .ZN(n625) );
  XNOR2_X1 U706 ( .A(KEYINPUT83), .B(n625), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G61), .A2(n581), .ZN(n626) );
  XOR2_X1 U708 ( .A(KEYINPUT82), .B(n626), .Z(n627) );
  NOR2_X1 U709 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U710 ( .A(KEYINPUT84), .B(n629), .Z(n630) );
  NOR2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U712 ( .A1(n648), .A2(G48), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G85), .A2(n652), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G72), .A2(n653), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U717 ( .A(KEYINPUT67), .B(n636), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n581), .A2(G60), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n648), .A2(G47), .ZN(n637) );
  AND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(G290) );
  NAND2_X1 U722 ( .A1(G49), .A2(n648), .ZN(n642) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n641) );
  NAND2_X1 U724 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U725 ( .A1(n581), .A2(n643), .ZN(n647) );
  NAND2_X1 U726 ( .A1(G87), .A2(n644), .ZN(n645) );
  XOR2_X1 U727 ( .A(KEYINPUT81), .B(n645), .Z(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U729 ( .A1(n648), .A2(G50), .ZN(n650) );
  NAND2_X1 U730 ( .A1(G62), .A2(n581), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U732 ( .A(KEYINPUT85), .B(n651), .ZN(n657) );
  NAND2_X1 U733 ( .A1(G88), .A2(n652), .ZN(n655) );
  NAND2_X1 U734 ( .A1(G75), .A2(n653), .ZN(n654) );
  AND2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(G303) );
  INV_X1 U737 ( .A(G303), .ZN(G166) );
  XOR2_X1 U738 ( .A(n667), .B(G290), .Z(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT19), .B(n941), .Z(n658) );
  XNOR2_X1 U740 ( .A(G288), .B(n658), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U742 ( .A(G305), .B(n661), .ZN(n663) );
  INV_X1 U743 ( .A(G299), .ZN(n730) );
  XNOR2_X1 U744 ( .A(n730), .B(G166), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n663), .B(n662), .ZN(n903) );
  XOR2_X1 U746 ( .A(n903), .B(n664), .Z(n665) );
  NAND2_X1 U747 ( .A1(G868), .A2(n665), .ZN(n669) );
  NAND2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U754 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U756 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  NOR2_X1 U757 ( .A1(G219), .A2(G220), .ZN(n674) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U759 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G96), .A2(n676), .ZN(n839) );
  AND2_X1 U761 ( .A1(G2106), .A2(n839), .ZN(n681) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n677) );
  NOR2_X1 U763 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U764 ( .A1(G108), .A2(n678), .ZN(n838) );
  NAND2_X1 U765 ( .A1(G567), .A2(n838), .ZN(n679) );
  XOR2_X1 U766 ( .A(KEYINPUT86), .B(n679), .Z(n680) );
  NOR2_X1 U767 ( .A1(n681), .A2(n680), .ZN(G319) );
  INV_X1 U768 ( .A(G319), .ZN(n683) );
  NAND2_X1 U769 ( .A1(G661), .A2(G483), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n683), .A2(n682), .ZN(n837) );
  NAND2_X1 U771 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U772 ( .A1(G119), .A2(n874), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G107), .A2(n875), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U775 ( .A(KEYINPUT89), .B(n686), .ZN(n690) );
  NAND2_X1 U776 ( .A1(G131), .A2(n882), .ZN(n688) );
  NAND2_X1 U777 ( .A1(G95), .A2(n880), .ZN(n687) );
  AND2_X1 U778 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U779 ( .A1(n690), .A2(n689), .ZN(n888) );
  XNOR2_X1 U780 ( .A(KEYINPUT90), .B(G1991), .ZN(n988) );
  NAND2_X1 U781 ( .A1(n888), .A2(n988), .ZN(n700) );
  NAND2_X1 U782 ( .A1(G129), .A2(n874), .ZN(n692) );
  NAND2_X1 U783 ( .A1(G117), .A2(n875), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n880), .A2(G105), .ZN(n693) );
  XOR2_X1 U786 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U788 ( .A(KEYINPUT91), .B(n696), .Z(n698) );
  NAND2_X1 U789 ( .A1(n882), .A2(G141), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n887) );
  NAND2_X1 U791 ( .A1(G1996), .A2(n887), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n1005) );
  NOR2_X1 U793 ( .A1(G164), .A2(G1384), .ZN(n705) );
  NAND2_X1 U794 ( .A1(G160), .A2(G40), .ZN(n704) );
  NOR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n829) );
  NAND2_X1 U796 ( .A1(n1005), .A2(n829), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n701), .B(KEYINPUT92), .ZN(n703) );
  XNOR2_X1 U798 ( .A(G1986), .B(G290), .ZN(n945) );
  NAND2_X1 U799 ( .A1(n945), .A2(n829), .ZN(n702) );
  NAND2_X1 U800 ( .A1(n703), .A2(n702), .ZN(n805) );
  INV_X1 U801 ( .A(n704), .ZN(n706) );
  INV_X1 U802 ( .A(G1996), .ZN(n978) );
  NOR2_X1 U803 ( .A1(n756), .A2(n978), .ZN(n707) );
  XNOR2_X1 U804 ( .A(n707), .B(KEYINPUT26), .ZN(n710) );
  AND2_X1 U805 ( .A1(n756), .A2(G1341), .ZN(n708) );
  OR2_X1 U806 ( .A1(n708), .A2(n941), .ZN(n709) );
  NAND2_X1 U807 ( .A1(n719), .A2(n923), .ZN(n711) );
  XNOR2_X1 U808 ( .A(n711), .B(KEYINPUT100), .ZN(n718) );
  NAND2_X1 U809 ( .A1(G1348), .A2(n756), .ZN(n712) );
  XOR2_X1 U810 ( .A(KEYINPUT101), .B(n712), .Z(n715) );
  INV_X1 U811 ( .A(KEYINPUT96), .ZN(n713) );
  XNOR2_X1 U812 ( .A(n756), .B(n713), .ZN(n723) );
  NAND2_X1 U813 ( .A1(G2067), .A2(n723), .ZN(n714) );
  NAND2_X1 U814 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U815 ( .A(KEYINPUT102), .B(n716), .ZN(n717) );
  NAND2_X1 U816 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U817 ( .A1(n923), .A2(n719), .ZN(n720) );
  XNOR2_X1 U818 ( .A(n720), .B(KEYINPUT103), .ZN(n721) );
  NAND2_X1 U819 ( .A1(n722), .A2(n721), .ZN(n728) );
  NAND2_X1 U820 ( .A1(G2072), .A2(n723), .ZN(n724) );
  XNOR2_X1 U821 ( .A(n724), .B(KEYINPUT27), .ZN(n726) );
  XOR2_X1 U822 ( .A(G1956), .B(KEYINPUT98), .Z(n950) );
  NOR2_X1 U823 ( .A1(n723), .A2(n950), .ZN(n725) );
  NOR2_X1 U824 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U825 ( .A1(n730), .A2(n729), .ZN(n727) );
  NAND2_X1 U826 ( .A1(n728), .A2(n727), .ZN(n734) );
  NOR2_X1 U827 ( .A1(n730), .A2(n729), .ZN(n732) );
  XNOR2_X1 U828 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n731) );
  XNOR2_X1 U829 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U830 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U831 ( .A(n736), .B(n735), .ZN(n741) );
  XNOR2_X1 U832 ( .A(G1961), .B(KEYINPUT95), .ZN(n968) );
  NAND2_X1 U833 ( .A1(n756), .A2(n968), .ZN(n738) );
  XNOR2_X1 U834 ( .A(G2078), .B(KEYINPUT25), .ZN(n977) );
  NAND2_X1 U835 ( .A1(n723), .A2(n977), .ZN(n737) );
  NAND2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n749) );
  AND2_X1 U837 ( .A1(n749), .A2(G171), .ZN(n739) );
  XNOR2_X1 U838 ( .A(n739), .B(KEYINPUT97), .ZN(n740) );
  NAND2_X1 U839 ( .A1(n741), .A2(n740), .ZN(n753) );
  NOR2_X1 U840 ( .A1(G1966), .A2(n799), .ZN(n743) );
  INV_X1 U841 ( .A(KEYINPUT94), .ZN(n742) );
  XNOR2_X1 U842 ( .A(n743), .B(n742), .ZN(n765) );
  INV_X1 U843 ( .A(G8), .ZN(n744) );
  NOR2_X1 U844 ( .A1(G2084), .A2(n756), .ZN(n766) );
  NOR2_X1 U845 ( .A1(n744), .A2(n766), .ZN(n745) );
  AND2_X1 U846 ( .A1(n765), .A2(n745), .ZN(n746) );
  NOR2_X1 U847 ( .A1(G171), .A2(n749), .ZN(n750) );
  NOR2_X1 U848 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U849 ( .A1(n753), .A2(n521), .ZN(n768) );
  NAND2_X1 U850 ( .A1(G286), .A2(n768), .ZN(n755) );
  NOR2_X1 U851 ( .A1(G1971), .A2(n799), .ZN(n758) );
  NOR2_X1 U852 ( .A1(G2090), .A2(n756), .ZN(n757) );
  NOR2_X1 U853 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U854 ( .A1(G303), .A2(n759), .ZN(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U856 ( .A1(n762), .A2(G8), .ZN(n764) );
  INV_X1 U857 ( .A(KEYINPUT32), .ZN(n763) );
  INV_X1 U858 ( .A(n765), .ZN(n770) );
  NAND2_X1 U859 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U862 ( .A(n771), .B(KEYINPUT104), .ZN(n779) );
  NOR2_X1 U863 ( .A1(n777), .A2(n779), .ZN(n774) );
  NAND2_X1 U864 ( .A1(G166), .A2(G8), .ZN(n772) );
  NOR2_X1 U865 ( .A1(G2090), .A2(n772), .ZN(n773) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U867 ( .A(n775), .B(KEYINPUT107), .ZN(n776) );
  NAND2_X1 U868 ( .A1(n776), .A2(n799), .ZN(n796) );
  INV_X1 U869 ( .A(n777), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G288), .A2(G1976), .ZN(n778) );
  XNOR2_X1 U871 ( .A(n778), .B(KEYINPUT106), .ZN(n925) );
  INV_X1 U872 ( .A(n925), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n780), .A2(n518), .ZN(n785) );
  NOR2_X1 U874 ( .A1(G1976), .A2(G288), .ZN(n924) );
  NOR2_X1 U875 ( .A1(G1971), .A2(G303), .ZN(n781) );
  NOR2_X1 U876 ( .A1(n924), .A2(n781), .ZN(n782) );
  OR2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n784) );
  AND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n924), .A2(KEYINPUT33), .ZN(n786) );
  NOR2_X1 U880 ( .A1(n786), .A2(n799), .ZN(n788) );
  XOR2_X1 U881 ( .A(G1981), .B(G305), .Z(n935) );
  INV_X1 U882 ( .A(n935), .ZN(n787) );
  NOR2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n792) );
  INV_X1 U884 ( .A(n792), .ZN(n789) );
  OR2_X1 U885 ( .A1(n799), .A2(n789), .ZN(n790) );
  AND2_X1 U886 ( .A1(n792), .A2(KEYINPUT33), .ZN(n793) );
  NOR2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U888 ( .A1(n796), .A2(n795), .ZN(n802) );
  NOR2_X1 U889 ( .A1(G1981), .A2(G305), .ZN(n797) );
  XNOR2_X1 U890 ( .A(n797), .B(KEYINPUT24), .ZN(n798) );
  XNOR2_X1 U891 ( .A(n798), .B(KEYINPUT93), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U894 ( .A(n803), .B(KEYINPUT108), .ZN(n804) );
  NOR2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n817) );
  NAND2_X1 U896 ( .A1(G140), .A2(n882), .ZN(n807) );
  NAND2_X1 U897 ( .A1(G104), .A2(n880), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n807), .A2(n806), .ZN(n809) );
  XOR2_X1 U899 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n808) );
  XNOR2_X1 U900 ( .A(n809), .B(n808), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G128), .A2(n874), .ZN(n811) );
  NAND2_X1 U902 ( .A1(G116), .A2(n875), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT35), .B(n812), .Z(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT36), .B(n815), .ZN(n900) );
  XNOR2_X1 U907 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U908 ( .A1(n900), .A2(n826), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n816), .B(KEYINPUT88), .ZN(n1017) );
  NAND2_X1 U910 ( .A1(n829), .A2(n1017), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n817), .A2(n824), .ZN(n831) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n887), .ZN(n1010) );
  NOR2_X1 U913 ( .A1(n988), .A2(n888), .ZN(n1006) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U915 ( .A1(n1006), .A2(n818), .ZN(n819) );
  XOR2_X1 U916 ( .A(KEYINPUT109), .B(n819), .Z(n820) );
  NOR2_X1 U917 ( .A1(n1005), .A2(n820), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n821), .B(KEYINPUT110), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n1010), .A2(n822), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT39), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n826), .A2(n900), .ZN(n1014) );
  NAND2_X1 U923 ( .A1(n827), .A2(n1014), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n831), .A2(n830), .ZN(n833) );
  XOR2_X1 U926 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n832) );
  XNOR2_X1 U927 ( .A(n833), .B(n832), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U930 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U934 ( .A(G120), .ZN(G236) );
  INV_X1 U935 ( .A(G96), .ZN(G221) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  XOR2_X1 U939 ( .A(KEYINPUT42), .B(G2084), .Z(n841) );
  XNOR2_X1 U940 ( .A(G2072), .B(G2078), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U942 ( .A(n842), .B(G2096), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(KEYINPUT43), .B(KEYINPUT113), .Z(n846) );
  XNOR2_X1 U946 ( .A(G2678), .B(G2100), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n848), .B(n847), .Z(G227) );
  XNOR2_X1 U949 ( .A(G1961), .B(G2474), .ZN(n858) );
  XOR2_X1 U950 ( .A(G1976), .B(G1971), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1986), .B(G1956), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U953 ( .A(G1981), .B(G1966), .Z(n852) );
  XNOR2_X1 U954 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U957 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U960 ( .A1(G124), .A2(n874), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n859), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n880), .A2(G100), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U964 ( .A1(G136), .A2(n882), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G112), .A2(n875), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U968 ( .A1(G130), .A2(n874), .ZN(n867) );
  NAND2_X1 U969 ( .A1(G118), .A2(n875), .ZN(n866) );
  NAND2_X1 U970 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U971 ( .A1(G142), .A2(n882), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G106), .A2(n880), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n870), .Z(n871) );
  NOR2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U976 ( .A(G160), .B(n873), .ZN(n899) );
  XNOR2_X1 U977 ( .A(KEYINPUT117), .B(KEYINPUT47), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G127), .A2(n874), .ZN(n877) );
  NAND2_X1 U979 ( .A1(G115), .A2(n875), .ZN(n876) );
  NAND2_X1 U980 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n880), .A2(G103), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n881), .B(KEYINPUT116), .ZN(n884) );
  NAND2_X1 U984 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  NOR2_X1 U986 ( .A1(n886), .A2(n885), .ZN(n999) );
  XNOR2_X1 U987 ( .A(n999), .B(n887), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n892) );
  XNOR2_X1 U989 ( .A(G164), .B(G162), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n890), .B(n1004), .ZN(n891) );
  XOR2_X1 U991 ( .A(n892), .B(n891), .Z(n897) );
  XOR2_X1 U992 ( .A(KEYINPUT115), .B(KEYINPUT118), .Z(n894) );
  XNOR2_X1 U993 ( .A(KEYINPUT119), .B(KEYINPUT46), .ZN(n893) );
  XNOR2_X1 U994 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U995 ( .A(KEYINPUT48), .B(n895), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1000 ( .A(G171), .B(G286), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n905), .B(n923), .ZN(n906) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n906), .ZN(G397) );
  XOR2_X1 U1004 ( .A(KEYINPUT112), .B(G2446), .Z(n908) );
  XNOR2_X1 U1005 ( .A(G2443), .B(G2454), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1007 ( .A(n909), .B(G2451), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G1341), .B(G1348), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1010 ( .A(G2435), .B(G2427), .Z(n913) );
  XNOR2_X1 U1011 ( .A(G2430), .B(G2438), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1013 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1014 ( .A1(G14), .A2(n916), .ZN(n922) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(G108), .ZN(G238) );
  INV_X1 U1023 ( .A(n922), .ZN(G401) );
  XNOR2_X1 U1024 ( .A(G16), .B(KEYINPUT56), .ZN(n949) );
  XNOR2_X1 U1025 ( .A(n923), .B(G1348), .ZN(n934) );
  INV_X1 U1026 ( .A(n924), .ZN(n926) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT125), .ZN(n930) );
  XNOR2_X1 U1029 ( .A(G171), .B(G1961), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(n928), .B(KEYINPUT124), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G1956), .B(G299), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n940) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G168), .ZN(n936) );
  NAND2_X1 U1036 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1037 ( .A(n937), .B(KEYINPUT57), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT123), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n947) );
  XOR2_X1 U1040 ( .A(n941), .B(G1341), .Z(n943) );
  XNOR2_X1 U1041 ( .A(G166), .B(G1971), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n1028) );
  XNOR2_X1 U1046 ( .A(n950), .B(G20), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(G6), .B(G1981), .ZN(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1051 ( .A(KEYINPUT59), .B(G1348), .Z(n955) );
  XNOR2_X1 U1052 ( .A(G4), .B(n955), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(KEYINPUT126), .B(n958), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(n959), .B(KEYINPUT60), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(G1986), .B(G24), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(G1971), .B(KEYINPUT127), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(n962), .B(G22), .ZN(n963) );
  NAND2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1062 ( .A(KEYINPUT58), .B(n965), .Z(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n972) );
  XOR2_X1 U1064 ( .A(G1966), .B(G21), .Z(n970) );
  XNOR2_X1 U1065 ( .A(n968), .B(G5), .ZN(n969) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NOR2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1068 ( .A(KEYINPUT61), .B(n973), .ZN(n975) );
  INV_X1 U1069 ( .A(G16), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n976), .A2(G11), .ZN(n1026) );
  XOR2_X1 U1072 ( .A(n977), .B(G27), .Z(n980) );
  XOR2_X1 U1073 ( .A(n978), .B(G32), .Z(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(KEYINPUT122), .B(n981), .ZN(n987) );
  XOR2_X1 U1076 ( .A(G2072), .B(G33), .Z(n982) );
  NAND2_X1 U1077 ( .A1(G28), .A2(n982), .ZN(n985) );
  XOR2_X1 U1078 ( .A(KEYINPUT121), .B(G2067), .Z(n983) );
  XNOR2_X1 U1079 ( .A(G26), .B(n983), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(G25), .B(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1084 ( .A(KEYINPUT53), .B(n991), .Z(n994) );
  XOR2_X1 U1085 ( .A(G34), .B(KEYINPUT54), .Z(n992) );
  XNOR2_X1 U1086 ( .A(G2084), .B(n992), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G35), .B(G2090), .ZN(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(G29), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(n998), .B(KEYINPUT55), .ZN(n1024) );
  XOR2_X1 U1092 ( .A(G2072), .B(n999), .Z(n1001) );
  XOR2_X1 U1093 ( .A(G164), .B(G2078), .Z(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1002), .ZN(n1020) );
  XOR2_X1 U1096 ( .A(G2084), .B(G160), .Z(n1003) );
  NOR2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1013) );
  XOR2_X1 U1100 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(n1011), .B(KEYINPUT51), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT120), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1021), .ZN(n1022) );
  NAND2_X1 U1109 ( .A1(G29), .A2(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1113 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

