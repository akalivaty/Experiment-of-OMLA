

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U325 ( .A(n343), .B(n342), .ZN(n365) );
  NOR2_X2 U326 ( .A1(n415), .A2(n521), .ZN(n416) );
  XNOR2_X1 U327 ( .A(n306), .B(n305), .ZN(n579) );
  XNOR2_X1 U328 ( .A(KEYINPUT125), .B(n572), .ZN(n580) );
  XOR2_X1 U329 ( .A(KEYINPUT65), .B(n416), .Z(n293) );
  INV_X1 U330 ( .A(KEYINPUT68), .ZN(n335) );
  XNOR2_X1 U331 ( .A(n336), .B(n335), .ZN(n338) );
  INV_X1 U332 ( .A(KEYINPUT32), .ZN(n298) );
  XNOR2_X1 U333 ( .A(n338), .B(n337), .ZN(n352) );
  XNOR2_X1 U334 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U335 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n372) );
  XNOR2_X1 U336 ( .A(n373), .B(n372), .ZN(n533) );
  BUF_X1 U337 ( .A(n533), .Z(n551) );
  NOR2_X1 U338 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U339 ( .A(n362), .B(KEYINPUT41), .ZN(n562) );
  XNOR2_X1 U340 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U341 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(G85GAT), .B(G92GAT), .Z(n295) );
  XNOR2_X1 U343 ( .A(G99GAT), .B(G106GAT), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n334) );
  XNOR2_X1 U345 ( .A(n334), .B(KEYINPUT33), .ZN(n297) );
  AND2_X1 U346 ( .A1(G230GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U348 ( .A(G176GAT), .B(G64GAT), .Z(n387) );
  XNOR2_X1 U349 ( .A(n387), .B(KEYINPUT31), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U351 ( .A(KEYINPUT13), .B(G57GAT), .Z(n309) );
  XNOR2_X1 U352 ( .A(n302), .B(n309), .ZN(n306) );
  XOR2_X1 U353 ( .A(G120GAT), .B(G71GAT), .Z(n442) );
  XOR2_X1 U354 ( .A(G78GAT), .B(G148GAT), .Z(n304) );
  XNOR2_X1 U355 ( .A(KEYINPUT70), .B(G204GAT), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n420) );
  XOR2_X1 U357 ( .A(n442), .B(n420), .Z(n305) );
  XOR2_X1 U358 ( .A(G211GAT), .B(G71GAT), .Z(n308) );
  XNOR2_X1 U359 ( .A(G183GAT), .B(G127GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n310) );
  XOR2_X1 U361 ( .A(n310), .B(n309), .Z(n312) );
  XNOR2_X1 U362 ( .A(G22GAT), .B(G155GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n317) );
  XNOR2_X1 U364 ( .A(G15GAT), .B(G1GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n313), .B(KEYINPUT69), .ZN(n356) );
  XOR2_X1 U366 ( .A(n356), .B(G64GAT), .Z(n315) );
  NAND2_X1 U367 ( .A1(G231GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U369 ( .A(n317), .B(n316), .Z(n325) );
  XOR2_X1 U370 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n319) );
  XNOR2_X1 U371 ( .A(G78GAT), .B(KEYINPUT79), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U373 ( .A(KEYINPUT12), .B(KEYINPUT78), .Z(n321) );
  XNOR2_X1 U374 ( .A(G8GAT), .B(KEYINPUT77), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(n325), .B(n324), .Z(n475) );
  INV_X1 U378 ( .A(n475), .ZN(n583) );
  XOR2_X1 U379 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT9), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT75), .B(KEYINPUT73), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(n428), .B(n328), .Z(n330) );
  NAND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n343) );
  XOR2_X1 U386 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n332) );
  XNOR2_X1 U387 ( .A(G134GAT), .B(KEYINPUT74), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U389 ( .A(n334), .B(n333), .Z(n341) );
  XNOR2_X1 U390 ( .A(G43GAT), .B(G29GAT), .ZN(n336) );
  XOR2_X1 U391 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n337) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(G190GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n339), .B(G218GAT), .ZN(n382) );
  XNOR2_X1 U394 ( .A(n352), .B(n382), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X2 U396 ( .A(n365), .B(KEYINPUT76), .Z(n545) );
  XNOR2_X1 U397 ( .A(KEYINPUT36), .B(n545), .ZN(n586) );
  NOR2_X1 U398 ( .A1(n583), .A2(n586), .ZN(n345) );
  XNOR2_X1 U399 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n359) );
  XOR2_X1 U401 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n347) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U404 ( .A(n348), .B(KEYINPUT67), .Z(n354) );
  XOR2_X1 U405 ( .A(G197GAT), .B(G113GAT), .Z(n350) );
  XNOR2_X1 U406 ( .A(G50GAT), .B(G36GAT), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U410 ( .A(G169GAT), .B(G8GAT), .Z(n388) );
  XOR2_X1 U411 ( .A(n355), .B(n388), .Z(n358) );
  XOR2_X1 U412 ( .A(G141GAT), .B(G22GAT), .Z(n429) );
  XNOR2_X1 U413 ( .A(n429), .B(n356), .ZN(n357) );
  XOR2_X1 U414 ( .A(n358), .B(n357), .Z(n507) );
  INV_X1 U415 ( .A(n507), .ZN(n573) );
  NAND2_X1 U416 ( .A1(n359), .A2(n573), .ZN(n360) );
  NOR2_X1 U417 ( .A1(n579), .A2(n360), .ZN(n361) );
  XNOR2_X1 U418 ( .A(KEYINPUT111), .B(n361), .ZN(n371) );
  XNOR2_X1 U419 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n579), .B(KEYINPUT64), .ZN(n362) );
  NOR2_X1 U421 ( .A1(n573), .A2(n562), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n367) );
  INV_X1 U423 ( .A(n365), .ZN(n560) );
  NOR2_X1 U424 ( .A1(n475), .A2(n365), .ZN(n366) );
  NAND2_X1 U425 ( .A1(n367), .A2(n366), .ZN(n369) );
  XOR2_X1 U426 ( .A(KEYINPUT47), .B(KEYINPUT110), .Z(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  NAND2_X1 U428 ( .A1(n370), .A2(n371), .ZN(n373) );
  XOR2_X1 U429 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n375) );
  XNOR2_X1 U430 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U432 ( .A(KEYINPUT18), .B(n376), .Z(n452) );
  XOR2_X1 U433 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n378) );
  XNOR2_X1 U434 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U436 ( .A(G197GAT), .B(n379), .Z(n433) );
  XNOR2_X1 U437 ( .A(n452), .B(n433), .ZN(n392) );
  XOR2_X1 U438 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n381) );
  XNOR2_X1 U439 ( .A(G204GAT), .B(G92GAT), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n386) );
  XOR2_X1 U441 ( .A(n382), .B(KEYINPUT93), .Z(n384) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U444 ( .A(n386), .B(n385), .Z(n390) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U447 ( .A(n392), .B(n391), .Z(n511) );
  INV_X1 U448 ( .A(n511), .ZN(n523) );
  NAND2_X1 U449 ( .A1(n533), .A2(n523), .ZN(n394) );
  XOR2_X1 U450 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n393) );
  XNOR2_X1 U451 ( .A(n394), .B(n393), .ZN(n415) );
  XOR2_X1 U452 ( .A(KEYINPUT0), .B(G134GAT), .Z(n396) );
  XNOR2_X1 U453 ( .A(KEYINPUT80), .B(G127GAT), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U455 ( .A(G113GAT), .B(n397), .ZN(n446) );
  XOR2_X1 U456 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n399) );
  XNOR2_X1 U457 ( .A(KEYINPUT6), .B(KEYINPUT91), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n413) );
  XOR2_X1 U459 ( .A(G148GAT), .B(G120GAT), .Z(n401) );
  XNOR2_X1 U460 ( .A(G29GAT), .B(G141GAT), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U462 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n403) );
  XNOR2_X1 U463 ( .A(G1GAT), .B(G57GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U465 ( .A(n405), .B(n404), .Z(n411) );
  XNOR2_X1 U466 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n406), .B(KEYINPUT3), .ZN(n421) );
  XOR2_X1 U468 ( .A(G85GAT), .B(G162GAT), .Z(n408) );
  NAND2_X1 U469 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n421), .B(n409), .ZN(n410) );
  XNOR2_X1 U472 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U473 ( .A(n413), .B(n412), .Z(n414) );
  XOR2_X1 U474 ( .A(n446), .B(n414), .Z(n550) );
  INV_X1 U475 ( .A(n550), .ZN(n521) );
  XOR2_X1 U476 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n418) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U478 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U479 ( .A(n419), .B(KEYINPUT23), .Z(n423) );
  XNOR2_X1 U480 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n425) );
  XNOR2_X1 U483 ( .A(G218GAT), .B(G106GAT), .ZN(n424) );
  XNOR2_X1 U484 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U485 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n468) );
  NAND2_X1 U489 ( .A1(n293), .A2(n468), .ZN(n435) );
  XOR2_X1 U490 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n453) );
  XOR2_X1 U492 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT84), .B(KEYINPUT83), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U495 ( .A(KEYINPUT81), .B(G15GAT), .Z(n439) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G43GAT), .ZN(n438) );
  XNOR2_X1 U497 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n450) );
  XOR2_X1 U499 ( .A(G99GAT), .B(G190GAT), .Z(n444) );
  XNOR2_X1 U500 ( .A(n442), .B(G176GAT), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U502 ( .A(n446), .B(n445), .ZN(n448) );
  NAND2_X1 U503 ( .A1(G227GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XOR2_X1 U506 ( .A(n452), .B(n451), .Z(n527) );
  INV_X1 U507 ( .A(n527), .ZN(n536) );
  NOR2_X1 U508 ( .A1(n453), .A2(n536), .ZN(n454) );
  XNOR2_X1 U509 ( .A(n454), .B(KEYINPUT119), .ZN(n568) );
  NOR2_X1 U510 ( .A1(n568), .A2(n545), .ZN(n458) );
  XNOR2_X1 U511 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n456) );
  INV_X1 U512 ( .A(G190GAT), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n573), .A2(n568), .ZN(n461) );
  INV_X1 U514 ( .A(KEYINPUT120), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n459), .B(G169GAT), .ZN(n460) );
  XNOR2_X1 U516 ( .A(n461), .B(n460), .ZN(G1348GAT) );
  NOR2_X1 U517 ( .A1(n573), .A2(n579), .ZN(n462) );
  XOR2_X1 U518 ( .A(KEYINPUT71), .B(n462), .Z(n492) );
  XOR2_X1 U519 ( .A(n511), .B(KEYINPUT95), .Z(n463) );
  XOR2_X1 U520 ( .A(n463), .B(KEYINPUT27), .Z(n470) );
  INV_X1 U521 ( .A(n470), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT28), .B(n468), .Z(n529) );
  INV_X1 U523 ( .A(n529), .ZN(n515) );
  NAND2_X1 U524 ( .A1(n521), .A2(n515), .ZN(n464) );
  NOR2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n534) );
  NAND2_X1 U526 ( .A1(n534), .A2(n536), .ZN(n474) );
  NAND2_X1 U527 ( .A1(n527), .A2(n523), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n468), .A2(n466), .ZN(n467) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n467), .Z(n471) );
  NOR2_X1 U530 ( .A1(n468), .A2(n527), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n469), .B(KEYINPUT26), .ZN(n571) );
  NAND2_X1 U532 ( .A1(n571), .A2(n470), .ZN(n549) );
  NAND2_X1 U533 ( .A1(n471), .A2(n549), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n550), .A2(n472), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n474), .A2(n473), .ZN(n488) );
  NAND2_X1 U536 ( .A1(n475), .A2(n545), .ZN(n476) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n476), .Z(n477) );
  AND2_X1 U538 ( .A1(n488), .A2(n477), .ZN(n508) );
  NAND2_X1 U539 ( .A1(n492), .A2(n508), .ZN(n478) );
  XNOR2_X1 U540 ( .A(KEYINPUT96), .B(n478), .ZN(n486) );
  NOR2_X1 U541 ( .A1(n486), .A2(n550), .ZN(n480) );
  XNOR2_X1 U542 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U545 ( .A1(n486), .A2(n511), .ZN(n482) );
  XOR2_X1 U546 ( .A(G8GAT), .B(n482), .Z(n483) );
  XNOR2_X1 U547 ( .A(KEYINPUT98), .B(n483), .ZN(G1325GAT) );
  NOR2_X1 U548 ( .A1(n486), .A2(n536), .ZN(n485) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n484) );
  XNOR2_X1 U550 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  NOR2_X1 U551 ( .A1(n515), .A2(n486), .ZN(n487) );
  XOR2_X1 U552 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NAND2_X1 U554 ( .A1(n583), .A2(n488), .ZN(n489) );
  NOR2_X1 U555 ( .A1(n586), .A2(n489), .ZN(n491) );
  XNOR2_X1 U556 ( .A(KEYINPUT37), .B(KEYINPUT99), .ZN(n490) );
  XNOR2_X1 U557 ( .A(n491), .B(n490), .ZN(n518) );
  NAND2_X1 U558 ( .A1(n518), .A2(n492), .ZN(n493) );
  XOR2_X1 U559 ( .A(KEYINPUT38), .B(n493), .Z(n502) );
  NAND2_X1 U560 ( .A1(n521), .A2(n502), .ZN(n494) );
  XNOR2_X1 U561 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n502), .A2(n523), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n496), .B(KEYINPUT100), .ZN(n497) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n497), .ZN(G1329GAT) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n501) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT40), .Z(n499) );
  NAND2_X1 U567 ( .A1(n527), .A2(n502), .ZN(n498) );
  XNOR2_X1 U568 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n501), .B(n500), .ZN(G1330GAT) );
  XOR2_X1 U570 ( .A(G50GAT), .B(KEYINPUT103), .Z(n504) );
  NAND2_X1 U571 ( .A1(n502), .A2(n529), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U575 ( .A(n506), .B(n505), .ZN(n510) );
  NOR2_X1 U576 ( .A1(n562), .A2(n507), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n519), .A2(n508), .ZN(n514) );
  NOR2_X1 U578 ( .A1(n550), .A2(n514), .ZN(n509) );
  XOR2_X1 U579 ( .A(n510), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U580 ( .A1(n511), .A2(n514), .ZN(n512) );
  XOR2_X1 U581 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U582 ( .A1(n536), .A2(n514), .ZN(n513) );
  XOR2_X1 U583 ( .A(G71GAT), .B(n513), .Z(G1334GAT) );
  NOR2_X1 U584 ( .A1(n515), .A2(n514), .ZN(n517) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U586 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U587 ( .A1(n519), .A2(n518), .ZN(n520) );
  XOR2_X1 U588 ( .A(KEYINPUT106), .B(n520), .Z(n530) );
  NAND2_X1 U589 ( .A1(n530), .A2(n521), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n525) );
  NAND2_X1 U592 ( .A1(n523), .A2(n530), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(G92GAT), .B(n526), .ZN(G1337GAT) );
  NAND2_X1 U595 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U596 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n531), .B(KEYINPUT44), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U600 ( .A1(n534), .A2(n551), .ZN(n535) );
  NOR2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT113), .B(n537), .ZN(n544) );
  NOR2_X1 U603 ( .A1(n573), .A2(n544), .ZN(n538) );
  XOR2_X1 U604 ( .A(G113GAT), .B(n538), .Z(G1340GAT) );
  NOR2_X1 U605 ( .A1(n562), .A2(n544), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  NOR2_X1 U608 ( .A1(n583), .A2(n544), .ZN(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT114), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U611 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U613 ( .A(KEYINPUT115), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NOR2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n552) );
  NAND2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n559) );
  NOR2_X1 U618 ( .A1(n573), .A2(n559), .ZN(n553) );
  XOR2_X1 U619 ( .A(G141GAT), .B(n553), .Z(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n555) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n562), .A2(n559), .ZN(n556) );
  XOR2_X1 U624 ( .A(n557), .B(n556), .Z(G1345GAT) );
  NOR2_X1 U625 ( .A1(n583), .A2(n559), .ZN(n558) );
  XOR2_X1 U626 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n568), .ZN(n567) );
  XOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n564) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U633 ( .A(KEYINPUT121), .B(n565), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n583), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(KEYINPUT123), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n571), .A2(n293), .ZN(n572) );
  INV_X1 U639 ( .A(n580), .ZN(n585) );
  NOR2_X1 U640 ( .A1(n573), .A2(n585), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n575) );
  XNOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n574) );
  XNOR2_X1 U643 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U644 ( .A(KEYINPUT59), .B(n576), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .Z(n582) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n583), .A2(n585), .ZN(n584) );
  XOR2_X1 U650 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

