

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U548 ( .A1(n615), .A2(n616), .ZN(n630) );
  NOR2_X1 U549 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U550 ( .A1(G651), .A2(n575), .ZN(n797) );
  NOR2_X1 U551 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U552 ( .A1(n793), .A2(G85), .ZN(n512) );
  XNOR2_X1 U553 ( .A(n512), .B(KEYINPUT68), .ZN(n514) );
  XOR2_X1 U554 ( .A(KEYINPUT0), .B(G543), .Z(n575) );
  INV_X1 U555 ( .A(G651), .ZN(n516) );
  NOR2_X1 U556 ( .A1(n575), .A2(n516), .ZN(n789) );
  NAND2_X1 U557 ( .A1(G72), .A2(n789), .ZN(n513) );
  NAND2_X1 U558 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U559 ( .A(KEYINPUT69), .B(n515), .ZN(n521) );
  NOR2_X1 U560 ( .A1(G543), .A2(n516), .ZN(n517) );
  XOR2_X1 U561 ( .A(KEYINPUT1), .B(n517), .Z(n790) );
  NAND2_X1 U562 ( .A1(G60), .A2(n790), .ZN(n519) );
  NAND2_X1 U563 ( .A1(G47), .A2(n797), .ZN(n518) );
  AND2_X1 U564 ( .A1(n519), .A2(n518), .ZN(n520) );
  NAND2_X1 U565 ( .A1(n521), .A2(n520), .ZN(G290) );
  AND2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U567 ( .A1(G114), .A2(n881), .ZN(n522) );
  XOR2_X1 U568 ( .A(KEYINPUT84), .B(n522), .Z(n525) );
  INV_X1 U569 ( .A(G2104), .ZN(n530) );
  AND2_X1 U570 ( .A1(n530), .A2(G2105), .ZN(n883) );
  NAND2_X1 U571 ( .A1(G126), .A2(n883), .ZN(n523) );
  XNOR2_X1 U572 ( .A(KEYINPUT83), .B(n523), .ZN(n524) );
  NOR2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n529) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X1 U575 ( .A(KEYINPUT17), .B(n526), .Z(n527) );
  XNOR2_X2 U576 ( .A(KEYINPUT66), .B(n527), .ZN(n877) );
  NAND2_X1 U577 ( .A1(G138), .A2(n877), .ZN(n528) );
  NAND2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n533) );
  NOR2_X1 U579 ( .A1(G2105), .A2(n530), .ZN(n876) );
  NAND2_X1 U580 ( .A1(G102), .A2(n876), .ZN(n531) );
  XNOR2_X1 U581 ( .A(KEYINPUT85), .B(n531), .ZN(n532) );
  NOR2_X1 U582 ( .A1(n533), .A2(n532), .ZN(G164) );
  NAND2_X1 U583 ( .A1(G113), .A2(n881), .ZN(n535) );
  NAND2_X1 U584 ( .A1(G125), .A2(n883), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n535), .A2(n534), .ZN(n538) );
  NAND2_X1 U586 ( .A1(G137), .A2(n877), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n536), .B(KEYINPUT67), .ZN(n537) );
  NOR2_X1 U588 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U589 ( .A1(n876), .A2(G101), .ZN(n540) );
  XNOR2_X1 U590 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n539) );
  XNOR2_X1 U591 ( .A(n540), .B(n539), .ZN(n541) );
  NAND2_X1 U592 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X2 U593 ( .A(n543), .B(KEYINPUT64), .Z(G160) );
  NAND2_X1 U594 ( .A1(G64), .A2(n790), .ZN(n545) );
  NAND2_X1 U595 ( .A1(G52), .A2(n797), .ZN(n544) );
  NAND2_X1 U596 ( .A1(n545), .A2(n544), .ZN(n550) );
  NAND2_X1 U597 ( .A1(G90), .A2(n793), .ZN(n547) );
  NAND2_X1 U598 ( .A1(G77), .A2(n789), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n548), .Z(n549) );
  NOR2_X1 U601 ( .A1(n550), .A2(n549), .ZN(G171) );
  NAND2_X1 U602 ( .A1(G91), .A2(n793), .ZN(n552) );
  NAND2_X1 U603 ( .A1(G78), .A2(n789), .ZN(n551) );
  NAND2_X1 U604 ( .A1(n552), .A2(n551), .ZN(n555) );
  NAND2_X1 U605 ( .A1(n797), .A2(G53), .ZN(n553) );
  XOR2_X1 U606 ( .A(KEYINPUT70), .B(n553), .Z(n554) );
  NOR2_X1 U607 ( .A1(n555), .A2(n554), .ZN(n557) );
  NAND2_X1 U608 ( .A1(n790), .A2(G65), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n557), .A2(n556), .ZN(G299) );
  NAND2_X1 U610 ( .A1(G89), .A2(n793), .ZN(n558) );
  XOR2_X1 U611 ( .A(KEYINPUT75), .B(n558), .Z(n559) );
  XNOR2_X1 U612 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G76), .A2(n789), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U615 ( .A(n562), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U616 ( .A1(G63), .A2(n790), .ZN(n564) );
  NAND2_X1 U617 ( .A1(G51), .A2(n797), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U619 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U620 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U621 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U622 ( .A1(G88), .A2(n793), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G75), .A2(n789), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U625 ( .A1(G62), .A2(n790), .ZN(n572) );
  NAND2_X1 U626 ( .A1(G50), .A2(n797), .ZN(n571) );
  NAND2_X1 U627 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U628 ( .A1(n574), .A2(n573), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  XOR2_X1 U630 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U631 ( .A1(n575), .A2(G87), .ZN(n576) );
  XNOR2_X1 U632 ( .A(KEYINPUT80), .B(n576), .ZN(n582) );
  NAND2_X1 U633 ( .A1(G49), .A2(n797), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G74), .A2(G651), .ZN(n577) );
  NAND2_X1 U635 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U636 ( .A1(n790), .A2(n579), .ZN(n580) );
  XOR2_X1 U637 ( .A(KEYINPUT79), .B(n580), .Z(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U639 ( .A1(G86), .A2(n793), .ZN(n584) );
  NAND2_X1 U640 ( .A1(G61), .A2(n790), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U642 ( .A1(n789), .A2(G73), .ZN(n585) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n585), .Z(n586) );
  NOR2_X1 U644 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U645 ( .A(KEYINPUT81), .B(n588), .Z(n590) );
  NAND2_X1 U646 ( .A1(n797), .A2(G48), .ZN(n589) );
  NAND2_X1 U647 ( .A1(n590), .A2(n589), .ZN(G305) );
  XOR2_X1 U648 ( .A(G1986), .B(G290), .Z(n970) );
  INV_X1 U649 ( .A(n970), .ZN(n591) );
  NOR2_X1 U650 ( .A1(G164), .A2(G1384), .ZN(n592) );
  NAND2_X1 U651 ( .A1(G40), .A2(G160), .ZN(n616) );
  NOR2_X1 U652 ( .A1(n592), .A2(n616), .ZN(n746) );
  NAND2_X1 U653 ( .A1(n591), .A2(n746), .ZN(n736) );
  INV_X1 U654 ( .A(G2084), .ZN(n593) );
  INV_X1 U655 ( .A(n592), .ZN(n615) );
  AND2_X1 U656 ( .A1(n593), .A2(n630), .ZN(n645) );
  NAND2_X1 U657 ( .A1(G8), .A2(n645), .ZN(n656) );
  OR2_X1 U658 ( .A1(n615), .A2(n616), .ZN(n596) );
  INV_X1 U659 ( .A(G8), .ZN(n594) );
  NOR2_X1 U660 ( .A1(n594), .A2(G1966), .ZN(n595) );
  AND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n654) );
  NOR2_X1 U662 ( .A1(n630), .A2(G1961), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n597), .B(KEYINPUT97), .ZN(n599) );
  XNOR2_X1 U664 ( .A(G2078), .B(KEYINPUT25), .ZN(n937) );
  NAND2_X1 U665 ( .A1(n630), .A2(n937), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n649) );
  NAND2_X1 U667 ( .A1(n649), .A2(G171), .ZN(n644) );
  INV_X1 U668 ( .A(G299), .ZN(n962) );
  NAND2_X1 U669 ( .A1(n630), .A2(G2072), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT27), .ZN(n602) );
  INV_X1 U671 ( .A(G1956), .ZN(n963) );
  NOR2_X1 U672 ( .A1(n963), .A2(n630), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n962), .A2(n605), .ZN(n604) );
  INV_X1 U675 ( .A(KEYINPUT28), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n604), .B(n603), .ZN(n641) );
  NAND2_X1 U677 ( .A1(n962), .A2(n605), .ZN(n639) );
  NAND2_X1 U678 ( .A1(G56), .A2(n790), .ZN(n606) );
  XOR2_X1 U679 ( .A(KEYINPUT14), .B(n606), .Z(n612) );
  NAND2_X1 U680 ( .A1(n793), .A2(G81), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT12), .ZN(n609) );
  NAND2_X1 U682 ( .A1(G68), .A2(n789), .ZN(n608) );
  NAND2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U684 ( .A(KEYINPUT13), .B(n610), .Z(n611) );
  NOR2_X1 U685 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n797), .A2(G43), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n966) );
  INV_X1 U688 ( .A(G1996), .ZN(n835) );
  OR2_X1 U689 ( .A1(n615), .A2(n835), .ZN(n617) );
  NOR2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U691 ( .A(n618), .B(KEYINPUT26), .Z(n620) );
  NAND2_X1 U692 ( .A1(n596), .A2(G1341), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n966), .A2(n621), .ZN(n634) );
  NAND2_X1 U695 ( .A1(G79), .A2(n789), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G54), .A2(n797), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n623), .A2(n622), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G92), .A2(n793), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G66), .A2(n790), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U701 ( .A(KEYINPUT74), .B(n626), .ZN(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U703 ( .A(n629), .B(KEYINPUT15), .Z(n971) );
  INV_X1 U704 ( .A(n971), .ZN(n768) );
  NAND2_X1 U705 ( .A1(G1348), .A2(n596), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G2067), .A2(n630), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n635) );
  NOR2_X1 U708 ( .A1(n768), .A2(n635), .ZN(n633) );
  OR2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U710 ( .A1(n768), .A2(n635), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U714 ( .A(n642), .B(KEYINPUT29), .Z(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n662) );
  NOR2_X1 U716 ( .A1(n654), .A2(n645), .ZN(n646) );
  NAND2_X1 U717 ( .A1(n646), .A2(G8), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n647), .B(KEYINPUT30), .ZN(n648) );
  NOR2_X1 U719 ( .A1(G168), .A2(n648), .ZN(n651) );
  NOR2_X1 U720 ( .A1(G171), .A2(n649), .ZN(n650) );
  XOR2_X1 U721 ( .A(KEYINPUT31), .B(n652), .Z(n661) );
  AND2_X1 U722 ( .A1(n662), .A2(n661), .ZN(n653) );
  NOR2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n670) );
  NAND2_X1 U725 ( .A1(G8), .A2(n596), .ZN(n727) );
  NOR2_X1 U726 ( .A1(G1971), .A2(n727), .ZN(n658) );
  NOR2_X1 U727 ( .A1(G2090), .A2(n596), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n659), .A2(G303), .ZN(n660) );
  OR2_X1 U730 ( .A1(n594), .A2(n660), .ZN(n664) );
  AND2_X1 U731 ( .A1(n661), .A2(n664), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n667) );
  INV_X1 U733 ( .A(n664), .ZN(n665) );
  OR2_X1 U734 ( .A1(n665), .A2(G286), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n668), .B(KEYINPUT32), .ZN(n669) );
  NAND2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT98), .B(n671), .ZN(n725) );
  NOR2_X1 U739 ( .A1(G1976), .A2(G288), .ZN(n674) );
  NOR2_X1 U740 ( .A1(G1971), .A2(G303), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n674), .A2(n672), .ZN(n969) );
  INV_X1 U742 ( .A(n727), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n675), .A2(KEYINPUT33), .ZN(n677) );
  AND2_X1 U745 ( .A1(n969), .A2(n677), .ZN(n676) );
  NAND2_X1 U746 ( .A1(n725), .A2(n676), .ZN(n682) );
  INV_X1 U747 ( .A(n677), .ZN(n680) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n960) );
  NOR2_X1 U749 ( .A1(n727), .A2(KEYINPUT33), .ZN(n678) );
  AND2_X1 U750 ( .A1(n960), .A2(n678), .ZN(n679) );
  OR2_X1 U751 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U753 ( .A(KEYINPUT99), .B(n683), .Z(n720) );
  XOR2_X1 U754 ( .A(G1981), .B(G305), .Z(n979) );
  NAND2_X1 U755 ( .A1(G95), .A2(n876), .ZN(n684) );
  XNOR2_X1 U756 ( .A(n684), .B(KEYINPUT88), .ZN(n691) );
  NAND2_X1 U757 ( .A1(G107), .A2(n881), .ZN(n686) );
  NAND2_X1 U758 ( .A1(G119), .A2(n883), .ZN(n685) );
  NAND2_X1 U759 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U760 ( .A1(G131), .A2(n877), .ZN(n687) );
  XNOR2_X1 U761 ( .A(KEYINPUT89), .B(n687), .ZN(n688) );
  NOR2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U763 ( .A1(n691), .A2(n690), .ZN(n870) );
  NAND2_X1 U764 ( .A1(G1991), .A2(n870), .ZN(n692) );
  XNOR2_X1 U765 ( .A(n692), .B(KEYINPUT90), .ZN(n703) );
  NAND2_X1 U766 ( .A1(G117), .A2(n881), .ZN(n694) );
  NAND2_X1 U767 ( .A1(G129), .A2(n883), .ZN(n693) );
  NAND2_X1 U768 ( .A1(n694), .A2(n693), .ZN(n698) );
  NAND2_X1 U769 ( .A1(G105), .A2(n876), .ZN(n695) );
  XNOR2_X1 U770 ( .A(n695), .B(KEYINPUT38), .ZN(n696) );
  XNOR2_X1 U771 ( .A(n696), .B(KEYINPUT91), .ZN(n697) );
  NOR2_X1 U772 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n699), .B(KEYINPUT92), .ZN(n701) );
  NAND2_X1 U774 ( .A1(G141), .A2(n877), .ZN(n700) );
  NAND2_X1 U775 ( .A1(n701), .A2(n700), .ZN(n895) );
  NAND2_X1 U776 ( .A1(G1996), .A2(n895), .ZN(n702) );
  NAND2_X1 U777 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U778 ( .A(KEYINPUT93), .B(n704), .Z(n932) );
  NAND2_X1 U779 ( .A1(n932), .A2(n746), .ZN(n705) );
  XOR2_X1 U780 ( .A(KEYINPUT94), .B(n705), .Z(n739) );
  XNOR2_X1 U781 ( .A(KEYINPUT95), .B(n739), .ZN(n717) );
  XNOR2_X1 U782 ( .A(KEYINPUT87), .B(KEYINPUT36), .ZN(n716) );
  NAND2_X1 U783 ( .A1(G116), .A2(n881), .ZN(n707) );
  NAND2_X1 U784 ( .A1(G128), .A2(n883), .ZN(n706) );
  NAND2_X1 U785 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U786 ( .A(KEYINPUT35), .B(n708), .ZN(n714) );
  NAND2_X1 U787 ( .A1(G104), .A2(n876), .ZN(n710) );
  NAND2_X1 U788 ( .A1(G140), .A2(n877), .ZN(n709) );
  NAND2_X1 U789 ( .A1(n710), .A2(n709), .ZN(n712) );
  XOR2_X1 U790 ( .A(KEYINPUT86), .B(KEYINPUT34), .Z(n711) );
  XNOR2_X1 U791 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U792 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U793 ( .A(n716), .B(n715), .ZN(n896) );
  XNOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NOR2_X1 U795 ( .A1(n896), .A2(n744), .ZN(n911) );
  NAND2_X1 U796 ( .A1(n746), .A2(n911), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n717), .A2(n742), .ZN(n732) );
  INV_X1 U798 ( .A(n732), .ZN(n718) );
  AND2_X1 U799 ( .A1(n979), .A2(n718), .ZN(n719) );
  NAND2_X1 U800 ( .A1(n720), .A2(n719), .ZN(n734) );
  NOR2_X1 U801 ( .A1(G1981), .A2(G305), .ZN(n721) );
  XOR2_X1 U802 ( .A(n721), .B(KEYINPUT24), .Z(n722) );
  XNOR2_X1 U803 ( .A(KEYINPUT96), .B(n722), .ZN(n723) );
  OR2_X1 U804 ( .A1(n727), .A2(n723), .ZN(n730) );
  NOR2_X1 U805 ( .A1(G2090), .A2(G303), .ZN(n724) );
  NAND2_X1 U806 ( .A1(G8), .A2(n724), .ZN(n726) );
  NAND2_X1 U807 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U808 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U809 ( .A1(n730), .A2(n729), .ZN(n731) );
  OR2_X1 U810 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U811 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U812 ( .A1(n736), .A2(n735), .ZN(n749) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n895), .ZN(n919) );
  NOR2_X1 U814 ( .A1(G1991), .A2(n870), .ZN(n924) );
  NOR2_X1 U815 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U816 ( .A1(n924), .A2(n737), .ZN(n738) );
  NOR2_X1 U817 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U818 ( .A1(n919), .A2(n740), .ZN(n741) );
  XNOR2_X1 U819 ( .A(n741), .B(KEYINPUT39), .ZN(n743) );
  NAND2_X1 U820 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U821 ( .A1(n896), .A2(n744), .ZN(n910) );
  NAND2_X1 U822 ( .A1(n745), .A2(n910), .ZN(n747) );
  NAND2_X1 U823 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n751) );
  XNOR2_X1 U825 ( .A(KEYINPUT100), .B(KEYINPUT40), .ZN(n750) );
  XNOR2_X1 U826 ( .A(n751), .B(n750), .ZN(G329) );
  INV_X1 U827 ( .A(G171), .ZN(G301) );
  XOR2_X1 U828 ( .A(KEYINPUT103), .B(G2454), .Z(n753) );
  XNOR2_X1 U829 ( .A(KEYINPUT102), .B(G2430), .ZN(n752) );
  XNOR2_X1 U830 ( .A(n753), .B(n752), .ZN(n763) );
  XOR2_X1 U831 ( .A(G2446), .B(G2451), .Z(n755) );
  XNOR2_X1 U832 ( .A(G1341), .B(G2435), .ZN(n754) );
  XNOR2_X1 U833 ( .A(n755), .B(n754), .ZN(n759) );
  XOR2_X1 U834 ( .A(G2438), .B(G2427), .Z(n757) );
  XNOR2_X1 U835 ( .A(KEYINPUT101), .B(KEYINPUT104), .ZN(n756) );
  XNOR2_X1 U836 ( .A(n757), .B(n756), .ZN(n758) );
  XOR2_X1 U837 ( .A(n759), .B(n758), .Z(n761) );
  XNOR2_X1 U838 ( .A(G1348), .B(G2443), .ZN(n760) );
  XNOR2_X1 U839 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U840 ( .A(n763), .B(n762), .ZN(n764) );
  AND2_X1 U841 ( .A1(n764), .A2(G14), .ZN(G401) );
  AND2_X1 U842 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  INV_X1 U844 ( .A(G82), .ZN(G220) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U846 ( .A(n765), .B(KEYINPUT72), .ZN(n766) );
  XOR2_X1 U847 ( .A(KEYINPUT10), .B(n766), .Z(n826) );
  NAND2_X1 U848 ( .A1(n826), .A2(G567), .ZN(n767) );
  XOR2_X1 U849 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  XNOR2_X1 U850 ( .A(G860), .B(KEYINPUT73), .ZN(n774) );
  OR2_X1 U851 ( .A1(n966), .A2(n774), .ZN(G153) );
  NAND2_X1 U852 ( .A1(G868), .A2(G301), .ZN(n770) );
  INV_X1 U853 ( .A(G868), .ZN(n810) );
  NAND2_X1 U854 ( .A1(n768), .A2(n810), .ZN(n769) );
  NAND2_X1 U855 ( .A1(n770), .A2(n769), .ZN(G284) );
  NOR2_X1 U856 ( .A1(G286), .A2(n810), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT76), .ZN(n773) );
  NOR2_X1 U858 ( .A1(G299), .A2(G868), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U860 ( .A1(n774), .A2(G559), .ZN(n775) );
  NAND2_X1 U861 ( .A1(n775), .A2(n971), .ZN(n776) );
  XNOR2_X1 U862 ( .A(n776), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U863 ( .A1(G868), .A2(n966), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G868), .A2(n971), .ZN(n777) );
  NOR2_X1 U865 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U866 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U867 ( .A1(G123), .A2(n883), .ZN(n780) );
  XOR2_X1 U868 ( .A(KEYINPUT77), .B(n780), .Z(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G111), .A2(n881), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n787) );
  NAND2_X1 U872 ( .A1(G99), .A2(n876), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G135), .A2(n877), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n923) );
  XNOR2_X1 U876 ( .A(n923), .B(G2096), .ZN(n788) );
  INV_X1 U877 ( .A(G2100), .ZN(n844) );
  NAND2_X1 U878 ( .A1(n788), .A2(n844), .ZN(G156) );
  NAND2_X1 U879 ( .A1(G80), .A2(n789), .ZN(n792) );
  NAND2_X1 U880 ( .A1(G67), .A2(n790), .ZN(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U882 ( .A1(n793), .A2(G93), .ZN(n794) );
  XOR2_X1 U883 ( .A(KEYINPUT78), .B(n794), .Z(n795) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U885 ( .A1(n797), .A2(G55), .ZN(n798) );
  NAND2_X1 U886 ( .A1(n799), .A2(n798), .ZN(n811) );
  NAND2_X1 U887 ( .A1(G559), .A2(n971), .ZN(n800) );
  XNOR2_X1 U888 ( .A(n966), .B(n800), .ZN(n808) );
  NOR2_X1 U889 ( .A1(G860), .A2(n808), .ZN(n801) );
  XOR2_X1 U890 ( .A(n811), .B(n801), .Z(G145) );
  XOR2_X1 U891 ( .A(KEYINPUT82), .B(KEYINPUT19), .Z(n802) );
  XNOR2_X1 U892 ( .A(G288), .B(n802), .ZN(n805) );
  XOR2_X1 U893 ( .A(G299), .B(G305), .Z(n803) );
  XNOR2_X1 U894 ( .A(n803), .B(n811), .ZN(n804) );
  XNOR2_X1 U895 ( .A(n805), .B(n804), .ZN(n807) );
  XOR2_X1 U896 ( .A(G290), .B(G303), .Z(n806) );
  XNOR2_X1 U897 ( .A(n807), .B(n806), .ZN(n899) );
  XNOR2_X1 U898 ( .A(n899), .B(n808), .ZN(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n813) );
  NOR2_X1 U900 ( .A1(G868), .A2(n811), .ZN(n812) );
  NOR2_X1 U901 ( .A1(n813), .A2(n812), .ZN(G295) );
  NAND2_X1 U902 ( .A1(G2078), .A2(G2084), .ZN(n814) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n814), .Z(n815) );
  NAND2_X1 U904 ( .A1(G2090), .A2(n815), .ZN(n816) );
  XNOR2_X1 U905 ( .A(KEYINPUT21), .B(n816), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n817), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U907 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U908 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U909 ( .A1(G120), .A2(G108), .ZN(n818) );
  NOR2_X1 U910 ( .A1(G237), .A2(n818), .ZN(n819) );
  NAND2_X1 U911 ( .A1(G69), .A2(n819), .ZN(n1019) );
  NAND2_X1 U912 ( .A1(n1019), .A2(G567), .ZN(n824) );
  NOR2_X1 U913 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U914 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U915 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G96), .A2(n822), .ZN(n1020) );
  NAND2_X1 U917 ( .A1(n1020), .A2(G2106), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(n831) );
  NAND2_X1 U919 ( .A1(G483), .A2(G661), .ZN(n825) );
  NOR2_X1 U920 ( .A1(n831), .A2(n825), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(G36), .ZN(G176) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n826), .ZN(G217) );
  INV_X1 U923 ( .A(n826), .ZN(G223) );
  AND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n827) );
  NAND2_X1 U925 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U926 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(n830), .Z(G188) );
  INV_X1 U929 ( .A(n831), .ZN(G319) );
  XOR2_X1 U930 ( .A(KEYINPUT107), .B(G2474), .Z(n833) );
  XOR2_X1 U931 ( .A(n963), .B(KEYINPUT41), .Z(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(n834), .B(G1961), .Z(n837) );
  XOR2_X1 U934 ( .A(n835), .B(G1991), .Z(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U936 ( .A(G1976), .B(G1981), .Z(n839) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1966), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1971), .B(KEYINPUT108), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(G229) );
  XNOR2_X1 U942 ( .A(n844), .B(G2096), .ZN(n846) );
  XNOR2_X1 U943 ( .A(G2090), .B(KEYINPUT43), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U945 ( .A(n847), .B(G2678), .Z(n849) );
  XNOR2_X1 U946 ( .A(G2072), .B(KEYINPUT42), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U948 ( .A(KEYINPUT106), .B(G2084), .Z(n851) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2078), .ZN(n850) );
  XNOR2_X1 U950 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(G227) );
  NAND2_X1 U952 ( .A1(G124), .A2(n883), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U954 ( .A1(n881), .A2(G112), .ZN(n855) );
  NAND2_X1 U955 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U956 ( .A1(G100), .A2(n876), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G136), .A2(n877), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U959 ( .A1(n860), .A2(n859), .ZN(G162) );
  NAND2_X1 U960 ( .A1(n883), .A2(G127), .ZN(n861) );
  XOR2_X1 U961 ( .A(KEYINPUT113), .B(n861), .Z(n863) );
  NAND2_X1 U962 ( .A1(n881), .A2(G115), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(KEYINPUT47), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G103), .A2(n876), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n877), .A2(G139), .ZN(n867) );
  XOR2_X1 U968 ( .A(KEYINPUT112), .B(n867), .Z(n868) );
  NOR2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n913) );
  XNOR2_X1 U970 ( .A(G162), .B(G160), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(n870), .ZN(n875) );
  XOR2_X1 U972 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n873) );
  XNOR2_X1 U973 ( .A(KEYINPUT114), .B(KEYINPUT111), .ZN(n872) );
  XNOR2_X1 U974 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U975 ( .A(n875), .B(n874), .Z(n892) );
  NAND2_X1 U976 ( .A1(G106), .A2(n876), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G142), .A2(n877), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(n880), .B(KEYINPUT45), .ZN(n888) );
  NAND2_X1 U980 ( .A1(n881), .A2(G118), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT109), .B(n882), .Z(n885) );
  NAND2_X1 U982 ( .A1(n883), .A2(G130), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U984 ( .A(KEYINPUT110), .B(n886), .Z(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n889), .B(n923), .ZN(n890) );
  XNOR2_X1 U987 ( .A(G164), .B(n890), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U989 ( .A(n913), .B(n893), .Z(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U993 ( .A(G286), .B(n899), .Z(n900) );
  XOR2_X1 U994 ( .A(n971), .B(n900), .Z(n902) );
  XNOR2_X1 U995 ( .A(n966), .B(G301), .ZN(n901) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U997 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n904), .B(KEYINPUT49), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G401), .A2(n905), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(G319), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT115), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n908) );
  NAND2_X1 U1004 ( .A1(n909), .A2(n908), .ZN(G225) );
  XOR2_X1 U1005 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  XNOR2_X1 U1006 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  INV_X1 U1008 ( .A(n910), .ZN(n912) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n930) );
  XNOR2_X1 U1010 ( .A(G164), .B(G2078), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(G2072), .B(n913), .ZN(n914) );
  XNOR2_X1 U1012 ( .A(n914), .B(KEYINPUT118), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n917), .B(KEYINPUT50), .ZN(n928) );
  XOR2_X1 U1015 ( .A(G160), .B(G2084), .Z(n922) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(KEYINPUT51), .B(n920), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n926) );
  NOR2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(KEYINPUT52), .B(n933), .ZN(n935) );
  INV_X1 U1026 ( .A(KEYINPUT55), .ZN(n934) );
  NAND2_X1 U1027 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1028 ( .A1(n936), .A2(G29), .ZN(n1017) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G35), .ZN(n951) );
  XOR2_X1 U1030 ( .A(n937), .B(G27), .Z(n939) );
  XNOR2_X1 U1031 ( .A(G1996), .B(G32), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(KEYINPUT120), .B(n940), .ZN(n946) );
  XOR2_X1 U1034 ( .A(G1991), .B(G25), .Z(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(G28), .ZN(n944) );
  XOR2_X1 U1036 ( .A(KEYINPUT119), .B(G2067), .Z(n942) );
  XNOR2_X1 U1037 ( .A(G26), .B(n942), .ZN(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1040 ( .A(G33), .B(G2072), .ZN(n947) );
  NOR2_X1 U1041 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1042 ( .A(KEYINPUT53), .B(n949), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1044 ( .A(KEYINPUT121), .B(n952), .Z(n955) );
  XOR2_X1 U1045 ( .A(G34), .B(KEYINPUT54), .Z(n953) );
  XNOR2_X1 U1046 ( .A(G2084), .B(n953), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1048 ( .A(KEYINPUT55), .B(n956), .Z(n958) );
  INV_X1 U1049 ( .A(G29), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(G11), .A2(n959), .ZN(n1015) );
  INV_X1 U1052 ( .A(G16), .ZN(n1011) );
  XOR2_X1 U1053 ( .A(n1011), .B(KEYINPUT56), .Z(n985) );
  XOR2_X1 U1054 ( .A(G301), .B(G1961), .Z(n961) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n977) );
  XOR2_X1 U1056 ( .A(n963), .B(n962), .Z(n965) );
  NAND2_X1 U1057 ( .A1(G1971), .A2(G303), .ZN(n964) );
  NAND2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n968) );
  XNOR2_X1 U1059 ( .A(G1341), .B(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n975) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1062 ( .A(G1348), .B(n971), .Z(n972) );
  NOR2_X1 U1063 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1066 ( .A(KEYINPUT122), .B(n978), .ZN(n983) );
  XNOR2_X1 U1067 ( .A(G1966), .B(G168), .ZN(n980) );
  NAND2_X1 U1068 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1069 ( .A(KEYINPUT57), .B(n981), .ZN(n982) );
  NAND2_X1 U1070 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n1013) );
  XOR2_X1 U1072 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n1009) );
  XNOR2_X1 U1073 ( .A(KEYINPUT123), .B(G1966), .ZN(n986) );
  XNOR2_X1 U1074 ( .A(n986), .B(G21), .ZN(n998) );
  XOR2_X1 U1075 ( .A(G20), .B(G1956), .Z(n990) );
  XNOR2_X1 U1076 ( .A(G1341), .B(G19), .ZN(n988) );
  XNOR2_X1 U1077 ( .A(G6), .B(G1981), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1080 ( .A(KEYINPUT59), .B(G1348), .Z(n991) );
  XNOR2_X1 U1081 ( .A(G4), .B(n991), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT60), .B(n994), .Z(n996) );
  XNOR2_X1 U1084 ( .A(G1961), .B(G5), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n1006) );
  XNOR2_X1 U1087 ( .A(G1971), .B(G22), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G23), .B(G1976), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1090 ( .A(G1986), .B(KEYINPUT124), .Z(n1001) );
  XNOR2_X1 U1091 ( .A(G24), .B(n1001), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT58), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(n1007), .B(KEYINPUT61), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1099 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1100 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1101 ( .A(KEYINPUT62), .B(n1018), .Z(G311) );
  XNOR2_X1 U1102 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1103 ( .A(G120), .ZN(G236) );
  INV_X1 U1104 ( .A(G96), .ZN(G221) );
  INV_X1 U1105 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(G325) );
  INV_X1 U1107 ( .A(G325), .ZN(G261) );
endmodule

