//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:53 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n451, new_n452,
    new_n454, new_n457, new_n458, new_n459, new_n460, new_n461, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n862, new_n863, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT64), .Z(G173));
  XOR2_X1   g024(.A(KEYINPUT65), .B(KEYINPUT1), .Z(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  AND2_X1   g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(G223));
  NAND2_X1  g028(.A1(new_n452), .A2(G567), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G234));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(G217));
  NOR4_X1   g031(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT2), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR4_X1   g034(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  AOI22_X1  g038(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n461), .ZN(G319));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G125), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT68), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n477), .A2(new_n478), .A3(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n473), .A2(KEYINPUT69), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT69), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(KEYINPUT3), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G137), .A3(new_n472), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n480), .A2(new_n482), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G101), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n470), .A2(new_n479), .B1(new_n487), .B2(new_n469), .ZN(G160));
  NAND2_X1  g063(.A1(new_n483), .A2(new_n472), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n483), .A2(KEYINPUT70), .A3(new_n472), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n469), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT71), .Z(new_n495));
  OAI21_X1  g070(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G112), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G136), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT4), .A2(G138), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n483), .A2(new_n472), .A3(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n472), .A2(new_n474), .A3(G138), .A4(new_n469), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT4), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(G102), .A2(G2105), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n510), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n506), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT73), .B1(new_n514), .B2(G543), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT5), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(new_n518), .B1(new_n514), .B2(G543), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT6), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(KEYINPUT72), .A3(KEYINPUT6), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n525), .A2(new_n526), .B1(new_n524), .B2(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT74), .B(G88), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n527), .A2(G543), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n522), .A2(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n534));
  XOR2_X1   g109(.A(new_n534), .B(KEYINPUT75), .Z(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  INV_X1    g112(.A(G51), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(new_n527), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT76), .B(G89), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n537), .B1(new_n531), .B2(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n535), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n521), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(KEYINPUT77), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(KEYINPUT77), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n519), .A2(new_n527), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n527), .A2(G543), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT78), .B(G52), .ZN(new_n549));
  AOI22_X1  g124(.A1(G90), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n514), .A2(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n516), .B1(KEYINPUT5), .B2(new_n517), .ZN(new_n555));
  NOR3_X1   g130(.A1(new_n514), .A2(KEYINPUT73), .A3(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n553), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n521), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n561), .B1(new_n560), .B2(new_n559), .ZN(new_n562));
  XOR2_X1   g137(.A(KEYINPUT80), .B(G81), .Z(new_n563));
  AOI22_X1  g138(.A1(new_n547), .A2(new_n563), .B1(new_n548), .B2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  AOI22_X1  g146(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(new_n521), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(G91), .B2(new_n547), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n548), .A2(new_n575), .A3(G53), .ZN(new_n576));
  INV_X1    g151(.A(G53), .ZN(new_n577));
  OAI21_X1  g152(.A(KEYINPUT9), .B1(new_n531), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(KEYINPUT81), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n576), .B2(new_n578), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n574), .B1(new_n580), .B2(new_n582), .ZN(G299));
  INV_X1    g158(.A(G168), .ZN(G286));
  OAI221_X1 g159(.A(new_n529), .B1(new_n531), .B2(new_n530), .C1(new_n520), .C2(new_n521), .ZN(G303));
  OAI21_X1  g160(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n527), .A2(G49), .A3(G543), .ZN(new_n587));
  INV_X1    g162(.A(G87), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n539), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n557), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n548), .B2(G48), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n539), .ZN(G305));
  AOI22_X1  g170(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(new_n521), .ZN(new_n597));
  INV_X1    g172(.A(G85), .ZN(new_n598));
  INV_X1    g173(.A(G47), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n539), .A2(new_n598), .B1(new_n531), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n597), .A2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n547), .A2(G92), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n603), .B(KEYINPUT10), .Z(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n557), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n607), .A2(G651), .B1(new_n548), .B2(G54), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n602), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n602), .B1(new_n610), .B2(G868), .ZN(G321));
  NAND2_X1  g187(.A1(G286), .A2(G868), .ZN(new_n613));
  INV_X1    g188(.A(G299), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(G297));
  XNOR2_X1  g190(.A(G297), .B(KEYINPUT82), .ZN(G280));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n610), .B1(G860), .B2(new_n617), .ZN(G148));
  NAND2_X1  g193(.A1(new_n610), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n566), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND3_X1   g197(.A1(new_n485), .A2(new_n467), .A3(new_n469), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(G2100), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n493), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n469), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  AND3_X1   g204(.A1(new_n499), .A2(KEYINPUT84), .A3(G135), .ZN(new_n630));
  AOI21_X1  g205(.A(KEYINPUT84), .B1(new_n499), .B2(G135), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2096), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n626), .A2(new_n633), .A3(new_n634), .ZN(G156));
  XOR2_X1   g210(.A(G2451), .B(G2454), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(KEYINPUT14), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n640), .B(new_n646), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n648), .ZN(G401));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  XNOR2_X1  g228(.A(G2067), .B(G2678), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT86), .ZN(new_n655));
  NOR2_X1   g230(.A1(G2072), .A2(G2078), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n444), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(KEYINPUT17), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  OAI211_X1 g235(.A(new_n653), .B(new_n654), .C1(new_n444), .C2(new_n656), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n655), .A3(new_n653), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2096), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n667), .B(new_n668), .Z(new_n669));
  XNOR2_X1  g244(.A(G1956), .B(G2474), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1961), .B(G1966), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT88), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  INV_X1    g251(.A(new_n669), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n676), .B1(new_n677), .B2(new_n672), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(KEYINPUT89), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(new_n684), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n686), .B1(new_n685), .B2(new_n687), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  NAND2_X1  g265(.A1(G115), .A2(G2104), .ZN(new_n691));
  INV_X1    g266(.A(G127), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n475), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(G2105), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT25), .ZN(new_n696));
  AOI211_X1 g271(.A(new_n694), .B(new_n696), .C1(new_n499), .C2(G139), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(KEYINPUT99), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(KEYINPUT99), .ZN(new_n700));
  OAI21_X1  g275(.A(G29), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G33), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT100), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT100), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n701), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n442), .A3(new_n707), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n702), .A2(G32), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n485), .A2(G105), .A3(new_n469), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT101), .Z(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT26), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n499), .A2(G141), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n493), .A2(G129), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n714), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n709), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT102), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT27), .B(G1996), .ZN(new_n720));
  INV_X1    g295(.A(G160), .ZN(new_n721));
  NAND2_X1  g296(.A1(KEYINPUT24), .A2(G34), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT24), .ZN(new_n723));
  INV_X1    g298(.A(G34), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n721), .A2(G29), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n719), .A2(new_n720), .B1(G2084), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n708), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n442), .B1(new_n705), .B2(new_n707), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT103), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n730), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT103), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n732), .A2(new_n733), .A3(new_n708), .A4(new_n728), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n727), .A2(G2084), .ZN(new_n735));
  NAND2_X1  g310(.A1(G164), .A2(G29), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G27), .B2(G29), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(new_n443), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n443), .ZN(new_n739));
  INV_X1    g314(.A(G28), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n742));
  OR2_X1    g317(.A1(KEYINPUT31), .A2(G11), .ZN(new_n743));
  NAND2_X1  g318(.A1(KEYINPUT31), .A2(G11), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n741), .A2(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n738), .A2(new_n739), .A3(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G16), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n747), .ZN(new_n749));
  AOI211_X1 g324(.A(new_n735), .B(new_n746), .C1(new_n749), .C2(G1961), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n747), .A2(G21), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G168), .B2(new_n747), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n752), .A2(G1966), .B1(new_n632), .B2(new_n702), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G1966), .B2(new_n752), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n750), .B(new_n754), .C1(G1961), .C2(new_n749), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n719), .A2(new_n720), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n731), .A2(new_n734), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT104), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT104), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n731), .A2(new_n734), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n702), .A2(G35), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n501), .B2(G29), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n702), .A2(G26), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT28), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n499), .A2(G140), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n493), .A2(G128), .ZN(new_n773));
  OR2_X1    g348(.A1(G104), .A2(G2105), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n772), .A2(new_n773), .A3(new_n775), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n771), .B1(new_n779), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2067), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT97), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n609), .B2(new_n747), .ZN(new_n784));
  INV_X1    g359(.A(G1348), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n747), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n566), .B2(new_n747), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1341), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2090), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n766), .A2(new_n791), .A3(new_n767), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n769), .A2(new_n781), .A3(new_n790), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n747), .A2(G20), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT23), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n614), .B2(new_n747), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT106), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT105), .B(G1956), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n759), .A2(new_n761), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n747), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n747), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT94), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1971), .ZN(new_n805));
  MUX2_X1   g380(.A(G23), .B(G288), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT33), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1976), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  MUX2_X1   g384(.A(G6), .B(G305), .S(G16), .Z(new_n810));
  OR2_X1    g385(.A1(new_n810), .A2(KEYINPUT93), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n810), .A2(KEYINPUT93), .ZN(new_n812));
  XNOR2_X1  g387(.A(KEYINPUT32), .B(G1981), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  INV_X1    g390(.A(new_n813), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n809), .A2(KEYINPUT34), .A3(new_n814), .A4(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n817), .A2(new_n814), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n805), .A2(new_n808), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n824));
  OAI21_X1  g399(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n825));
  INV_X1    g400(.A(G107), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(G2105), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n827), .B1(new_n493), .B2(G119), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n499), .A2(G131), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT91), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(KEYINPUT91), .B1(new_n499), .B2(G131), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT92), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n835), .B(new_n828), .C1(new_n831), .C2(new_n832), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G29), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n702), .A2(G25), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT90), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT90), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G1991), .Z(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n844), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n747), .A2(G24), .ZN(new_n847));
  INV_X1    g422(.A(G290), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n747), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1986), .ZN(new_n850));
  NOR3_X1   g425(.A1(new_n845), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  AND3_X1   g426(.A1(new_n823), .A2(new_n824), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n824), .B1(new_n823), .B2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT36), .ZN(new_n854));
  OAI22_X1  g429(.A1(new_n852), .A2(new_n853), .B1(KEYINPUT95), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n823), .A2(new_n851), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(KEYINPUT96), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n854), .A2(KEYINPUT95), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n823), .A2(new_n824), .A3(new_n851), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n801), .B1(new_n855), .B2(new_n860), .ZN(G311));
  NAND2_X1  g436(.A1(new_n855), .A2(new_n860), .ZN(new_n862));
  INV_X1    g437(.A(new_n801), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(G150));
  AOI22_X1  g439(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(new_n521), .ZN(new_n866));
  INV_X1    g441(.A(G93), .ZN(new_n867));
  INV_X1    g442(.A(G55), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n539), .A2(new_n867), .B1(new_n531), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G860), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n610), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT107), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT38), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n565), .B(new_n870), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n878), .A2(KEYINPUT39), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n871), .B1(new_n878), .B2(KEYINPUT39), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(G145));
  INV_X1    g456(.A(KEYINPUT40), .ZN(new_n882));
  INV_X1    g457(.A(new_n779), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(G164), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n779), .A2(new_n512), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n499), .A2(G142), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n493), .A2(G130), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n889), .B(G2104), .C1(G118), .C2(new_n469), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n884), .A2(new_n891), .A3(new_n885), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n700), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(KEYINPUT109), .A3(new_n698), .ZN(new_n897));
  INV_X1    g472(.A(new_n717), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n624), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n837), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n834), .A2(KEYINPUT110), .A3(new_n836), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n902), .A2(new_n903), .A3(new_n900), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n897), .B(new_n717), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n908), .A2(new_n904), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n895), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g486(.A1(G162), .A2(new_n632), .ZN(new_n912));
  XNOR2_X1  g487(.A(G160), .B(KEYINPUT108), .ZN(new_n913));
  NAND2_X1  g488(.A1(G162), .A2(new_n632), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n909), .B1(new_n908), .B2(new_n904), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n905), .A2(new_n899), .A3(new_n906), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n918), .A2(new_n919), .A3(new_n893), .A4(new_n894), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n911), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n917), .B1(new_n911), .B2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n882), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n924), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n926), .A2(KEYINPUT40), .A3(new_n922), .A4(new_n921), .ZN(new_n927));
  AND2_X1   g502(.A1(new_n925), .A2(new_n927), .ZN(G395));
  XOR2_X1   g503(.A(G288), .B(KEYINPUT111), .Z(new_n929));
  XNOR2_X1  g504(.A(new_n929), .B(G305), .ZN(new_n930));
  XNOR2_X1  g505(.A(G290), .B(G166), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n930), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n619), .B(new_n877), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n609), .B(G299), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(KEYINPUT41), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n935), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n934), .B2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n933), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(G868), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n944), .B1(G868), .B2(new_n870), .ZN(G295));
  OAI21_X1  g520(.A(new_n944), .B1(G868), .B2(new_n870), .ZN(G331));
  NAND2_X1  g521(.A1(new_n877), .A2(G286), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n566), .A2(new_n870), .ZN(new_n948));
  AND3_X1   g523(.A1(new_n562), .A2(new_n564), .A3(new_n870), .ZN(new_n949));
  OAI21_X1  g524(.A(G168), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n947), .A2(new_n950), .A3(G171), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G171), .B1(new_n947), .B2(new_n950), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n936), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n877), .A2(G286), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n948), .A2(G168), .A3(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(G301), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n938), .A2(new_n957), .A3(new_n940), .A4(new_n951), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n932), .ZN(new_n960));
  INV_X1    g535(.A(new_n932), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n965), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n966), .A3(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(G397));
  NAND2_X1  g546(.A1(new_n470), .A2(new_n479), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n487), .A2(new_n469), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(G40), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n975));
  INV_X1    g550(.A(G1384), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n512), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n512), .A2(new_n976), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(KEYINPUT50), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT122), .B(G2084), .Z(new_n982));
  NAND3_X1  g557(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT45), .B1(new_n512), .B2(new_n976), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT120), .B1(new_n974), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT120), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n987), .A2(new_n988), .A3(G40), .A4(G160), .ZN(new_n989));
  INV_X1    g564(.A(new_n979), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(new_n989), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT121), .ZN(new_n993));
  INV_X1    g568(.A(G1966), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n993), .B1(new_n992), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n983), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(G168), .A2(G8), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1000));
  NAND3_X1  g575(.A1(G303), .A2(G8), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(G303), .B2(G8), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT113), .B1(new_n979), .B2(new_n986), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT113), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n512), .A2(new_n1006), .A3(KEYINPUT45), .A4(new_n976), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n974), .A2(new_n984), .ZN(new_n1009));
  AOI21_X1  g584(.A(G1971), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR4_X1   g585(.A1(new_n980), .A2(new_n974), .A3(G2090), .A4(new_n977), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1004), .B(G8), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n547), .A2(G87), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(G1976), .A3(new_n586), .A4(new_n587), .ZN(new_n1014));
  OAI211_X1 g589(.A(G8), .B(new_n1014), .C1(new_n974), .C2(new_n979), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT52), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n990), .A2(G160), .A3(G40), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1017), .A2(new_n1019), .A3(G8), .A4(new_n1014), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1017), .A2(G8), .ZN(new_n1022));
  XOR2_X1   g597(.A(KEYINPUT115), .B(G1981), .Z(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n593), .B(new_n1024), .C1(new_n594), .C2(new_n539), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n527), .A2(G48), .A3(G543), .ZN(new_n1026));
  XOR2_X1   g601(.A(KEYINPUT116), .B(G86), .Z(new_n1027));
  NAND3_X1  g602(.A1(new_n519), .A2(new_n527), .A3(new_n1027), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1026), .B(new_n1028), .C1(new_n1029), .C2(new_n521), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n1030), .A2(new_n1031), .A3(G1981), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n1030), .B2(G1981), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1025), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1022), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1025), .B(KEYINPUT49), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1021), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT63), .ZN(new_n1039));
  OAI21_X1  g614(.A(G8), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1004), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n999), .A2(new_n1012), .A3(new_n1038), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n997), .A2(new_n998), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT119), .B1(new_n979), .B2(KEYINPUT50), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n512), .A2(new_n1047), .A3(new_n975), .A4(new_n976), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1049), .A2(new_n978), .A3(new_n791), .ZN(new_n1050));
  OAI21_X1  g625(.A(G8), .B1(new_n1050), .B2(new_n1010), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(new_n1041), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(new_n1038), .A3(new_n1012), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1045), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT63), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT123), .B1(new_n1045), .B2(new_n1053), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1044), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1022), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1037), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1021), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1012), .A3(new_n1062), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1049), .A2(new_n978), .ZN(new_n1065));
  OAI22_X1  g640(.A1(new_n1064), .A2(G1971), .B1(new_n1065), .B2(G2090), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1004), .B1(new_n1066), .B2(G8), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n999), .A2(new_n1055), .A3(new_n1068), .ZN(new_n1069));
  AND4_X1   g644(.A1(new_n1044), .A2(new_n1069), .A3(new_n1039), .A4(new_n1057), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1043), .B1(new_n1058), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT127), .ZN(new_n1072));
  OAI211_X1 g647(.A(G168), .B(new_n983), .C1(new_n995), .C2(new_n996), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT51), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1073), .A2(new_n1074), .A3(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n997), .A2(G286), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1076), .A2(G8), .A3(new_n1073), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1077), .B2(KEYINPUT51), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1072), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1064), .A2(new_n443), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n978), .A2(new_n981), .ZN(new_n1084));
  INV_X1    g659(.A(G1961), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1083), .B(new_n1086), .C1(new_n992), .C2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1068), .A2(G171), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1089), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1073), .A2(G8), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1074), .B1(new_n1091), .B2(new_n1076), .ZN(new_n1092));
  OAI211_X1 g667(.A(KEYINPUT127), .B(KEYINPUT62), .C1(new_n1092), .C2(new_n1075), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1080), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1025), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G288), .A2(G1976), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1095), .B1(new_n1061), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(new_n1022), .B(KEYINPUT118), .Z(new_n1098));
  INV_X1    g673(.A(new_n1038), .ZN(new_n1099));
  OAI22_X1  g674(.A1(new_n1097), .A2(new_n1098), .B1(new_n1099), .B2(new_n1012), .ZN(new_n1100));
  XNOR2_X1  g675(.A(G301), .B(KEYINPUT54), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1088), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1103));
  INV_X1    g678(.A(G40), .ZN(new_n1104));
  AOI211_X1 g679(.A(new_n1104), .B(new_n1087), .C1(new_n477), .C2(G2105), .ZN(new_n1105));
  AND4_X1   g680(.A1(new_n973), .A2(new_n1008), .A3(new_n987), .A4(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1102), .B(new_n1068), .C1(new_n1103), .C2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT126), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1084), .A2(new_n785), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1017), .ZN(new_n1111));
  INV_X1    g686(.A(G2067), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT60), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1109), .B1(new_n1114), .B2(new_n609), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1084), .A2(new_n785), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1116));
  OAI211_X1 g691(.A(KEYINPUT126), .B(new_n610), .C1(new_n1116), .C2(KEYINPUT60), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(KEYINPUT60), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n574), .A2(new_n1121), .ZN(new_n1122));
  AOI22_X1  g697(.A1(G299), .A2(KEYINPUT57), .B1(new_n1122), .B2(new_n579), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(KEYINPUT56), .B(G2072), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1064), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(G1956), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1065), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1123), .A2(new_n1126), .A3(KEYINPUT61), .A4(new_n1128), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1124), .A2(new_n1129), .ZN(new_n1132));
  OR2_X1    g707(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1130), .B(new_n1131), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1996), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1064), .A2(new_n1135), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  NAND2_X1  g712(.A1(new_n1017), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n565), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT59), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1139), .B(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1120), .A2(new_n1134), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1130), .B1(new_n609), .B2(new_n1116), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1124), .B2(new_n1129), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1108), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1078), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1100), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1071), .A2(new_n1094), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n974), .A2(new_n987), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1135), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n1151), .A2(new_n717), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n1152), .B(KEYINPUT112), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n779), .B(new_n1112), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1154), .B1(new_n1135), .B2(new_n898), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1153), .B1(new_n1155), .B2(new_n1150), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1150), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n837), .B(new_n843), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OR2_X1    g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G290), .A2(G1986), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1149), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1156), .A2(new_n843), .A3(new_n834), .A4(new_n836), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n883), .A2(new_n1112), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1157), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1160), .A2(new_n1157), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT48), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1159), .A2(new_n1169), .ZN(new_n1170));
  XOR2_X1   g745(.A(new_n1151), .B(KEYINPUT46), .Z(new_n1171));
  NAND2_X1  g746(.A1(new_n1154), .A2(new_n898), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1172), .B2(new_n1150), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1173), .B(KEYINPUT47), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1167), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1164), .A2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g751(.A(G319), .ZN(new_n1178));
  NOR3_X1   g752(.A1(G401), .A2(new_n1178), .A3(G227), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n688), .B2(new_n689), .ZN(new_n1180));
  AOI21_X1  g754(.A(new_n1180), .B1(new_n964), .B2(new_n966), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n926), .A2(new_n922), .A3(new_n921), .ZN(new_n1182));
  AND2_X1   g756(.A1(new_n1181), .A2(new_n1182), .ZN(G308));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(G225));
endmodule


