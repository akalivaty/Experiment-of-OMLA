//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1115,
    new_n1116, new_n1117, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1142, new_n1143, new_n1144, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT64), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND3_X1  g0023(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n209), .B1(new_n220), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XOR2_X1   g0027(.A(G238), .B(G244), .Z(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n244));
  NOR2_X1   g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n216), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT66), .ZN(new_n249));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  AND3_X1   g0050(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT8), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G33), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n248), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n207), .A2(G1), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n260), .B(KEYINPUT68), .ZN(new_n261));
  INV_X1    g0061(.A(new_n244), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n247), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI211_X1 g0064(.A(new_n245), .B(new_n259), .C1(G50), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(KEYINPUT9), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT71), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n265), .A2(KEYINPUT9), .ZN(new_n269));
  INV_X1    g0069(.A(G200), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G222), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G77), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G223), .ZN(new_n276));
  OAI221_X1 g0076(.A(new_n273), .B1(new_n274), .B2(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(G274), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n280), .A2(new_n285), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(G226), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n270), .B1(new_n281), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n281), .A2(new_n289), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NOR3_X1   g0093(.A1(new_n269), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n268), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n291), .A2(G179), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n297), .B(new_n265), .C1(new_n298), .C2(new_n291), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT75), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n288), .A2(G232), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n286), .B2(new_n282), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n271), .A2(G226), .A3(G1698), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n271), .A2(G223), .A3(new_n272), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G87), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n279), .B1(new_n308), .B2(KEYINPUT74), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT74), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n305), .A2(new_n306), .A3(new_n310), .A4(new_n307), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n304), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n312), .A2(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n302), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n312), .A2(new_n313), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n317), .B(KEYINPUT75), .C1(G169), .C2(new_n312), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G68), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n250), .A2(new_n320), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n321), .A2(new_n201), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT7), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n271), .B2(G20), .ZN(new_n327));
  INV_X1    g0127(.A(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT3), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT3), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G33), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n320), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  OR3_X1    g0134(.A1(new_n324), .A2(new_n325), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n325), .B1(new_n324), .B2(new_n334), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n247), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n253), .A2(new_n244), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(new_n264), .B2(new_n253), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n319), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT18), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n316), .A2(new_n318), .B1(new_n337), .B2(new_n339), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n312), .A2(new_n270), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n312), .A2(G190), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n337), .A3(new_n339), .A4(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT17), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n342), .A2(new_n345), .A3(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n255), .A2(G77), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n257), .A2(G50), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n207), .A2(G68), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(KEYINPUT72), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(KEYINPUT72), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n247), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT11), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n244), .A2(KEYINPUT70), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n244), .A2(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(new_n247), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n363), .A2(G68), .A3(new_n261), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n356), .A2(new_n357), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT73), .B(KEYINPUT12), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n361), .B2(G68), .ZN(new_n367));
  INV_X1    g0167(.A(G13), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(G1), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT12), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n353), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n358), .A2(new_n364), .A3(new_n365), .A4(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G97), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n271), .A2(new_n272), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n374), .B1(new_n328), .B2(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n280), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n287), .B1(G238), .B2(new_n288), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT13), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G169), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .B1(new_n313), .B2(new_n382), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n373), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n382), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n373), .B1(new_n387), .B2(G190), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n270), .B2(new_n387), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n288), .A2(G244), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n271), .A2(G232), .A3(new_n272), .ZN(new_n392));
  INV_X1    g0192(.A(G107), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT69), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT69), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G107), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(G238), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n392), .B1(new_n398), .B2(new_n271), .C1(new_n275), .C2(new_n399), .ZN(new_n400));
  AOI211_X1 g0200(.A(new_n287), .B(new_n391), .C1(new_n400), .C2(new_n280), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n401), .A2(new_n313), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n363), .A2(G77), .A3(new_n261), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G20), .A2(G77), .ZN(new_n404));
  INV_X1    g0204(.A(new_n257), .ZN(new_n405));
  XNOR2_X1  g0205(.A(KEYINPUT15), .B(G87), .ZN(new_n406));
  OAI221_X1 g0206(.A(new_n404), .B1(new_n252), .B2(new_n405), .C1(new_n254), .C2(new_n406), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n407), .A2(new_n247), .B1(new_n362), .B2(new_n274), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n403), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n401), .B2(G169), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n402), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(G190), .B2(new_n401), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(new_n270), .B2(new_n401), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n301), .A2(new_n350), .A3(new_n390), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT6), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n417), .A2(new_n375), .A3(G107), .ZN(new_n418));
  XNOR2_X1  g0218(.A(G97), .B(G107), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  OAI22_X1  g0220(.A1(new_n420), .A2(new_n207), .B1(new_n274), .B2(new_n405), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n398), .B1(new_n327), .B2(new_n333), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n247), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n262), .A2(new_n375), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n206), .A2(G33), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n244), .A2(new_n425), .A3(new_n216), .A4(new_n246), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(G97), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n329), .A2(new_n331), .A3(G244), .A4(new_n272), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT4), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n271), .A2(KEYINPUT4), .A3(G244), .A4(new_n272), .ZN(new_n433));
  NAND2_X1  g0233(.A1(G33), .A2(G283), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n280), .ZN(new_n437));
  XNOR2_X1  g0237(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n438));
  OAI211_X1 g0238(.A(G274), .B(new_n279), .C1(new_n438), .C2(G41), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n206), .A2(G45), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT76), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G41), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT76), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n206), .A4(G45), .ZN(new_n447));
  AND3_X1   g0247(.A1(new_n443), .A2(KEYINPUT77), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT77), .B1(new_n443), .B2(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n440), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n443), .A2(new_n447), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n438), .A2(G41), .ZN(new_n452));
  OAI211_X1 g0252(.A(G257), .B(new_n279), .C1(new_n451), .C2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n437), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n429), .B1(G200), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n292), .B2(new_n454), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n254), .A2(KEYINPUT19), .A3(new_n375), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n207), .B1(new_n328), .B2(new_n375), .ZN(new_n458));
  INV_X1    g0258(.A(G87), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n375), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n397), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n457), .B1(new_n461), .B2(KEYINPUT19), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n329), .A2(new_n331), .A3(new_n207), .A4(G68), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT79), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n271), .A2(KEYINPUT79), .A3(new_n207), .A4(G68), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n247), .B1(new_n462), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n362), .A2(new_n406), .ZN(new_n469));
  INV_X1    g0269(.A(new_n406), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT80), .B1(new_n427), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT80), .ZN(new_n472));
  NOR3_X1   g0272(.A1(new_n426), .A2(new_n472), .A3(new_n406), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  AND3_X1   g0274(.A1(new_n468), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n329), .A2(new_n331), .A3(G244), .A4(G1698), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n329), .A2(new_n331), .A3(G238), .A4(new_n272), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n477), .C1(new_n328), .C2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n280), .ZN(new_n480));
  INV_X1    g0280(.A(G250), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(new_n284), .B2(G1), .ZN(new_n482));
  INV_X1    g0282(.A(G274), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n206), .A2(new_n483), .A3(G45), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n279), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n298), .B1(new_n480), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n485), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n313), .B(new_n487), .C1(new_n479), .C2(new_n280), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(G200), .B1(new_n480), .B2(new_n485), .ZN(new_n490));
  AOI211_X1 g0290(.A(G190), .B(new_n487), .C1(new_n479), .C2(new_n280), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n427), .A2(G87), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n468), .A2(new_n469), .A3(new_n493), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n475), .A2(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n454), .A2(new_n298), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n437), .A2(new_n450), .A3(new_n313), .A4(new_n453), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n429), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n456), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n271), .A2(G257), .A3(G1698), .ZN(new_n501));
  INV_X1    g0301(.A(G294), .ZN(new_n502));
  OAI221_X1 g0302(.A(new_n501), .B1(new_n328), .B2(new_n502), .C1(new_n376), .C2(new_n481), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n280), .ZN(new_n504));
  OAI211_X1 g0304(.A(G264), .B(new_n279), .C1(new_n451), .C2(new_n452), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT85), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT85), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n504), .A2(new_n508), .A3(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n450), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n270), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT86), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT86), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n513), .A3(new_n270), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n504), .A2(new_n292), .A3(new_n450), .A4(new_n505), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n512), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n271), .A2(new_n207), .A3(G87), .ZN(new_n517));
  XNOR2_X1  g0317(.A(new_n517), .B(KEYINPUT22), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n393), .A2(G20), .ZN(new_n519));
  OAI22_X1  g0319(.A1(KEYINPUT23), .A2(new_n519), .B1(new_n254), .B2(new_n478), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n398), .A2(G20), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(KEYINPUT23), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n523), .A2(KEYINPUT24), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(KEYINPUT24), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n247), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n369), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(new_n519), .ZN(new_n528));
  XOR2_X1   g0328(.A(KEYINPUT84), .B(KEYINPUT25), .Z(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n530), .B1(G107), .B2(new_n427), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n500), .B1(new_n516), .B2(new_n533), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n507), .A2(G179), .A3(new_n450), .A4(new_n509), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT77), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n451), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n443), .A2(KEYINPUT77), .A3(new_n447), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n439), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(G169), .B1(new_n506), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n535), .A2(new_n540), .B1(new_n526), .B2(new_n531), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G270), .B(new_n279), .C1(new_n451), .C2(new_n452), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT81), .B1(new_n545), .B2(new_n539), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT81), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n450), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n362), .A2(new_n478), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n361), .A2(G116), .A3(new_n248), .A4(new_n425), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n434), .B(new_n207), .C1(G33), .C2(new_n375), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n552), .B(new_n247), .C1(new_n207), .C2(G116), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT20), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n551), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n271), .A2(G257), .A3(new_n272), .ZN(new_n558));
  INV_X1    g0358(.A(G303), .ZN(new_n559));
  INV_X1    g0359(.A(G264), .ZN(new_n560));
  OAI221_X1 g0360(.A(new_n558), .B1(new_n559), .B2(new_n271), .C1(new_n275), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n280), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n313), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n549), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n546), .B2(new_n548), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n557), .A2(KEYINPUT21), .A3(G169), .ZN(new_n567));
  NOR3_X1   g0367(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT82), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n450), .A2(new_n547), .A3(new_n544), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n547), .B1(new_n450), .B2(new_n544), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n562), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n557), .A2(KEYINPUT21), .A3(G169), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n565), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT83), .ZN(new_n576));
  INV_X1    g0376(.A(new_n557), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(new_n298), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT21), .B1(new_n578), .B2(new_n572), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n565), .B(new_n581), .C1(new_n568), .C2(new_n574), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n557), .B1(new_n572), .B2(G200), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n292), .B2(new_n572), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(new_n580), .A3(new_n582), .A4(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n543), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g0386(.A1(new_n416), .A2(new_n586), .ZN(G372));
  NAND2_X1  g0387(.A1(new_n389), .A2(new_n411), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n588), .A2(new_n386), .ZN(new_n589));
  INV_X1    g0389(.A(new_n349), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n342), .B(new_n345), .C1(new_n589), .C2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n299), .B1(new_n591), .B2(new_n296), .ZN(new_n592));
  INV_X1    g0392(.A(new_n416), .ZN(new_n593));
  INV_X1    g0393(.A(new_n475), .ZN(new_n594));
  INV_X1    g0394(.A(new_n489), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT26), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n495), .B2(new_n499), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n495), .A2(new_n499), .A3(new_n597), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OR3_X1    g0401(.A1(new_n575), .A2(KEYINPUT87), .A3(new_n579), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT87), .B1(new_n575), .B2(new_n579), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n542), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n604), .B2(new_n534), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n592), .B1(new_n593), .B2(new_n605), .ZN(G369));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n603), .ZN(new_n607));
  OR3_X1    g0407(.A1(new_n527), .A2(KEYINPUT27), .A3(G20), .ZN(new_n608));
  OAI21_X1  g0408(.A(KEYINPUT27), .B1(new_n527), .B2(G20), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(G213), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(G343), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n577), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n585), .B2(new_n614), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(G330), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n532), .A2(new_n612), .ZN(new_n619));
  XNOR2_X1  g0419(.A(new_n619), .B(KEYINPUT88), .ZN(new_n620));
  AOI211_X1 g0420(.A(new_n541), .B(new_n620), .C1(new_n533), .C2(new_n516), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n542), .A2(new_n613), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n576), .A2(new_n580), .A3(new_n582), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n625), .A2(new_n613), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n621), .A2(new_n626), .B1(new_n541), .B2(new_n613), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(G399));
  INV_X1    g0428(.A(new_n210), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n629), .A2(G41), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n397), .A2(G116), .A3(new_n460), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G1), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n214), .B2(new_n631), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT28), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n541), .A2(new_n579), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n576), .A2(new_n582), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT91), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n534), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT89), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n600), .B1(new_n640), .B2(new_n598), .ZN(new_n641));
  NOR4_X1   g0441(.A1(new_n495), .A2(new_n499), .A3(KEYINPUT89), .A4(new_n597), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n596), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(KEYINPUT90), .B(new_n596), .C1(new_n641), .C2(new_n642), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n639), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n638), .B1(new_n637), .B2(new_n534), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n613), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT29), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n605), .A2(KEYINPUT29), .A3(new_n612), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n586), .A2(new_n613), .ZN(new_n654));
  INV_X1    g0454(.A(new_n454), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n487), .B1(new_n479), .B2(new_n280), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n564), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n507), .A2(new_n509), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(new_n658), .A3(new_n549), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT30), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n655), .A2(G179), .A3(new_n656), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n510), .A3(new_n572), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n612), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT31), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n654), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n668), .A2(G330), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n653), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n635), .B1(new_n670), .B2(G1), .ZN(G364));
  NOR2_X1   g0471(.A1(new_n368), .A2(G20), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n206), .B1(new_n672), .B2(G45), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n630), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n618), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(G330), .B2(new_n616), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n216), .B1(G20), .B2(new_n298), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n292), .A2(G179), .A3(G200), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n207), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n207), .A2(new_n313), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G200), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n684), .A2(new_n292), .ZN(new_n685));
  AOI22_X1  g0485(.A1(G294), .A2(new_n682), .B1(new_n685), .B2(G326), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT95), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(G190), .A3(new_n270), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n207), .A2(G179), .ZN(new_n690));
  NOR2_X1   g0490(.A1(G190), .A2(G200), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n689), .A2(G322), .B1(new_n693), .B2(G329), .ZN(new_n694));
  INV_X1    g0494(.A(G311), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n683), .A2(new_n691), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n694), .B(new_n332), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n684), .A2(G190), .ZN(new_n698));
  INV_X1    g0498(.A(G317), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT33), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n699), .A2(KEYINPUT33), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G283), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n690), .A2(new_n292), .A3(G200), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n690), .A2(G190), .A3(G200), .ZN(new_n705));
  OAI221_X1 g0505(.A(new_n702), .B1(new_n703), .B2(new_n704), .C1(new_n559), .C2(new_n705), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n687), .A2(new_n697), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n704), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G107), .ZN(new_n709));
  INV_X1    g0509(.A(G159), .ZN(new_n710));
  OAI21_X1  g0510(.A(KEYINPUT32), .B1(new_n692), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n705), .ZN(new_n713));
  AOI211_X1 g0513(.A(new_n332), .B(new_n712), .C1(G87), .C2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n685), .ZN(new_n715));
  INV_X1    g0515(.A(new_n698), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n202), .A2(new_n715), .B1(new_n716), .B2(new_n320), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n692), .A2(KEYINPUT32), .A3(new_n710), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n681), .A2(new_n375), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  OAI22_X1  g0520(.A1(new_n688), .A2(new_n250), .B1(new_n696), .B2(new_n274), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT94), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n679), .B1(new_n707), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n726), .A2(KEYINPUT93), .A3(G20), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT93), .B1(new_n726), .B2(G20), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n678), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n629), .A2(new_n332), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n732), .A2(G355), .B1(new_n478), .B2(new_n629), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n239), .A2(new_n284), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n210), .A2(new_n332), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n736), .B1(new_n284), .B2(new_n215), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n733), .A2(KEYINPUT92), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n731), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n675), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n724), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n729), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n742), .B1(new_n616), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n677), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(G396));
  NOR2_X1   g0546(.A1(new_n412), .A2(new_n612), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n409), .A2(new_n612), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n414), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n412), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  OR3_X1    g0552(.A1(new_n605), .A2(new_n612), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n752), .B1(new_n605), .B2(new_n612), .ZN(new_n756));
  XOR2_X1   g0556(.A(new_n755), .B(new_n756), .Z(new_n757));
  OR2_X1    g0557(.A1(new_n757), .A2(new_n669), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n669), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n758), .A2(new_n741), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n678), .A2(new_n725), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n741), .B1(new_n274), .B2(new_n761), .ZN(new_n762));
  AOI22_X1  g0562(.A1(new_n698), .A2(G283), .B1(new_n685), .B2(G303), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n393), .B2(new_n705), .ZN(new_n764));
  AOI22_X1  g0564(.A1(new_n689), .A2(G294), .B1(new_n693), .B2(G311), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n765), .B(new_n332), .C1(new_n478), .C2(new_n696), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n704), .A2(new_n459), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n764), .A2(new_n766), .A3(new_n719), .A4(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n696), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n689), .A2(G143), .B1(new_n769), .B2(G159), .ZN(new_n770));
  INV_X1    g0570(.A(G137), .ZN(new_n771));
  INV_X1    g0571(.A(G150), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n770), .B1(new_n715), .B2(new_n771), .C1(new_n772), .C2(new_n716), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT34), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n202), .A2(new_n705), .B1(new_n704), .B2(new_n320), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n777));
  INV_X1    g0577(.A(G132), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n271), .B1(new_n692), .B2(new_n778), .C1(new_n681), .C2(new_n250), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n768), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n752), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n762), .B1(new_n679), .B2(new_n781), .C1(new_n782), .C2(new_n726), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n760), .A2(new_n783), .ZN(G384));
  INV_X1    g0584(.A(new_n420), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT35), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT35), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n786), .A2(G116), .A3(new_n217), .A4(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT36), .Z(new_n789));
  OR3_X1    g0589(.A1(new_n214), .A2(new_n274), .A3(new_n321), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n202), .A2(G68), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n206), .B(G13), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n610), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n340), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n348), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT37), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n341), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(KEYINPUT37), .B1(new_n343), .B2(new_n796), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n350), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n802), .B2(new_n795), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT38), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n795), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n350), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(KEYINPUT38), .A3(new_n801), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n805), .A2(KEYINPUT39), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT99), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n798), .B1(new_n797), .B2(new_n341), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n350), .A2(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n799), .A2(KEYINPUT99), .A3(new_n800), .ZN(new_n813));
  AOI21_X1  g0613(.A(KEYINPUT38), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n807), .A2(KEYINPUT38), .A3(new_n801), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n809), .B1(new_n816), .B2(KEYINPUT39), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n386), .A2(new_n612), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n373), .A2(new_n612), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT98), .Z(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n390), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n386), .A2(new_n389), .A3(new_n821), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n753), .B2(new_n748), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n805), .A2(new_n808), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n345), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n343), .A2(new_n344), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n610), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n819), .A2(new_n829), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n592), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n653), .B2(new_n416), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n833), .B(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT40), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n805), .A2(new_n837), .A3(new_n808), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n752), .B1(new_n654), .B2(new_n667), .ZN(new_n839));
  NAND2_X1  g0639(.A1(KEYINPUT100), .A2(KEYINPUT40), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n838), .A2(new_n839), .A3(new_n825), .A4(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT31), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n666), .B(new_n842), .ZN(new_n843));
  NOR3_X1   g0643(.A1(new_n543), .A2(new_n585), .A3(new_n612), .ZN(new_n844));
  OAI211_X1 g0644(.A(new_n825), .B(new_n782), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n816), .B1(KEYINPUT100), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n841), .B1(new_n846), .B2(new_n837), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n416), .A2(new_n668), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n848), .ZN(new_n850));
  AND3_X1   g0650(.A1(new_n849), .A2(G330), .A3(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n836), .A2(new_n851), .B1(new_n206), .B2(new_n672), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n836), .A2(new_n851), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n793), .B1(new_n852), .B2(new_n853), .ZN(G367));
  AND2_X1   g0654(.A1(new_n621), .A2(new_n626), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n429), .A2(new_n612), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n456), .A2(new_n499), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n499), .B2(new_n613), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n499), .B1(new_n542), .B2(new_n857), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n859), .A2(KEYINPUT42), .B1(new_n613), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(KEYINPUT42), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n494), .A2(new_n612), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n496), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n864), .B1(new_n596), .B2(new_n863), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT43), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(KEYINPUT43), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n624), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT101), .B1(new_n870), .B2(new_n858), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AND3_X1   g0672(.A1(new_n870), .A2(KEYINPUT101), .A3(new_n858), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n630), .B(KEYINPUT41), .Z(new_n875));
  NAND2_X1  g0675(.A1(new_n627), .A2(new_n858), .ZN(new_n876));
  XOR2_X1   g0676(.A(new_n876), .B(KEYINPUT45), .Z(new_n877));
  NOR2_X1   g0677(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n627), .A2(new_n858), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n878), .B1(new_n627), .B2(new_n858), .ZN(new_n880));
  NAND2_X1  g0680(.A1(KEYINPUT102), .A2(KEYINPUT44), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n877), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n870), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT103), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n883), .A2(KEYINPUT103), .A3(new_n870), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n623), .A2(new_n626), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n855), .ZN(new_n889));
  XNOR2_X1  g0689(.A(new_n889), .B(new_n617), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n670), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n877), .B(new_n624), .C1(new_n879), .C2(new_n882), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n886), .A2(new_n887), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n875), .B1(new_n894), .B2(new_n670), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n872), .B(new_n874), .C1(new_n895), .C2(new_n674), .ZN(new_n896));
  INV_X1    g0696(.A(new_n235), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n730), .B1(new_n210), .B2(new_n406), .C1(new_n897), .C2(new_n736), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT104), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n741), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n271), .B1(new_n692), .B2(new_n771), .C1(new_n688), .C2(new_n772), .ZN(new_n902));
  INV_X1    g0702(.A(G143), .ZN(new_n903));
  OAI22_X1  g0703(.A1(new_n715), .A2(new_n903), .B1(new_n705), .B2(new_n250), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n681), .A2(new_n320), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n704), .A2(new_n274), .ZN(new_n906));
  OR4_X1    g0706(.A1(new_n902), .A2(new_n904), .A3(new_n905), .A4(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n698), .A2(G159), .B1(new_n769), .B2(G50), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT105), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n698), .A2(G294), .B1(new_n708), .B2(G97), .ZN(new_n910));
  OAI221_X1 g0710(.A(new_n910), .B1(new_n695), .B2(new_n715), .C1(new_n398), .C2(new_n681), .ZN(new_n911));
  AOI22_X1  g0711(.A1(G283), .A2(new_n769), .B1(new_n693), .B2(G317), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n271), .B1(new_n689), .B2(G303), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n713), .A2(KEYINPUT46), .A3(G116), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT46), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n705), .B2(new_n478), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n912), .A2(new_n913), .A3(new_n914), .A4(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n907), .A2(new_n909), .B1(new_n911), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT47), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n901), .B1(new_n919), .B2(new_n678), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n865), .B2(new_n743), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n896), .A2(new_n921), .ZN(G387));
  NAND2_X1  g0722(.A1(new_n890), .A2(new_n674), .ZN(new_n923));
  XOR2_X1   g0723(.A(new_n923), .B(KEYINPUT106), .Z(new_n924));
  NOR2_X1   g0724(.A1(new_n623), .A2(new_n743), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n689), .A2(G317), .B1(new_n769), .B2(G303), .ZN(new_n926));
  INV_X1    g0726(.A(G322), .ZN(new_n927));
  OAI221_X1 g0727(.A(new_n926), .B1(new_n715), .B2(new_n927), .C1(new_n695), .C2(new_n716), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT48), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n682), .A2(G283), .B1(new_n713), .B2(G294), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n934), .A2(KEYINPUT49), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n271), .B1(new_n693), .B2(G326), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n478), .B2(new_n704), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(KEYINPUT49), .B2(new_n934), .ZN(new_n939));
  XNOR2_X1  g0739(.A(KEYINPUT107), .B(G150), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n696), .A2(new_n320), .B1(new_n692), .B2(new_n940), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n332), .B(new_n941), .C1(G50), .C2(new_n689), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n681), .A2(new_n406), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G97), .B2(new_n708), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n685), .A2(G159), .B1(new_n713), .B2(G77), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n253), .A2(new_n698), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n942), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n679), .B1(new_n939), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n232), .A2(G45), .ZN(new_n949));
  INV_X1    g0749(.A(new_n732), .ZN(new_n950));
  OAI22_X1  g0750(.A1(new_n949), .A2(new_n736), .B1(new_n632), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n252), .A2(G50), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT50), .ZN(new_n953));
  AOI21_X1  g0753(.A(G45), .B1(G68), .B2(G77), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n632), .A3(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n951), .A2(new_n955), .B1(new_n393), .B2(new_n629), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n675), .B1(new_n956), .B2(new_n731), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n925), .A2(new_n948), .A3(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n924), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n892), .A2(new_n631), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n670), .B2(new_n890), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n961), .ZN(G393));
  NAND2_X1  g0762(.A1(new_n884), .A2(new_n893), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n631), .B1(new_n963), .B2(new_n891), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n894), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT112), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n884), .A2(new_n674), .A3(new_n893), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n730), .B1(new_n375), .B2(new_n210), .C1(new_n242), .C2(new_n736), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n741), .B1(new_n968), .B2(KEYINPUT108), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(KEYINPUT108), .B2(new_n968), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n681), .A2(new_n274), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n271), .B1(new_n696), .B2(new_n252), .C1(new_n459), .C2(new_n704), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(G50), .C2(new_n698), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n715), .A2(new_n772), .B1(new_n710), .B2(new_n688), .ZN(new_n974));
  XOR2_X1   g0774(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n975));
  OR2_X1    g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n705), .A2(new_n320), .B1(new_n692), .B2(new_n903), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n974), .A2(new_n975), .B1(new_n977), .B2(KEYINPUT110), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n973), .A2(new_n976), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n709), .B(new_n332), .C1(new_n927), .C2(new_n692), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G283), .B2(new_n713), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT111), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n715), .A2(new_n699), .B1(new_n695), .B2(new_n688), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT52), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n681), .A2(new_n478), .B1(new_n696), .B2(new_n502), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G303), .B2(new_n698), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n980), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n970), .B1(new_n989), .B2(new_n678), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n858), .B2(new_n743), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n967), .A2(new_n991), .ZN(new_n992));
  AND3_X1   g0792(.A1(new_n965), .A2(new_n966), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n966), .B1(new_n965), .B2(new_n992), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(G390));
  INV_X1    g0796(.A(new_n818), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n817), .B1(new_n827), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT113), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n613), .B(new_n751), .C1(new_n647), .C2(new_n648), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n748), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n825), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n818), .B1(new_n814), .B2(new_n815), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n999), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n826), .B1(new_n1000), .B2(new_n748), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1006), .A2(KEYINPUT113), .A3(new_n1003), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n998), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n839), .A2(G330), .A3(new_n825), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n669), .A2(new_n416), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n592), .B(new_n1012), .C1(new_n652), .C2(new_n593), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n668), .A2(G330), .A3(new_n782), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n826), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n1009), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n753), .A2(new_n748), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n748), .A3(new_n1009), .A4(new_n1000), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1013), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n998), .B(new_n1009), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1011), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1011), .A2(new_n1021), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1020), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1023), .A2(KEYINPUT114), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT114), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n630), .B(new_n1022), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT115), .B1(new_n1023), .B2(new_n673), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT115), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1011), .A2(new_n1029), .A3(new_n674), .A4(new_n1021), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n817), .A2(new_n725), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n761), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n675), .B1(new_n253), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n716), .A2(new_n771), .B1(new_n704), .B2(new_n202), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n685), .A2(G128), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n710), .B2(new_n681), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(KEYINPUT54), .B(G143), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n688), .A2(new_n778), .B1(new_n696), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(G125), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n271), .B1(new_n692), .B2(new_n1039), .ZN(new_n1040));
  NOR4_X1   g0840(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n705), .A2(new_n940), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT53), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n715), .A2(new_n703), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n971), .B(new_n1044), .C1(new_n397), .C2(new_n698), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n320), .A2(new_n704), .B1(new_n705), .B2(new_n459), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n332), .B1(new_n688), .B2(new_n478), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n696), .A2(new_n375), .B1(new_n692), .B2(new_n502), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1046), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1041), .A2(new_n1043), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1033), .B1(new_n1051), .B2(new_n678), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1028), .A2(new_n1030), .B1(new_n1031), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1027), .A2(new_n1053), .ZN(G378));
  INV_X1    g0854(.A(new_n1013), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1022), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(KEYINPUT119), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT119), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1022), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n265), .A2(new_n610), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT55), .Z(new_n1062));
  XNOR2_X1  g0862(.A(new_n301), .B(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1063), .B(new_n1065), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n847), .A2(new_n1066), .A3(G330), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n847), .B2(G330), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n833), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n847), .A2(G330), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n1066), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n819), .A2(new_n829), .A3(new_n832), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n847), .A2(new_n1066), .A3(G330), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1069), .A2(new_n1075), .A3(KEYINPUT118), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT118), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1077), .B(new_n833), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(KEYINPUT57), .B1(new_n1060), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT57), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1069), .B2(new_n1075), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1022), .A2(new_n1058), .A3(new_n1055), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1058), .B1(new_n1022), .B2(new_n1055), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n630), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1080), .A2(new_n1086), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1039), .A2(new_n715), .B1(new_n716), .B2(new_n778), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n689), .A2(G128), .B1(new_n769), .B2(G137), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n705), .B2(new_n1037), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1088), .B(new_n1090), .C1(G150), .C2(new_n682), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OR2_X1    g0892(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(KEYINPUT59), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n708), .A2(G159), .ZN(new_n1095));
  AOI211_X1 g0895(.A(G33), .B(G41), .C1(new_n693), .C2(G124), .ZN(new_n1096));
  AND4_X1   g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n271), .A2(G41), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n703), .B2(new_n692), .C1(new_n406), .C2(new_n696), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n905), .B(new_n1099), .C1(G77), .C2(new_n713), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n716), .A2(new_n375), .B1(new_n704), .B2(new_n250), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G116), .B2(new_n685), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n688), .A2(new_n393), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT116), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT58), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g0907(.A(G50), .B(new_n1098), .C1(new_n328), .C2(new_n283), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1109));
  NOR4_X1   g0909(.A1(new_n1097), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n675), .B1(G50), .B2(new_n1032), .C1(new_n1110), .C2(new_n679), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1071), .B2(new_n725), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n1079), .B2(new_n674), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1087), .A2(new_n1113), .ZN(G375));
  NAND2_X1  g0914(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n674), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n698), .A2(G116), .B1(new_n685), .B2(G294), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n375), .B2(new_n705), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n271), .B1(new_n693), .B2(G303), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n703), .B2(new_n688), .C1(new_n398), .C2(new_n696), .ZN(new_n1120));
  NOR4_X1   g0920(.A1(new_n1118), .A2(new_n1120), .A3(new_n906), .A4(new_n943), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n332), .B1(new_n693), .B2(G128), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n771), .B2(new_n688), .C1(new_n772), .C2(new_n696), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n682), .A2(G50), .B1(new_n713), .B2(G159), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n778), .B2(new_n715), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n716), .A2(new_n1037), .B1(new_n704), .B2(new_n250), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1123), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n678), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n741), .B1(new_n320), .B2(new_n761), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n825), .C2(new_n726), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1116), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n875), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1024), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1115), .A2(new_n1055), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(G381));
  INV_X1    g0935(.A(G384), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n959), .A2(new_n745), .A3(new_n1136), .A4(new_n961), .ZN(new_n1137));
  NOR4_X1   g0937(.A1(G390), .A2(G387), .A3(G381), .A4(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(G378), .ZN(new_n1139));
  INV_X1    g0939(.A(G375), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(G407));
  NAND2_X1  g0941(.A1(new_n611), .A2(G213), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT120), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1139), .A3(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(G407), .A2(G213), .A3(new_n1144), .ZN(G409));
  OR2_X1    g0945(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n1024), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(KEYINPUT122), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT122), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1146), .A2(new_n1149), .A3(new_n1024), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1134), .A2(KEYINPUT60), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n630), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G384), .B(new_n1131), .C1(new_n1151), .C2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1153), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1131), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1136), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1143), .A2(G2897), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT124), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1142), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1154), .A2(G2897), .A3(new_n1157), .A4(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1161), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(G378), .B(new_n1113), .C1(new_n1080), .C2(new_n1086), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1079), .B(new_n1132), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1112), .B1(new_n1169), .B2(new_n674), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(new_n1139), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1167), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT121), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT121), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1167), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1174), .A2(new_n1142), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(G387), .A2(new_n995), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n896), .B(new_n921), .C1(new_n993), .C2(new_n994), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(G393), .B(new_n745), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT61), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1179), .A2(new_n1182), .A3(new_n1180), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1143), .B1(new_n1167), .B2(new_n1172), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1158), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1189), .A2(KEYINPUT63), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1187), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1174), .A2(new_n1142), .A3(new_n1189), .A4(new_n1176), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1194));
  OAI211_X1 g0994(.A(new_n1178), .B(new_n1191), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1160), .A2(new_n1163), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1185), .B1(new_n1196), .B2(new_n1188), .ZN(new_n1197));
  AND3_X1   g0997(.A1(new_n1188), .A2(new_n1189), .A3(KEYINPUT62), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT62), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1192), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT125), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1198), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1192), .A2(KEYINPUT125), .A3(new_n1199), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1184), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1186), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1195), .B1(new_n1204), .B2(new_n1207), .ZN(G405));
  NAND2_X1  g1008(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1158), .A2(KEYINPUT126), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1209), .B(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1167), .B1(new_n1158), .B2(KEYINPUT126), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1139), .B2(G375), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1212), .B(new_n1214), .ZN(G402));
endmodule


