//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT1), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n188), .A2(new_n190), .A3(new_n191), .A4(G128), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n189), .A2(G146), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n187), .B2(G143), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n189), .A2(KEYINPUT65), .A3(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(new_n188), .B2(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n192), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT66), .A2(G134), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT66), .A2(G134), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n201), .A2(new_n202), .A3(G137), .ZN(new_n203));
  INV_X1    g017(.A(G137), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT67), .B1(new_n204), .B2(G134), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G137), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n203), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(KEYINPUT11), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n201), .B2(new_n202), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n204), .A2(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n200), .A2(new_n210), .A3(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n195), .A2(new_n196), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n188), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT0), .A2(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(KEYINPUT0), .A2(G128), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n188), .A2(new_n190), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n222), .A2(new_n226), .B1(new_n227), .B2(new_n223), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT66), .B(G134), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n214), .B1(new_n229), .B2(new_n211), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n213), .B1(new_n230), .B2(new_n216), .ZN(new_n231));
  INV_X1    g045(.A(new_n217), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n234), .B(new_n235), .Z(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n200), .A2(new_n210), .A3(KEYINPUT68), .A4(new_n217), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n220), .A2(new_n233), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT30), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n220), .A2(new_n238), .A3(new_n233), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n200), .A2(new_n210), .A3(new_n217), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n188), .A2(new_n190), .A3(new_n223), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n197), .B2(new_n225), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n247), .B2(new_n217), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT64), .B1(new_n243), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n241), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  AOI211_X1 g064(.A(KEYINPUT64), .B(KEYINPUT30), .C1(new_n233), .C2(new_n218), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n240), .B1(new_n252), .B2(new_n236), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n255));
  INV_X1    g069(.A(G237), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n255), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT26), .B(G101), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n254), .A2(KEYINPUT71), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT29), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n264));
  INV_X1    g078(.A(new_n261), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n253), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n233), .A2(new_n237), .A3(new_n218), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n233), .A2(new_n218), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n236), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n269), .B(new_n271), .C1(new_n268), .C2(new_n239), .ZN(new_n272));
  OR2_X1    g086(.A1(new_n272), .A2(new_n261), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n262), .A2(new_n263), .A3(new_n266), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n269), .A2(KEYINPUT72), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n242), .A2(new_n236), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n276), .A2(new_n239), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n277), .B2(new_n268), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n239), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(KEYINPUT72), .A3(KEYINPUT28), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n278), .A2(KEYINPUT29), .A3(new_n265), .A4(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(KEYINPUT73), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n274), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G472), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n250), .A2(new_n237), .A3(new_n251), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n240), .A2(new_n261), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n251), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n247), .A2(new_n217), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n219), .A2(new_n218), .B1(new_n298), .B2(new_n228), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n238), .A2(new_n299), .B1(new_n270), .B2(KEYINPUT64), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(new_n236), .C1(new_n300), .C2(new_n241), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT31), .A3(new_n294), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n272), .A2(new_n261), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n291), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n304), .ZN(new_n306));
  AOI211_X1 g120(.A(KEYINPUT70), .B(new_n306), .C1(new_n296), .C2(new_n302), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n290), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT32), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT74), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT32), .B(new_n290), .C1(new_n305), .C2(new_n307), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n290), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n293), .A2(new_n295), .A3(new_n292), .ZN(new_n315));
  AOI21_X1  g129(.A(KEYINPUT31), .B1(new_n301), .B2(new_n294), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n304), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n303), .A2(new_n291), .A3(new_n304), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n314), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n289), .B1(new_n313), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT76), .B1(new_n323), .B2(G128), .ZN(new_n324));
  OR2_X1    g138(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(KEYINPUT23), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n325), .B(new_n326), .C1(G119), .C2(new_n198), .ZN(new_n327));
  XNOR2_X1  g141(.A(G119), .B(G128), .ZN(new_n328));
  XOR2_X1   g142(.A(KEYINPUT24), .B(G110), .Z(new_n329));
  OAI22_X1  g143(.A1(new_n327), .A2(G110), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(G125), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT77), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n331), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n338), .A2(KEYINPUT16), .ZN(new_n341));
  OAI21_X1  g155(.A(G146), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n330), .B(new_n342), .C1(G146), .C2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n341), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n335), .A2(new_n337), .A3(G140), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(KEYINPUT77), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n347), .B1(new_n333), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n187), .B(new_n346), .C1(new_n349), .C2(new_n331), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n327), .A2(G110), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n329), .A2(new_n328), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT75), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n354), .B1(new_n353), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n345), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G137), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n345), .B(new_n362), .C1(new_n357), .C2(new_n358), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G217), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(G234), .B2(new_n282), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(G902), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT79), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n364), .A2(new_n282), .A3(new_n365), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT25), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n364), .A2(new_n374), .A3(new_n282), .A4(new_n365), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n373), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n366), .A2(new_n377), .A3(new_n369), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n198), .A2(G143), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT92), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n380), .B(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n189), .A2(G128), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT13), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n189), .A2(KEYINPUT13), .A3(G128), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT93), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n380), .A2(new_n381), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT92), .B1(new_n198), .B2(G143), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n383), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n229), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g208(.A(G116), .B(G122), .ZN(new_n395));
  INV_X1    g209(.A(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OR2_X1    g211(.A1(new_n395), .A2(new_n396), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT93), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n387), .A2(new_n400), .A3(G134), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n389), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT94), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n392), .B(new_n393), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT14), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n395), .A2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G122), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G116), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n396), .B1(new_n408), .B2(KEYINPUT14), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n406), .A2(new_n409), .B1(new_n396), .B2(new_n395), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n403), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n229), .B1(new_n382), .B2(new_n383), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n403), .B(new_n410), .C1(new_n412), .C2(new_n394), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n402), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT9), .B(G234), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n417), .A2(new_n367), .A3(G953), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n402), .B(new_n418), .C1(new_n411), .C2(new_n414), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n282), .ZN(new_n423));
  INV_X1    g237(.A(G478), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT95), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(KEYINPUT15), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n424), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n423), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n256), .A2(new_n257), .A3(G214), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(new_n189), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT17), .A3(G131), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n342), .A2(new_n350), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT90), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(new_n431), .B(G143), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n437), .B(G131), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n342), .A2(new_n350), .A3(KEYINPUT90), .A4(new_n433), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n436), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n344), .A2(G146), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n336), .A2(new_n339), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(G146), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n446), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT18), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n432), .B1(new_n450), .B2(new_n213), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n437), .A2(KEYINPUT18), .A3(G131), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(G104), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n442), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n457), .B1(new_n442), .B2(new_n454), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n282), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G475), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n430), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n457), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n344), .A2(KEYINPUT19), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n466), .B1(new_n444), .B2(KEYINPUT19), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n467), .A2(new_n187), .ZN(new_n468));
  INV_X1    g282(.A(new_n342), .ZN(new_n469));
  NOR3_X1   g283(.A1(new_n468), .A2(new_n438), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g284(.A1(new_n447), .A2(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n458), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(G475), .A2(G902), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  XOR2_X1   g289(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(KEYINPUT91), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT91), .ZN(new_n478));
  INV_X1    g292(.A(new_n474), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n458), .B2(new_n472), .ZN(new_n480));
  INV_X1    g294(.A(new_n476), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n464), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G952), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n487), .A2(KEYINPUT96), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(KEYINPUT96), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n257), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(G234), .B2(G237), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n491), .B(KEYINPUT97), .Z(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G898), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT98), .ZN(new_n494));
  AOI211_X1 g308(.A(new_n282), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n486), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT87), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n200), .A2(new_n337), .ZN(new_n500));
  OAI211_X1 g314(.A(G125), .B(new_n244), .C1(new_n197), .C2(new_n225), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(G224), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(G953), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n502), .B(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT80), .ZN(new_n507));
  XNOR2_X1  g321(.A(G104), .B(G107), .ZN(new_n508));
  INV_X1    g322(.A(G101), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n396), .A2(G104), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n456), .A2(G107), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(KEYINPUT80), .A3(G101), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT3), .B1(new_n456), .B2(G107), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n396), .A3(G104), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n515), .A2(new_n517), .A3(new_n509), .A4(new_n512), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n510), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT5), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n323), .A3(G116), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT82), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(G113), .A3(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n235), .ZN(new_n525));
  OR2_X1    g339(.A1(new_n525), .A2(new_n234), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n519), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n515), .A2(new_n517), .A3(new_n512), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(G101), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT4), .A3(new_n518), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT4), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n531), .A3(G101), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n236), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT83), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(G110), .B(G122), .Z(new_n537));
  NAND3_X1  g351(.A1(new_n527), .A2(new_n533), .A3(KEYINPUT83), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT6), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(KEYINPUT6), .A3(new_n537), .A4(new_n538), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n534), .A2(new_n537), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n506), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n505), .A2(KEYINPUT84), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n500), .A2(new_n546), .A3(new_n501), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n505), .A2(KEYINPUT7), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n524), .A2(new_n526), .ZN(new_n550));
  INV_X1    g364(.A(new_n519), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n527), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n537), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT85), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT85), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n549), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n559), .A3(new_n543), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n545), .A2(new_n560), .A3(new_n282), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT86), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n499), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n563), .ZN(new_n566));
  INV_X1    g380(.A(new_n563), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n545), .A2(new_n560), .A3(new_n282), .A4(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n565), .B1(new_n569), .B2(KEYINPUT87), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n192), .B1(new_n227), .B2(new_n199), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n571), .A2(new_n518), .A3(new_n514), .A4(new_n510), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n519), .B2(new_n200), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n298), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT12), .ZN(new_n575));
  XNOR2_X1  g389(.A(G110), .B(G140), .ZN(new_n576));
  INV_X1    g390(.A(G227), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(G953), .ZN(new_n578));
  XOR2_X1   g392(.A(new_n576), .B(new_n578), .Z(new_n579));
  INV_X1    g393(.A(KEYINPUT10), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n519), .A2(KEYINPUT10), .A3(new_n200), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n228), .A2(new_n530), .A3(new_n532), .ZN(new_n583));
  INV_X1    g397(.A(new_n298), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n581), .A2(new_n582), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n573), .A2(new_n586), .A3(new_n298), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n575), .A2(new_n579), .A3(new_n585), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n298), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n590), .A2(new_n585), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT81), .B(new_n588), .C1(new_n591), .C2(new_n579), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n588), .A2(KEYINPUT81), .ZN(new_n593));
  INV_X1    g407(.A(G469), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n592), .A2(new_n593), .A3(new_n594), .A4(new_n282), .ZN(new_n595));
  NAND2_X1  g409(.A1(G469), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n579), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n591), .A2(new_n597), .ZN(new_n598));
  AND4_X1   g412(.A1(new_n597), .A2(new_n575), .A3(new_n585), .A4(new_n587), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n595), .B(new_n596), .C1(new_n594), .C2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G214), .B1(G237), .B2(G902), .ZN(new_n602));
  INV_X1    g416(.A(G221), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n416), .B2(new_n282), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n602), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n498), .A2(new_n570), .A3(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n322), .A2(new_n379), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n509), .ZN(G3));
  OAI21_X1  g424(.A(new_n282), .B1(new_n305), .B2(new_n307), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n320), .B1(G472), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n379), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n601), .A2(new_n605), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n602), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n566), .B2(new_n568), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n420), .A2(KEYINPUT33), .A3(new_n421), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT33), .B1(new_n420), .B2(new_n421), .ZN(new_n620));
  OAI21_X1  g434(.A(G478), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n422), .A2(new_n424), .A3(new_n282), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n424), .A2(new_n282), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n485), .B2(new_n462), .ZN(new_n626));
  INV_X1    g440(.A(new_n497), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n618), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n616), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT99), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n477), .A2(new_n633), .A3(new_n482), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n480), .A2(new_n481), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n633), .B1(new_n477), .B2(new_n482), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT101), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n477), .A2(new_n482), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(KEYINPUT100), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n635), .A4(new_n634), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n430), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n463), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n627), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n643), .A2(KEYINPUT102), .A3(new_n627), .A4(new_n645), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n569), .A2(new_n606), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n650), .A2(new_n613), .A3(new_n612), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT35), .B(G107), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G9));
  NOR2_X1   g468(.A1(new_n363), .A2(KEYINPUT36), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n359), .B(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n369), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n376), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n612), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n660), .A2(new_n608), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT103), .B(KEYINPUT37), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G110), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n313), .A2(new_n321), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n288), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n659), .ZN(new_n667));
  INV_X1    g481(.A(new_n651), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n495), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n492), .A2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n643), .A2(new_n645), .A3(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n667), .A2(new_n668), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n198), .ZN(G30));
  NAND2_X1  g489(.A1(new_n566), .A2(new_n568), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n564), .B1(new_n676), .B2(new_n499), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT38), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n485), .A2(new_n462), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n644), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n671), .B(KEYINPUT39), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n615), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n683), .B1(new_n686), .B2(KEYINPUT40), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n680), .A2(new_n659), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n253), .A2(new_n261), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n282), .B1(new_n279), .B2(new_n265), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n665), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n617), .B1(new_n686), .B2(KEYINPUT40), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  INV_X1    g509(.A(new_n625), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n681), .A2(new_n696), .A3(new_n672), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n626), .A2(KEYINPUT104), .A3(new_n672), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n667), .A2(new_n668), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n187), .ZN(G48));
  NAND3_X1  g517(.A1(new_n592), .A2(new_n593), .A3(new_n282), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n605), .A3(new_n595), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT105), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n705), .A2(new_n708), .A3(new_n605), .A4(new_n595), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n628), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n666), .A2(new_n613), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND3_X1  g528(.A1(new_n707), .A2(new_n618), .A3(new_n709), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n613), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n322), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n650), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G116), .ZN(G18));
  NOR3_X1   g534(.A1(new_n715), .A2(new_n497), .A3(new_n486), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n666), .A2(new_n659), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  AND4_X1   g537(.A1(new_n627), .A2(new_n707), .A3(new_n618), .A4(new_n709), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n278), .A2(new_n280), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n261), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n314), .B1(new_n726), .B2(new_n303), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n611), .B2(G472), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n613), .A3(new_n683), .A4(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n728), .A2(new_n613), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT106), .A3(new_n683), .A4(new_n724), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G122), .ZN(G24));
  AND2_X1   g549(.A1(new_n728), .A2(new_n659), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n699), .A2(new_n700), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n736), .A2(new_n737), .A3(new_n738), .A4(new_n716), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n728), .A2(new_n699), .A3(new_n659), .A4(new_n700), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT107), .B1(new_n740), .B2(new_n715), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  AOI211_X1 g557(.A(new_n617), .B(new_n564), .C1(new_n676), .C2(new_n499), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n615), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n701), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n666), .A2(new_n746), .A3(new_n613), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n320), .B2(KEYINPUT32), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n308), .A2(KEYINPUT108), .A3(new_n309), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n288), .A3(new_n751), .A4(new_n312), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n752), .A2(KEYINPUT42), .A3(new_n613), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n747), .A2(new_n748), .B1(new_n746), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n213), .ZN(G33));
  INV_X1    g569(.A(new_n673), .ZN(new_n756));
  INV_X1    g570(.A(new_n745), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n666), .A2(new_n613), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NAND2_X1  g573(.A1(new_n682), .A2(new_n696), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n612), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n763), .A3(new_n659), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT109), .Z(new_n767));
  OAI21_X1  g581(.A(new_n744), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n600), .B(KEYINPUT45), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(G469), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n596), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n595), .ZN(new_n773));
  AOI21_X1  g587(.A(KEYINPUT46), .B1(new_n771), .B2(new_n596), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n605), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n775), .A2(new_n684), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n769), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  XOR2_X1   g593(.A(new_n775), .B(KEYINPUT47), .Z(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n744), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n701), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(new_n322), .A3(new_n379), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G140), .ZN(G42));
  NOR3_X1   g599(.A1(new_n679), .A2(new_n604), .A3(new_n760), .ZN(new_n786));
  INV_X1    g600(.A(new_n692), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n705), .A2(new_n595), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n613), .B1(new_n788), .B2(KEYINPUT49), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(KEYINPUT49), .B2(new_n788), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n602), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n673), .A2(new_n668), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n701), .A2(new_n668), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n666), .B(new_n659), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n682), .A2(new_n659), .A3(new_n644), .A4(new_n671), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n692), .A2(new_n651), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n742), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n794), .A2(new_n742), .A3(KEYINPUT52), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n430), .A2(new_n463), .A3(new_n671), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n615), .A2(new_n744), .A3(new_n643), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n666), .A2(new_n803), .A3(new_n659), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n746), .A2(new_n736), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n758), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n758), .A2(new_n804), .A3(KEYINPUT111), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n608), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n666), .A2(new_n613), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n681), .A2(new_n696), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n644), .B2(new_n681), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n570), .A2(new_n814), .A3(new_n627), .A4(new_n602), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n616), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n812), .A2(new_n816), .A3(new_n817), .A4(new_n661), .ZN(new_n818));
  OAI22_X1  g632(.A1(new_n616), .A2(new_n815), .B1(new_n608), .B2(new_n660), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT110), .B1(new_n609), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n719), .A2(new_n734), .A3(new_n722), .A4(new_n712), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n754), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n801), .A2(new_n810), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n822), .ZN(new_n827));
  INV_X1    g641(.A(new_n754), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n827), .A2(new_n828), .A3(new_n821), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n801), .A4(new_n810), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT54), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT115), .ZN(new_n836));
  INV_X1    g650(.A(new_n492), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n762), .A2(new_n837), .A3(new_n732), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n716), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n833), .A2(new_n835), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n782), .A2(new_n710), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n787), .A2(new_n613), .A3(new_n837), .A4(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n490), .B1(new_n843), .B2(new_n626), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT51), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n707), .A2(new_n617), .A3(new_n709), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n679), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n838), .B(new_n849), .C1(new_n847), .C2(new_n848), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT50), .Z(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT113), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n841), .A2(new_n837), .A3(new_n762), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n736), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n843), .A2(new_n682), .A3(new_n625), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n781), .B1(new_n605), .B2(new_n788), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n838), .A2(new_n744), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n846), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n858), .A2(KEYINPUT114), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(new_n858), .B2(KEYINPUT114), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n846), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n856), .A3(new_n854), .A4(new_n851), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n752), .A2(new_n613), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n853), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n861), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n839), .A2(new_n836), .ZN(new_n871));
  AND2_X1   g685(.A1(KEYINPUT116), .A2(KEYINPUT48), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n867), .A2(new_n868), .A3(new_n872), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n845), .A2(new_n870), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(G952), .A2(G953), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n791), .B1(new_n874), .B2(new_n875), .ZN(G75));
  OR2_X1    g690(.A1(new_n541), .A2(new_n544), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(new_n506), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n282), .B1(new_n826), .B2(new_n830), .ZN(new_n880));
  AOI211_X1 g694(.A(KEYINPUT56), .B(new_n879), .C1(new_n880), .C2(new_n563), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT118), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n257), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n880), .A2(new_n563), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n885), .B2(KEYINPUT117), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n879), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n882), .A2(new_n884), .A3(new_n889), .ZN(G51));
  NAND2_X1  g704(.A1(new_n596), .A2(KEYINPUT57), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n833), .A2(new_n835), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n596), .A2(KEYINPUT57), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n592), .B(new_n593), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n880), .A2(G469), .A3(new_n770), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT119), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n883), .B1(new_n894), .B2(new_n896), .ZN(G54));
  NAND3_X1  g711(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(new_n473), .Z(new_n899));
  NOR2_X1   g713(.A1(new_n899), .A2(new_n883), .ZN(G60));
  XOR2_X1   g714(.A(new_n623), .B(KEYINPUT59), .Z(new_n901));
  NAND3_X1  g715(.A1(new_n833), .A2(new_n835), .A3(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n619), .A2(new_n620), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n902), .A2(new_n903), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n883), .ZN(G63));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n366), .B(KEYINPUT121), .Z(new_n908));
  NAND2_X1  g722(.A1(G217), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT60), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n831), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n907), .B1(new_n912), .B2(new_n883), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n910), .B1(new_n826), .B2(new_n830), .ZN(new_n914));
  OAI211_X1 g728(.A(KEYINPUT122), .B(new_n884), .C1(new_n914), .C2(new_n908), .ZN(new_n915));
  INV_X1    g729(.A(new_n657), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n914), .A2(KEYINPUT120), .A3(new_n916), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n913), .A2(new_n915), .A3(new_n919), .A4(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT123), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n922), .B1(new_n912), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(KEYINPUT123), .B1(new_n914), .B2(new_n908), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n925), .A2(new_n884), .A3(new_n917), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT124), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n923), .A2(new_n930), .A3(new_n927), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(G66));
  OAI21_X1  g746(.A(G953), .B1(new_n494), .B2(new_n503), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n822), .B1(new_n818), .B2(new_n820), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(G953), .ZN(new_n935));
  INV_X1    g749(.A(G898), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n877), .B1(new_n936), .B2(G953), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n935), .B(new_n937), .Z(G69));
  OAI21_X1  g752(.A(G953), .B1(new_n577), .B2(new_n669), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n794), .A2(new_n742), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n694), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT62), .Z(new_n942));
  NOR3_X1   g756(.A1(new_n322), .A2(new_n379), .A3(new_n745), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n943), .A2(new_n685), .A3(new_n814), .ZN(new_n944));
  AND4_X1   g758(.A1(new_n778), .A2(new_n942), .A3(new_n784), .A4(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n939), .B1(new_n945), .B2(G953), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n252), .B(new_n467), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n784), .A2(new_n940), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n866), .A2(new_n618), .A3(new_n683), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n777), .B1(new_n769), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n950), .A2(new_n828), .A3(new_n952), .A4(new_n758), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT125), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n949), .B1(new_n954), .B2(new_n257), .ZN(new_n955));
  OAI21_X1  g769(.A(G953), .B1(new_n669), .B2(G227), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(G72));
  XNOR2_X1  g771(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n958));
  AND2_X1   g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n958), .B(new_n959), .Z(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n954), .B2(new_n934), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n961), .A2(new_n265), .A3(new_n254), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n262), .B(new_n266), .C1(new_n293), .C2(new_n295), .ZN(new_n963));
  INV_X1    g777(.A(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT127), .Z(new_n966));
  NOR2_X1   g780(.A1(new_n832), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n960), .B1(new_n945), .B2(new_n934), .ZN(new_n968));
  INV_X1    g782(.A(new_n689), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n884), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n962), .A2(new_n967), .A3(new_n970), .ZN(G57));
endmodule


