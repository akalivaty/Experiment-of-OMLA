//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n977, new_n978;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n202), .B1(KEYINPUT23), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT25), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G176gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G169gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G183gat), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT64), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G183gat), .B2(G190gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n212), .A2(new_n215), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n205), .A2(new_n209), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT68), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n222), .B1(G183gat), .B2(G190gat), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n221), .A2(new_n223), .A3(new_n218), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n210), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n202), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n232), .A2(new_n207), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n204), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n220), .B1(new_n235), .B2(KEYINPUT25), .ZN(new_n236));
  INV_X1    g035(.A(new_n203), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n237), .B1(new_n232), .B2(KEYINPUT26), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(KEYINPUT26), .B2(new_n232), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n239), .A2(new_n210), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT27), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n241), .A2(G183gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n243));
  NOR4_X1   g042(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT28), .A4(G190gat), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n242), .B2(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n213), .A2(KEYINPUT27), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(G183gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT69), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n214), .A3(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n244), .B1(new_n250), .B2(KEYINPUT28), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n240), .B1(new_n251), .B2(KEYINPUT70), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT70), .ZN(new_n253));
  AOI211_X1 g052(.A(new_n253), .B(new_n244), .C1(new_n250), .C2(KEYINPUT28), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n236), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(G127gat), .B(G134gat), .Z(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G120gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n258));
  XOR2_X1   g057(.A(G113gat), .B(G120gat), .Z(new_n259));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260));
  XNOR2_X1  g059(.A(G127gat), .B(G134gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n255), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT28), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n247), .A2(new_n248), .A3(KEYINPUT69), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT69), .B1(new_n247), .B2(new_n248), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n267), .B1(new_n270), .B2(new_n214), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n253), .B1(new_n271), .B2(new_n244), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n251), .A2(KEYINPUT70), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n240), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n263), .A4(new_n236), .ZN(new_n275));
  INV_X1    g074(.A(G227gat), .ZN(new_n276));
  INV_X1    g075(.A(G233gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n266), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(G71gat), .B(G99gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n280), .B(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  OR2_X1    g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(KEYINPUT32), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n279), .A2(KEYINPUT72), .A3(KEYINPUT32), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n282), .B1(new_n279), .B2(KEYINPUT32), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n279), .A2(new_n283), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n278), .B1(new_n266), .B2(new_n275), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT34), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n295), .A2(new_n294), .A3(new_n296), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  AOI22_X1  g102(.A1(new_n287), .A2(new_n288), .B1(new_n291), .B2(new_n290), .ZN(new_n304));
  NOR3_X1   g103(.A1(new_n300), .A2(new_n297), .A3(new_n298), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT36), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n303), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n302), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n305), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT36), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  XOR2_X1   g110(.A(G8gat), .B(G36gat), .Z(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(KEYINPUT75), .ZN(new_n313));
  XNOR2_X1  g112(.A(G64gat), .B(G92gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G226gat), .A2(G233gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n235), .A2(KEYINPUT25), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n205), .A2(new_n209), .A3(new_n219), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n239), .A2(new_n210), .ZN(new_n321));
  INV_X1    g120(.A(new_n244), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n268), .A2(new_n269), .A3(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(new_n267), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(new_n253), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n320), .B1(new_n325), .B2(new_n273), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n317), .B1(new_n326), .B2(KEYINPUT29), .ZN(new_n327));
  XNOR2_X1  g126(.A(G197gat), .B(G204gat), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  INV_X1    g128(.A(G211gat), .ZN(new_n330));
  INV_X1    g129(.A(G218gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(G211gat), .B(G218gat), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n328), .A3(new_n332), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n317), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n255), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n327), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT29), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n339), .B1(new_n255), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n326), .B2(new_n317), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n255), .A2(KEYINPUT74), .A3(new_n339), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n316), .B(new_n341), .C1(new_n347), .C2(new_n338), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n341), .B1(new_n347), .B2(new_n338), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n315), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n255), .A2(KEYINPUT74), .A3(new_n339), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT74), .B1(new_n255), .B2(new_n339), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n327), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n338), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n316), .A4(new_n341), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n350), .A2(new_n352), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(G141gat), .A2(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT2), .ZN(new_n362));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  INV_X1    g164(.A(G155gat), .ZN(new_n366));
  INV_X1    g165(.A(G162gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n361), .A2(KEYINPUT76), .A3(new_n363), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n371));
  AND2_X1   g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n368), .A2(new_n374), .A3(new_n365), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n370), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AND2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT77), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n362), .B2(new_n377), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n369), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT3), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n369), .C1(new_n376), .C2(new_n380), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n384), .A3(new_n263), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT5), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n258), .A2(new_n262), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n365), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n390), .A2(KEYINPUT77), .B1(KEYINPUT2), .B2(new_n365), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n391), .A2(new_n370), .A3(new_n375), .A4(new_n373), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n389), .A2(new_n369), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT4), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT4), .B1(new_n381), .B2(new_n263), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT78), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n369), .C1(new_n376), .C2(new_n380), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n398), .A2(new_n399), .A3(new_n389), .A4(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n395), .A2(new_n397), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n389), .A4(new_n401), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n399), .B1(new_n381), .B2(new_n263), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n405), .A2(new_n385), .A3(new_n387), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n263), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n387), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n386), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G1gat), .B(G29gat), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(KEYINPUT6), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n413), .A2(KEYINPUT82), .A3(KEYINPUT6), .A4(new_n418), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n403), .A2(new_n388), .B1(new_n407), .B2(new_n411), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT6), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT80), .B1(new_n413), .B2(new_n418), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT80), .ZN(new_n427));
  AOI211_X1 g226(.A(new_n427), .B(new_n417), .C1(new_n404), .C2(new_n412), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n423), .B1(KEYINPUT81), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n425), .C1(new_n426), .C2(new_n428), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n359), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT84), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT3), .B1(new_n338), .B2(new_n342), .ZN(new_n435));
  INV_X1    g234(.A(new_n381), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G228gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n384), .A2(new_n342), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n356), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n435), .B1(new_n398), .B2(new_n401), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n440), .B2(new_n356), .ZN(new_n445));
  AOI211_X1 g244(.A(KEYINPUT83), .B(new_n338), .C1(new_n384), .C2(new_n342), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n443), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n442), .B1(new_n447), .B2(new_n439), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(G22gat), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(new_n442), .C1(new_n447), .C2(new_n439), .ZN(new_n451));
  XNOR2_X1  g250(.A(G78gat), .B(G106gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(KEYINPUT31), .B(G50gat), .ZN(new_n453));
  XOR2_X1   g252(.A(new_n452), .B(new_n453), .Z(new_n454));
  AND4_X1   g253(.A1(new_n434), .A2(new_n449), .A3(new_n451), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(KEYINPUT84), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n456), .A2(new_n454), .B1(new_n449), .B2(new_n451), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OAI22_X1  g257(.A1(new_n308), .A2(new_n311), .B1(new_n433), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n387), .B1(new_n403), .B2(new_n385), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT39), .B1(new_n409), .B2(new_n410), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n417), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n403), .A2(new_n385), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT85), .B(KEYINPUT39), .Z(new_n465));
  AND3_X1   g264(.A1(new_n464), .A2(new_n410), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n460), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n464), .A2(new_n410), .ZN(new_n468));
  INV_X1    g267(.A(new_n462), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n460), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n461), .A2(new_n465), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n470), .A2(new_n417), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n413), .A2(new_n418), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n467), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n359), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n458), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n351), .A2(KEYINPUT37), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(KEYINPUT88), .A3(new_n315), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n357), .A2(new_n480), .A3(new_n341), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n316), .B1(new_n351), .B2(KEYINPUT37), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(KEYINPUT88), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT38), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n425), .A2(new_n474), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n486), .A2(new_n348), .A3(new_n421), .A4(new_n422), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n338), .B1(new_n327), .B2(new_n340), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n347), .A2(new_n338), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n488), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n347), .A2(KEYINPUT87), .A3(new_n338), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT37), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT38), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n481), .A2(new_n495), .A3(new_n315), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n487), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n477), .B1(new_n485), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n309), .A2(new_n458), .A3(new_n310), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(new_n433), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n486), .A2(new_n421), .A3(new_n422), .ZN(new_n503));
  OR3_X1    g302(.A1(new_n359), .A2(new_n503), .A3(KEYINPUT35), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n309), .A2(new_n458), .A3(new_n310), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI22_X1  g305(.A1(new_n459), .A2(new_n499), .B1(new_n502), .B2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(G190gat), .B(G218gat), .Z(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(G99gat), .B(G106gat), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512));
  INV_X1    g311(.A(G85gat), .ZN(new_n513));
  INV_X1    g312(.A(G92gat), .ZN(new_n514));
  AOI22_X1  g313(.A1(KEYINPUT8), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT102), .Z(new_n516));
  INV_X1    g315(.A(KEYINPUT7), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n517), .B1(G85gat), .B2(G92gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT100), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(G85gat), .A3(G92gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT101), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n511), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n516), .A2(new_n522), .A3(new_n511), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G43gat), .B(G50gat), .Z(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G29gat), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n531), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT14), .B(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n536), .A2(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(KEYINPUT89), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n528), .A2(new_n529), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n540), .B(KEYINPUT90), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n530), .A2(new_n535), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n545));
  AOI21_X1  g344(.A(new_n527), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n539), .A2(new_n543), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT17), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n547), .B2(KEYINPUT17), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n546), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n547), .B2(new_n526), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT103), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(KEYINPUT103), .B(new_n552), .C1(new_n547), .C2(new_n526), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n509), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT99), .ZN(new_n561));
  XNOR2_X1  g360(.A(G134gat), .B(G162gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n551), .A2(new_n557), .A3(new_n509), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n563), .ZN(new_n566));
  INV_X1    g365(.A(new_n564), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(new_n558), .ZN(new_n568));
  XNOR2_X1  g367(.A(G15gat), .B(G22gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G1gat), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT16), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n571), .A2(new_n572), .B1(new_n573), .B2(new_n569), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n572), .B2(new_n571), .ZN(new_n575));
  INV_X1    g374(.A(G8gat), .ZN(new_n576));
  OR3_X1    g375(.A1(new_n575), .A2(KEYINPUT93), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(G8gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n575), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G64gat), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n583), .A2(G57gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(G57gat), .ZN(new_n585));
  AND2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  OAI22_X1  g385(.A1(new_n584), .A2(new_n585), .B1(KEYINPUT9), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G71gat), .B(G78gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT21), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT98), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n582), .A2(new_n593), .A3(new_n590), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(new_n366), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n592), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n589), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT97), .B(KEYINPUT21), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(G231gat), .A3(G233gat), .ZN(new_n606));
  INV_X1    g405(.A(G127gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n603), .A2(new_n608), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n606), .B2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n602), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  INV_X1    g413(.A(new_n602), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n598), .A2(new_n613), .A3(new_n616), .A4(new_n600), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n565), .A2(new_n568), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT104), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT104), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n565), .A2(new_n568), .A3(new_n620), .A4(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  AOI22_X1  g424(.A1(new_n544), .A2(new_n545), .B1(new_n577), .B2(new_n581), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n549), .B2(new_n550), .ZN(new_n627));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT95), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n544), .A2(new_n581), .A3(new_n577), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT18), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT96), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n632), .A2(KEYINPUT96), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g436(.A1(new_n627), .A2(KEYINPUT18), .A3(new_n630), .A4(new_n631), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n582), .A2(new_n547), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n631), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n629), .B(KEYINPUT13), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G113gat), .B(G141gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(G197gat), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT11), .B(G169gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n638), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n633), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n642), .A3(new_n638), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n637), .A2(new_n649), .B1(new_n651), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(G230gat), .A2(G233gat), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n526), .A2(new_n603), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n524), .A2(new_n589), .A3(new_n525), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n657), .A2(new_n656), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n657), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n654), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(G176gat), .B(G204gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  OR2_X1    g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n658), .A2(new_n659), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n653), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(new_n665), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n661), .A2(new_n654), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT105), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n625), .A2(new_n652), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n507), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT106), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n507), .A2(new_n677), .A3(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n429), .A2(KEYINPUT81), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n421), .A2(new_n422), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n680), .A2(new_n432), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  AND3_X1   g484(.A1(new_n350), .A2(new_n352), .A3(new_n358), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n686), .B1(new_n676), .B2(new_n678), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n576), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n690), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n686), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT107), .B1(new_n679), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696));
  INV_X1    g495(.A(new_n694), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n696), .B(new_n697), .C1(new_n676), .C2(new_n678), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n692), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI211_X1 g500(.A(new_n686), .B(new_n693), .C1(new_n676), .C2(new_n678), .ZN(new_n702));
  OAI22_X1  g501(.A1(new_n702), .A2(KEYINPUT42), .B1(new_n576), .B2(new_n687), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n695), .A2(new_n698), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT108), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n679), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n309), .A2(new_n310), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n707), .A2(G15gat), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n307), .B1(new_n303), .B2(new_n306), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n309), .A2(KEYINPUT36), .A3(new_n310), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n707), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n709), .A2(new_n713), .ZN(G1326gat));
  OR2_X1    g513(.A1(new_n455), .A2(new_n457), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n679), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT43), .B(G22gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n682), .A2(new_n686), .ZN(new_n720));
  AOI22_X1  g519(.A1(new_n710), .A2(new_n711), .B1(new_n720), .B2(new_n715), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n715), .B1(new_n359), .B2(new_n475), .ZN(new_n722));
  INV_X1    g521(.A(new_n481), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n723), .B1(KEYINPUT88), .B2(new_n483), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n478), .A2(new_n315), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT88), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n495), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n480), .B1(new_n491), .B2(new_n492), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n348), .B(new_n503), .C1(new_n729), .C2(new_n496), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n722), .B1(new_n728), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT35), .B1(new_n720), .B2(new_n505), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n359), .A2(new_n503), .A3(KEYINPUT35), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n501), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n721), .A2(new_n731), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n565), .A2(new_n568), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n719), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n507), .A2(KEYINPUT44), .A3(new_n736), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n652), .A2(new_n620), .A3(new_n673), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n738), .A2(new_n739), .A3(new_n743), .A4(new_n740), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n683), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G29gat), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n735), .A2(new_n737), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n747), .A2(new_n531), .A3(new_n683), .A4(new_n740), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n746), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1328gat));
  NAND3_X1  g553(.A1(new_n742), .A2(new_n359), .A3(new_n744), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G36gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n747), .A2(new_n534), .A3(new_n359), .A4(new_n740), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT46), .Z(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(new_n758), .A3(KEYINPUT111), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1329gat));
  AND2_X1   g562(.A1(new_n747), .A2(new_n740), .ZN(new_n764));
  INV_X1    g563(.A(G43gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n708), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n712), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n742), .A2(new_n768), .A3(new_n744), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n767), .B1(new_n769), .B2(G43gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n741), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n765), .B1(new_n773), .B2(new_n768), .ZN(new_n774));
  OAI22_X1  g573(.A1(new_n770), .A2(KEYINPUT47), .B1(new_n772), .B2(new_n774), .ZN(G1330gat));
  INV_X1    g574(.A(G50gat), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n764), .A2(new_n776), .A3(new_n715), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n742), .A2(new_n715), .A3(new_n744), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(G50gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n776), .B1(new_n773), .B2(new_n715), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n779), .A2(KEYINPUT48), .B1(new_n781), .B2(new_n782), .ZN(G1331gat));
  INV_X1    g582(.A(new_n652), .ZN(new_n784));
  INV_X1    g583(.A(new_n673), .ZN(new_n785));
  NOR4_X1   g584(.A1(new_n735), .A2(new_n784), .A3(new_n625), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n683), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n359), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n790));
  XOR2_X1   g589(.A(KEYINPUT49), .B(G64gat), .Z(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n789), .B2(new_n791), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n793), .A3(new_n766), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n786), .A2(new_n768), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n793), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n796), .B(new_n797), .Z(G1334gat));
  NAND2_X1  g597(.A1(new_n786), .A2(new_n715), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n620), .A3(new_n785), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n738), .A2(new_n739), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G85gat), .B1(new_n802), .B2(new_n682), .ZN(new_n803));
  INV_X1    g602(.A(new_n620), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n507), .A2(new_n652), .A3(new_n804), .A4(new_n736), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n683), .A2(new_n513), .A3(new_n673), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  NOR3_X1   g609(.A1(new_n785), .A2(G92gat), .A3(new_n686), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n738), .A2(new_n739), .A3(new_n359), .A4(new_n801), .ZN(new_n812));
  AOI22_X1  g611(.A1(new_n807), .A2(new_n811), .B1(G92gat), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT52), .Z(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n802), .B2(new_n712), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n785), .A2(new_n708), .A3(G99gat), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n808), .B2(new_n816), .ZN(G1338gat));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n785), .A2(new_n458), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n807), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(G106gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n458), .A2(new_n823), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n738), .A2(new_n739), .A3(new_n801), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n818), .A2(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n820), .B1(new_n824), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g629(.A(new_n819), .B(new_n828), .C1(new_n822), .C2(new_n823), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(G1339gat));
  AOI21_X1  g631(.A(new_n630), .B1(new_n627), .B2(new_n631), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n640), .A2(new_n641), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n646), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(KEYINPUT114), .B(new_n646), .C1(new_n833), .C2(new_n834), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n636), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n649), .B1(new_n840), .B2(new_n634), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n841), .A3(new_n673), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n665), .B1(new_n660), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n668), .A2(KEYINPUT54), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n667), .A2(new_n653), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n847), .A2(new_n848), .B1(new_n671), .B2(new_n669), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT55), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n842), .B(new_n737), .C1(new_n652), .C2(new_n851), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n839), .A2(new_n841), .A3(new_n849), .A4(new_n850), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n620), .B1(new_n853), .B2(new_n736), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n622), .A2(new_n624), .A3(new_n785), .ZN(new_n855));
  AOI22_X1  g654(.A1(new_n852), .A2(new_n854), .B1(new_n855), .B2(new_n652), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n505), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n682), .A2(new_n359), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n784), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n673), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g662(.A1(new_n859), .A2(new_n620), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g664(.A1(new_n859), .A2(new_n736), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(G134gat), .ZN(new_n867));
  XOR2_X1   g666(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(G134gat), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(G1343gat));
  NAND2_X1  g671(.A1(new_n712), .A2(new_n858), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n856), .A2(new_n458), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n784), .ZN(new_n875));
  NOR2_X1   g674(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT57), .B1(new_n856), .B2(new_n458), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n854), .A2(new_n852), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n622), .A2(new_n652), .A3(new_n624), .A4(new_n785), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n458), .A2(KEYINPUT57), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n873), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(G141gat), .A3(new_n784), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n877), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(KEYINPUT116), .A2(KEYINPUT58), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1344gat));
  INV_X1    g687(.A(G148gat), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n889), .A3(new_n673), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT59), .B(new_n889), .C1(new_n884), .C2(new_n673), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT118), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n880), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n893), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n882), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n873), .B(KEYINPUT117), .Z(new_n898));
  NAND4_X1  g697(.A1(new_n878), .A2(new_n897), .A3(new_n673), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n892), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n890), .B1(new_n891), .B2(new_n900), .ZN(G1345gat));
  AOI21_X1  g700(.A(KEYINPUT119), .B1(new_n874), .B2(new_n620), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(G155gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n874), .A2(KEYINPUT119), .A3(new_n620), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n804), .A2(new_n366), .ZN(new_n905));
  AOI22_X1  g704(.A1(new_n903), .A2(new_n904), .B1(new_n884), .B2(new_n905), .ZN(G1346gat));
  NAND3_X1  g705(.A1(new_n878), .A2(new_n883), .A3(new_n736), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(KEYINPUT120), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n878), .A2(new_n883), .A3(new_n909), .A4(new_n736), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(G162gat), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n874), .A2(new_n367), .A3(new_n736), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT121), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n911), .A2(new_n915), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n683), .A2(new_n686), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n857), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n652), .ZN(new_n920));
  XOR2_X1   g719(.A(new_n920), .B(G169gat), .Z(G1348gat));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n785), .ZN(new_n922));
  MUX2_X1   g721(.A(G176gat), .B(new_n206), .S(new_n922), .Z(G1349gat));
  INV_X1    g722(.A(KEYINPUT60), .ZN(new_n924));
  OR3_X1    g723(.A1(new_n919), .A2(new_n270), .A3(new_n804), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n213), .B1(new_n919), .B2(new_n804), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT122), .B(new_n924), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n929));
  AND4_X1   g728(.A1(new_n928), .A2(new_n925), .A3(new_n926), .A4(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n927), .A2(new_n930), .ZN(G1350gat));
  OAI22_X1  g730(.A1(new_n919), .A2(new_n737), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n932));
  NAND2_X1  g731(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n932), .B(new_n933), .ZN(G1351gat));
  NAND3_X1  g733(.A1(new_n712), .A2(new_n715), .A3(new_n918), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n856), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n784), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT57), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n881), .B2(new_n715), .ZN(new_n940));
  INV_X1    g739(.A(new_n882), .ZN(new_n941));
  AOI22_X1  g740(.A1(new_n854), .A2(new_n852), .B1(new_n880), .B2(new_n893), .ZN(new_n942));
  INV_X1    g741(.A(new_n896), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n938), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n878), .A2(new_n897), .A3(KEYINPUT123), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n712), .A2(new_n918), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(new_n652), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n937), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT124), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n951), .B(new_n952), .ZN(G1352gat));
  XNOR2_X1  g752(.A(KEYINPUT125), .B(G204gat), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n948), .A2(new_n785), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n954), .B1(new_n947), .B2(new_n955), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n936), .A2(new_n673), .A3(new_n954), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n957), .B(KEYINPUT62), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT126), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n957), .B(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  INV_X1    g761(.A(new_n955), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n963), .B1(new_n945), .B2(new_n946), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n961), .B(new_n962), .C1(new_n954), .C2(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n959), .A2(new_n965), .ZN(G1353gat));
  NAND3_X1  g765(.A1(new_n936), .A2(new_n330), .A3(new_n620), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n948), .A2(new_n804), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n878), .A2(new_n897), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g773(.A(KEYINPUT127), .B(new_n967), .C1(new_n970), .C2(new_n971), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1354gat));
  AOI21_X1  g775(.A(G218gat), .B1(new_n936), .B2(new_n736), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n948), .A2(new_n331), .A3(new_n737), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n947), .B2(new_n978), .ZN(G1355gat));
endmodule


