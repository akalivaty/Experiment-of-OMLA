//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1327, new_n1329, new_n1330, new_n1331, new_n1332, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1411, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n207), .B2(new_n220), .C1(new_n202), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n214), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OR2_X1    g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT66), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n229), .A2(new_n212), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n206), .A2(new_n207), .ZN(new_n231));
  AOI22_X1  g0031(.A1(new_n226), .A2(KEYINPUT1), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g0032(.A1(new_n218), .A2(new_n228), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND3_X1  g0049(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n250), .A2(new_n251), .A3(new_n229), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(new_n250), .B2(new_n229), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n202), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n212), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n255), .B1(new_n256), .B2(new_n257), .C1(new_n259), .C2(new_n207), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n254), .A2(new_n260), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT11), .ZN(new_n262));
  INV_X1    g0062(.A(G13), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n265), .A2(G68), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT12), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(KEYINPUT74), .A3(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n267), .B(new_n270), .C1(new_n269), .C2(new_n268), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n211), .A2(G13), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n212), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n250), .A2(new_n229), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n212), .A2(G1), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n275), .A2(G68), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n261), .A2(KEYINPUT11), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n262), .A2(new_n271), .A3(new_n278), .A4(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT14), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n220), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n235), .A2(G1698), .ZN(new_n286));
  AND2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(G33), .A2(G97), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G41), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  AOI21_X1  g0097(.A(G1), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n298), .A2(new_n293), .A3(G274), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n293), .A2(G238), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n283), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n293), .B1(new_n289), .B2(new_n290), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n299), .A2(new_n301), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT13), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n282), .B(G169), .C1(new_n303), .C2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n295), .A2(new_n302), .A3(new_n283), .ZN(new_n308));
  OAI21_X1  g0108(.A(KEYINPUT13), .B1(new_n304), .B2(new_n305), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G179), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n309), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n282), .B1(new_n312), .B2(G169), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT75), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n303), .A2(new_n306), .ZN(new_n315));
  INV_X1    g0115(.A(G169), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT14), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT75), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n317), .A2(new_n318), .A3(new_n310), .A4(new_n307), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n281), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n312), .A2(G200), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n315), .A2(G190), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n281), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT3), .B(G33), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n327), .A2(G222), .A3(new_n284), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT67), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n328), .B(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n327), .A2(G1698), .ZN(new_n331));
  INV_X1    g0131(.A(G223), .ZN(new_n332));
  OAI22_X1  g0132(.A1(new_n331), .A2(new_n332), .B1(new_n257), .B2(new_n327), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n293), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n293), .A2(new_n300), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n299), .B1(new_n220), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n316), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n208), .A2(G20), .B1(G150), .B2(new_n258), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT8), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(G58), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT70), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT69), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n256), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n254), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n252), .A2(new_n253), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n265), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n277), .A2(G50), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(G50), .B2(new_n265), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  INV_X1    g0155(.A(new_n337), .ZN(new_n356));
  OR2_X1    g0156(.A1(new_n328), .A2(new_n329), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n328), .A2(new_n329), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n333), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n355), .B(new_n356), .C1(new_n359), .C2(new_n293), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n338), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n343), .A2(new_n346), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n339), .B1(new_n363), .B2(new_n256), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n352), .B1(new_n364), .B2(new_n254), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n362), .B1(new_n365), .B2(KEYINPUT9), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n354), .A2(KEYINPUT73), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G200), .B1(new_n335), .B2(new_n337), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n348), .A2(new_n353), .A3(KEYINPUT9), .ZN(new_n371));
  OAI211_X1 g0171(.A(G190), .B(new_n356), .C1(new_n359), .C2(new_n293), .ZN(new_n372));
  AND3_X1   g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT10), .ZN(new_n374));
  AND3_X1   g0174(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n369), .B2(new_n373), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n361), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n343), .A2(new_n346), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n277), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n379), .A2(new_n350), .B1(new_n265), .B2(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(new_n274), .ZN(new_n381));
  OR2_X1    g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NAND2_X1  g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n383), .ZN(new_n384));
  NOR3_X1   g0184(.A1(new_n287), .A2(new_n288), .A3(G20), .ZN(new_n385));
  OR2_X1    g0185(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n384), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n203), .A2(new_n205), .A3(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G20), .B1(G159), .B2(new_n258), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n381), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n382), .A2(new_n212), .A3(new_n383), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n397), .B2(new_n388), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n393), .B(KEYINPUT16), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n380), .B1(new_n396), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n220), .A2(G1698), .ZN(new_n403));
  OAI221_X1 g0203(.A(new_n403), .B1(G223), .B2(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n293), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n293), .A2(G232), .A3(new_n300), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n299), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G179), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n406), .B2(new_n408), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(KEYINPUT18), .B1(new_n402), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(G190), .ZN(new_n415));
  OAI21_X1  g0215(.A(G200), .B1(new_n406), .B2(new_n408), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n402), .A2(KEYINPUT17), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n397), .A2(new_n386), .A3(new_n387), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n202), .B1(new_n419), .B2(new_n384), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n392), .A2(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n258), .A2(G159), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n395), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n274), .A3(new_n401), .ZN(new_n425));
  INV_X1    g0225(.A(new_n350), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n276), .B1(new_n343), .B2(new_n346), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n363), .B2(new_n273), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n425), .A2(new_n428), .A3(new_n415), .A4(new_n416), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n428), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(new_n412), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n414), .A2(new_n418), .A3(new_n431), .A4(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n287), .A2(new_n288), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n235), .A2(new_n284), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n221), .A2(G1698), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n294), .B1(new_n327), .B2(G107), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(G244), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n299), .B1(new_n442), .B2(new_n336), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(G200), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(new_n443), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(KEYINPUT71), .A3(G190), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n259), .A2(KEYINPUT72), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n342), .A2(new_n344), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n259), .A2(KEYINPUT72), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g0251(.A(KEYINPUT15), .B(G87), .ZN(new_n452));
  OAI221_X1 g0252(.A(new_n451), .B1(new_n212), .B2(new_n257), .C1(new_n256), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n274), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n276), .A2(new_n257), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n275), .A2(new_n455), .B1(new_n257), .B2(new_n273), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n445), .A2(new_n447), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(KEYINPUT71), .B1(new_n446), .B2(G190), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n454), .A2(new_n456), .B1(new_n444), .B2(new_n316), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n446), .A2(new_n355), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n459), .A2(new_n462), .ZN(new_n463));
  NOR4_X1   g0263(.A1(new_n326), .A2(new_n377), .A3(new_n435), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT85), .ZN(new_n465));
  OAI211_X1 g0265(.A(G257), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT83), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT83), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n327), .A2(new_n468), .A3(G257), .A4(new_n284), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n327), .A2(G264), .A3(G1698), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n436), .A2(G303), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n294), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n211), .B(G45), .C1(new_n296), .C2(KEYINPUT5), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(KEYINPUT79), .ZN(new_n475));
  INV_X1    g0275(.A(G274), .ZN(new_n476));
  INV_X1    g0276(.A(new_n229), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(new_n292), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n297), .A2(G1), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT5), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G41), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n296), .A2(KEYINPUT5), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n475), .A2(new_n478), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(new_n484), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G270), .A3(new_n293), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n473), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G200), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n294), .B2(new_n472), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G190), .ZN(new_n493));
  INV_X1    g0293(.A(G116), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n250), .A2(new_n229), .B1(G20), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  INV_X1    g0296(.A(G97), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n212), .C1(G33), .C2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT20), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n495), .A2(KEYINPUT20), .A3(new_n498), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n211), .A2(G33), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G116), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n212), .A2(G116), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n275), .A2(new_n505), .B1(new_n264), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n491), .A2(new_n493), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n491), .A2(new_n493), .A3(KEYINPUT84), .A4(new_n509), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT21), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n495), .A2(KEYINPUT20), .A3(new_n498), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n499), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n264), .A2(new_n506), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n381), .A2(new_n265), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n519), .B2(new_n504), .ZN(new_n520));
  OAI21_X1  g0320(.A(G169), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n515), .B1(new_n492), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n316), .B1(new_n502), .B2(new_n507), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n490), .A2(new_n523), .A3(KEYINPUT21), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n492), .A2(G179), .A3(new_n508), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n465), .B1(new_n514), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n514), .A2(new_n465), .A3(new_n526), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n389), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(KEYINPUT77), .B(G107), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n497), .A2(new_n534), .A3(KEYINPUT6), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G97), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(G20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n258), .A2(G77), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n531), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n274), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n265), .A2(G97), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n349), .A2(new_n265), .A3(new_n503), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n545), .B1(new_n547), .B2(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n442), .A2(G1698), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(KEYINPUT4), .C1(new_n288), .C2(new_n287), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT78), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT78), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n327), .A2(new_n553), .A3(KEYINPUT4), .A4(new_n550), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G250), .B(G1698), .C1(new_n287), .C2(new_n288), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n284), .A2(G244), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n382), .B2(new_n383), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n496), .B(new_n556), .C1(new_n558), .C2(KEYINPUT4), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n294), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n486), .A2(G257), .A3(new_n293), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n485), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n316), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n550), .B1(new_n287), .B2(new_n288), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n566), .A2(new_n567), .B1(G33), .B2(G283), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n568), .A2(new_n552), .A3(new_n556), .A4(new_n554), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n562), .B1(new_n569), .B2(new_n294), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n355), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n549), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n549), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT80), .B1(new_n564), .B2(G200), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT80), .ZN(new_n575));
  INV_X1    g0375(.A(G200), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n570), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n570), .A2(KEYINPUT81), .A3(G190), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT81), .B1(new_n570), .B2(G190), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n572), .B1(new_n578), .B2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(G250), .B(new_n284), .C1(new_n287), .C2(new_n288), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT88), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g0386(.A(KEYINPUT89), .B(G294), .Z(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G33), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n327), .A2(KEYINPUT88), .A3(G250), .A4(new_n284), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n327), .A2(G257), .A3(G1698), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n586), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n294), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n486), .A2(G264), .A3(new_n293), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n485), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(G169), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT90), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n486), .A2(KEYINPUT90), .A3(G264), .A4(new_n293), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n591), .A2(new_n294), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(G179), .A3(new_n485), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT23), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n212), .B2(G107), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n534), .A2(KEYINPUT23), .A3(G20), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(G33), .A2(G116), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n212), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n212), .B(G87), .C1(new_n287), .C2(new_n288), .ZN(new_n614));
  NOR2_X1   g0414(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n613), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n327), .A2(new_n212), .A3(G87), .A4(new_n615), .ZN(new_n618));
  AOI211_X1 g0418(.A(KEYINPUT24), .B(new_n611), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT24), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n614), .A2(new_n616), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(new_n618), .A3(new_n612), .ZN(new_n622));
  INV_X1    g0422(.A(new_n611), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n620), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n274), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n273), .A2(new_n534), .ZN(new_n626));
  XNOR2_X1  g0426(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n626), .B(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(G107), .B2(new_n547), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n603), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(G200), .B1(new_n601), .B2(new_n485), .ZN(new_n632));
  INV_X1    g0432(.A(G190), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n592), .A2(new_n633), .A3(new_n595), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n625), .B(new_n629), .C1(new_n632), .C2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n221), .A2(new_n284), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n442), .A2(G1698), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(new_n287), .C2(new_n288), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n608), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n294), .ZN(new_n640));
  INV_X1    g0440(.A(G250), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n297), .B2(G1), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n211), .A2(new_n476), .A3(G45), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n293), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT82), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n293), .B1(new_n638), .B2(new_n608), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT82), .ZN(new_n647));
  INV_X1    g0447(.A(new_n644), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n316), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n647), .B1(new_n646), .B2(new_n648), .ZN(new_n651));
  NOR2_X1   g0451(.A1(G238), .A2(G1698), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n652), .B1(new_n442), .B2(G1698), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n609), .B1(new_n653), .B2(new_n327), .ZN(new_n654));
  OAI211_X1 g0454(.A(KEYINPUT82), .B(new_n644), .C1(new_n654), .C2(new_n293), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n651), .A2(new_n655), .A3(new_n355), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT19), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n212), .B1(new_n290), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(G87), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n659), .A2(new_n497), .A3(new_n534), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n212), .B(G68), .C1(new_n287), .C2(new_n288), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n657), .B1(new_n256), .B2(new_n497), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n274), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n273), .A2(new_n452), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n665), .B(new_n666), .C1(new_n546), .C2(new_n452), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n650), .A2(new_n656), .A3(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(G200), .B1(new_n645), .B2(new_n649), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n651), .A2(new_n655), .A3(G190), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n349), .A2(G87), .A3(new_n265), .A4(new_n503), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n671), .A2(new_n665), .A3(new_n666), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n631), .A2(new_n635), .A3(new_n668), .A4(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n583), .A2(new_n674), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n464), .A2(new_n530), .A3(new_n675), .ZN(G372));
  INV_X1    g0476(.A(KEYINPUT93), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n432), .A2(new_n433), .A3(new_n412), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n433), .B1(new_n432), .B2(new_n412), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n414), .A2(KEYINPUT93), .A3(new_n434), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n462), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n320), .B1(new_n323), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n418), .A2(new_n431), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT73), .B1(new_n354), .B2(new_n367), .ZN(new_n687));
  AOI211_X1 g0487(.A(new_n362), .B(KEYINPUT9), .C1(new_n348), .C2(new_n353), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n690));
  OAI21_X1  g0490(.A(KEYINPUT10), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n369), .A2(new_n373), .A3(new_n374), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(new_n361), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n549), .A2(new_n565), .A3(new_n571), .ZN(new_n696));
  INV_X1    g0496(.A(new_n581), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n579), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n575), .B1(new_n570), .B2(new_n576), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n564), .A2(KEYINPUT80), .A3(G200), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n549), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n696), .B1(new_n698), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n640), .A2(new_n644), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n656), .B(new_n667), .C1(G169), .C2(new_n704), .ZN(new_n705));
  OAI211_X1 g0505(.A(new_n670), .B(new_n672), .C1(new_n576), .C2(new_n704), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n599), .A2(new_n600), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n592), .A2(new_n485), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n594), .B1(new_n294), .B2(new_n591), .ZN(new_n709));
  AOI22_X1  g0509(.A1(new_n708), .A2(new_n576), .B1(new_n709), .B2(new_n633), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n705), .B(new_n706), .C1(new_n710), .C2(new_n630), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n526), .A2(new_n631), .A3(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n597), .A2(new_n602), .B1(new_n625), .B2(new_n629), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT91), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n702), .A2(new_n712), .A3(new_n714), .A4(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n705), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n696), .A2(new_n668), .A3(new_n673), .A4(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT26), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n706), .A2(new_n705), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(new_n572), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n718), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n464), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n695), .A2(new_n728), .ZN(G369));
  OR3_X1    g0529(.A1(new_n272), .A2(KEYINPUT27), .A3(G20), .ZN(new_n730));
  OAI21_X1  g0530(.A(KEYINPUT27), .B1(new_n272), .B2(G20), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(G213), .A3(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G343), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n630), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n631), .A2(new_n635), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n715), .A2(new_n734), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n734), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n509), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n528), .B2(new_n529), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n716), .A2(new_n740), .ZN(new_n742));
  OAI211_X1 g0542(.A(G330), .B(new_n738), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n631), .A2(new_n635), .A3(new_n716), .A4(new_n739), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n715), .A2(new_n739), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT94), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n744), .A2(KEYINPUT94), .A3(new_n745), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n743), .B1(new_n746), .B2(new_n748), .ZN(G399));
  OR2_X1    g0549(.A1(new_n660), .A2(G116), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  INV_X1    g0551(.A(new_n215), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G41), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n751), .A2(new_n753), .A3(new_n211), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n754), .B1(new_n231), .B2(new_n753), .ZN(new_n755));
  XOR2_X1   g0555(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  AOI21_X1  g0556(.A(new_n734), .B1(new_n718), .B2(new_n726), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(KEYINPUT29), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT98), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n670), .A2(new_n672), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n576), .B1(new_n651), .B2(new_n655), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n656), .A2(new_n667), .ZN(new_n762));
  AOI21_X1  g0562(.A(G169), .B1(new_n651), .B2(new_n655), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n759), .B(new_n720), .C1(new_n764), .C2(new_n572), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n544), .A2(new_n548), .B1(new_n570), .B2(new_n355), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n767), .A2(new_n668), .A3(new_n673), .A4(new_n565), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n759), .B1(new_n768), .B2(new_n720), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n724), .A2(new_n572), .A3(new_n723), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n766), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n724), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n772), .B(new_n635), .C1(new_n715), .C2(new_n716), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n705), .B1(new_n773), .B2(new_n583), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n739), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT99), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n715), .A2(new_n716), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n711), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n719), .B1(new_n779), .B2(new_n702), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n720), .B1(new_n764), .B2(new_n572), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(KEYINPUT98), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n772), .A2(new_n696), .A3(KEYINPUT26), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n782), .A2(new_n765), .A3(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n780), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(KEYINPUT99), .A3(new_n739), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n777), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n758), .B1(new_n787), .B2(KEYINPUT29), .ZN(new_n788));
  INV_X1    g0588(.A(G330), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT30), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n570), .A2(new_n601), .A3(new_n651), .A4(new_n655), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n492), .A2(G179), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND4_X1   g0593(.A1(new_n560), .A2(new_n563), .A3(new_n651), .A4(new_n655), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n490), .A2(new_n355), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT30), .A4(new_n601), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT96), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n490), .A2(new_n797), .A3(new_n355), .A4(new_n703), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n703), .A2(new_n355), .ZN(new_n799));
  OAI21_X1  g0599(.A(KEYINPUT96), .B1(new_n492), .B2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n601), .A2(new_n485), .B1(new_n560), .B2(new_n563), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n798), .B(new_n800), .C1(new_n801), .C2(KEYINPUT97), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n801), .A2(KEYINPUT97), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n793), .B(new_n796), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AND3_X1   g0604(.A1(new_n804), .A2(KEYINPUT31), .A3(new_n734), .ZN(new_n805));
  AOI21_X1  g0605(.A(KEYINPUT31), .B1(new_n804), .B2(new_n734), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(KEYINPUT85), .B(new_n716), .C1(new_n512), .C2(new_n513), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n675), .B(new_n739), .C1(new_n808), .C2(new_n527), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n789), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n788), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n756), .B1(new_n811), .B2(G1), .ZN(G364));
  NOR2_X1   g0612(.A1(new_n741), .A2(new_n742), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(new_n789), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n263), .A2(G20), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G45), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G1), .ZN(new_n818));
  OR3_X1    g0618(.A1(new_n753), .A2(KEYINPUT100), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(KEYINPUT100), .B1(new_n753), .B2(new_n818), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n813), .A2(new_n789), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n815), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G13), .A2(G33), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(G20), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n813), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n821), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n215), .A2(new_n327), .ZN(new_n829));
  INV_X1    g0629(.A(G355), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n829), .A2(new_n830), .B1(G116), .B2(new_n215), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n752), .A2(new_n327), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n833), .B1(new_n231), .B2(new_n297), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n835), .A2(KEYINPUT101), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(KEYINPUT101), .B1(G45), .B2(new_n245), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n831), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n229), .B1(G20), .B2(new_n316), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n826), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n828), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(G179), .A2(G200), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT104), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n212), .A2(G190), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(G159), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT32), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n212), .A2(new_n633), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n355), .A2(G200), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n853), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n845), .A2(new_n851), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n859), .A2(KEYINPUT103), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(KEYINPUT103), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n858), .A2(G58), .B1(new_n863), .B2(G77), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n844), .A2(G190), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n865), .A2(new_n212), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(G97), .ZN(new_n868));
  NAND3_X1  g0668(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n869), .A2(G190), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n633), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n871), .A2(new_n202), .B1(new_n873), .B2(new_n207), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n576), .A2(G179), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n850), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(new_n659), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n845), .A2(new_n875), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n327), .B1(new_n878), .B2(new_n534), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n874), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n849), .A2(new_n864), .A3(new_n868), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n867), .A2(new_n587), .ZN(new_n882));
  INV_X1    g0682(.A(new_n846), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n858), .A2(G322), .B1(G329), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(G303), .ZN(new_n885));
  INV_X1    g0685(.A(G311), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n876), .A2(new_n885), .B1(new_n859), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n878), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n327), .B(new_n887), .C1(G283), .C2(new_n888), .ZN(new_n889));
  XNOR2_X1  g0689(.A(KEYINPUT33), .B(G317), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n890), .A2(new_n870), .B1(new_n872), .B2(G326), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n882), .A2(new_n884), .A3(new_n889), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n881), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n842), .B1(new_n839), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n827), .A2(new_n894), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n823), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(G396));
  AOI22_X1  g0697(.A1(new_n870), .A2(G150), .B1(new_n872), .B2(G137), .ZN(new_n898));
  INV_X1    g0698(.A(G143), .ZN(new_n899));
  OAI221_X1 g0699(.A(new_n898), .B1(new_n862), .B2(new_n847), .C1(new_n899), .C2(new_n857), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT34), .Z(new_n901));
  OAI21_X1  g0701(.A(new_n327), .B1(new_n878), .B2(new_n202), .ZN(new_n902));
  INV_X1    g0702(.A(new_n876), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n902), .B1(G50), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(G132), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n904), .B1(new_n905), .B2(new_n846), .C1(new_n866), .C2(new_n201), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n858), .A2(G294), .B1(new_n863), .B2(G116), .ZN(new_n907));
  INV_X1    g0707(.A(G283), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n436), .B1(new_n876), .B2(new_n534), .C1(new_n908), .C2(new_n871), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(G303), .B2(new_n872), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n907), .A2(new_n868), .A3(new_n910), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n846), .A2(new_n886), .B1(new_n659), .B2(new_n878), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(KEYINPUT105), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n901), .A2(new_n906), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n839), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n839), .A2(new_n824), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n821), .B1(new_n257), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n462), .A2(new_n734), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n454), .A2(new_n456), .ZN(new_n920));
  OAI22_X1  g0720(.A1(new_n457), .A2(new_n458), .B1(new_n920), .B2(new_n739), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n462), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n915), .B(new_n917), .C1(new_n924), .C2(new_n825), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n757), .B(new_n924), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n807), .A2(new_n809), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G330), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n828), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n926), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n925), .B1(new_n930), .B2(new_n931), .ZN(G384));
  NAND2_X1  g0732(.A1(new_n539), .A2(new_n540), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT35), .ZN(new_n934));
  OAI211_X1 g0734(.A(G116), .B(new_n230), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n935), .B1(new_n934), .B2(new_n933), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n231), .A2(G77), .A3(new_n391), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n207), .A2(G68), .ZN(new_n939));
  AOI211_X1 g0739(.A(new_n211), .B(G13), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n732), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n682), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n918), .B1(new_n757), .B2(new_n924), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n281), .A2(new_n739), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n314), .A2(new_n319), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n280), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n948), .B2(new_n323), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n320), .A2(new_n324), .A3(new_n945), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n401), .A2(new_n254), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n398), .B(G68), .C1(new_n397), .C2(new_n388), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT16), .B1(new_n954), .B2(new_n393), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n428), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n942), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n412), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n957), .A2(new_n958), .A3(new_n429), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT37), .ZN(new_n960));
  AOI221_X4 g0760(.A(KEYINPUT106), .B1(new_n410), .B2(new_n411), .C1(new_n425), .C2(new_n428), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT106), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n432), .B2(new_n412), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n432), .A2(new_n942), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT37), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n965), .A2(new_n966), .A3(new_n429), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n960), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n957), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n435), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT38), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n968), .A2(new_n970), .A3(KEYINPUT38), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n943), .B1(new_n952), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n948), .A2(new_n734), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n973), .A2(KEYINPUT39), .A3(new_n974), .ZN(new_n978));
  AND3_X1   g0778(.A1(new_n968), .A2(new_n970), .A3(KEYINPUT38), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n965), .B(new_n429), .C1(new_n402), .C2(new_n413), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT37), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n964), .B2(new_n967), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n685), .B1(new_n680), .B2(new_n681), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(new_n965), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n979), .B1(new_n984), .B2(new_n972), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n977), .B(new_n978), .C1(new_n985), .C2(KEYINPUT39), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n695), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(new_n788), .B2(new_n464), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n988), .B(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n325), .A2(new_n946), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n945), .B1(new_n320), .B2(new_n324), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n923), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n927), .A2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(KEYINPUT40), .B1(new_n995), .B2(new_n985), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT40), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n975), .A2(new_n927), .A3(new_n997), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n464), .A2(new_n927), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n789), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n1000), .B2(new_n999), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n991), .A2(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n211), .B2(new_n816), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n991), .A2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n941), .B1(new_n1004), .B2(new_n1005), .ZN(G367));
  INV_X1    g0806(.A(KEYINPUT108), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n549), .A2(new_n734), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n702), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n696), .A2(new_n734), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1009), .A2(KEYINPUT107), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(KEYINPUT107), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n715), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n734), .B1(new_n1013), .B2(new_n572), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n702), .A2(new_n1008), .B1(new_n696), .B2(new_n734), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1015), .A2(new_n744), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT42), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1007), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1018), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT107), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1015), .A2(KEYINPUT107), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n696), .B1(new_n1025), .B2(new_n715), .ZN(new_n1026));
  OAI211_X1 g0826(.A(KEYINPUT108), .B(new_n1020), .C1(new_n1026), .C2(new_n734), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1019), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n743), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n1025), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n672), .A2(new_n739), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n719), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n724), .B2(new_n1032), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n1029), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1031), .B1(new_n1029), .B2(new_n1035), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(KEYINPUT43), .B2(new_n1034), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n1031), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1034), .A2(KEYINPUT43), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1029), .A2(new_n1031), .A3(new_n1035), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n818), .B(KEYINPUT109), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(KEYINPUT99), .B1(new_n785), .B2(new_n739), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n776), .B(new_n734), .C1(new_n780), .C2(new_n784), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT29), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n758), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n928), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n746), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(new_n1015), .A3(new_n747), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT44), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1021), .B1(new_n748), .B2(new_n746), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT45), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1021), .B(KEYINPUT45), .C1(new_n748), .C2(new_n746), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1056), .A2(new_n1061), .A3(new_n743), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n743), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n716), .A2(new_n739), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n744), .B1(new_n738), .B2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n814), .B(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1052), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n753), .B(KEYINPUT41), .Z(new_n1070));
  OAI21_X1  g0870(.A(new_n1046), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1038), .A2(new_n1044), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n867), .A2(G68), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n863), .A2(G50), .B1(G137), .B2(new_n883), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n858), .A2(G150), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n871), .A2(new_n847), .B1(new_n873), .B2(new_n899), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n876), .A2(new_n201), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n878), .A2(new_n257), .ZN(new_n1078));
  NOR4_X1   g0878(.A1(new_n1076), .A2(new_n436), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(KEYINPUT46), .B1(new_n903), .B2(G116), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n903), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n873), .B2(new_n886), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n1081), .B(new_n1083), .C1(new_n587), .C2(new_n870), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n858), .A2(G303), .B1(new_n863), .B2(G283), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1084), .B(new_n1085), .C1(new_n534), .C2(new_n866), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n436), .B1(new_n878), .B2(new_n497), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT110), .B(G317), .Z(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n883), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT111), .Z(new_n1090));
  OAI21_X1  g0890(.A(new_n1080), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT47), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n839), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n832), .A2(new_n241), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n452), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n841), .B1(new_n752), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n821), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n826), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1093), .B(new_n1097), .C1(new_n1098), .C2(new_n1034), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1072), .A2(new_n1099), .ZN(G387));
  INV_X1    g0900(.A(KEYINPUT114), .ZN(new_n1101));
  OR3_X1    g0901(.A1(new_n811), .A2(new_n1068), .A3(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n811), .A2(new_n1068), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1101), .B1(new_n811), .B2(new_n1068), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1102), .A2(new_n753), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n736), .A2(new_n737), .A3(new_n826), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n751), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n1107), .A2(new_n829), .B1(G107), .B2(new_n215), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n751), .A2(KEYINPUT112), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n751), .A2(KEYINPUT112), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n449), .A2(new_n207), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(KEYINPUT50), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n297), .B1(new_n202), .B2(new_n257), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1111), .B2(KEYINPUT50), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n833), .B1(new_n238), .B2(G45), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1108), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n828), .B1(new_n1117), .B2(new_n841), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n876), .A2(new_n257), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n883), .B2(G150), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT113), .Z(new_n1121));
  NAND2_X1  g0921(.A1(new_n867), .A2(new_n1095), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n327), .B1(new_n878), .B2(new_n497), .C1(new_n202), .C2(new_n859), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G159), .B2(new_n872), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n858), .A2(G50), .B1(new_n378), .B2(new_n870), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1122), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n883), .A2(G326), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n327), .B1(new_n888), .B2(G116), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n903), .A2(new_n587), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n866), .B2(new_n908), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n858), .A2(new_n1088), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n870), .A2(G311), .B1(new_n872), .B2(G322), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n885), .C2(new_n862), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT48), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1134), .B2(new_n1133), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT49), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1127), .B(new_n1128), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1126), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1118), .B1(new_n1140), .B2(new_n839), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1068), .A2(new_n1045), .B1(new_n1106), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1105), .A2(new_n1142), .ZN(G393));
  OAI221_X1 g0943(.A(new_n840), .B1(new_n497), .B2(new_n215), .C1(new_n833), .C2(new_n248), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT117), .B1(new_n828), .B2(new_n1144), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n828), .A2(KEYINPUT117), .A3(new_n1144), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n858), .A2(G311), .B1(G317), .B2(new_n872), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT52), .Z(new_n1148));
  OAI221_X1 g0948(.A(new_n436), .B1(new_n878), .B2(new_n534), .C1(new_n908), .C2(new_n876), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G322), .B2(new_n883), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT119), .Z(new_n1151));
  INV_X1    g0951(.A(G294), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n871), .A2(new_n885), .B1(new_n859), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n867), .B2(G116), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1148), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G150), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n857), .A2(new_n847), .B1(new_n1156), .B2(new_n873), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT51), .Z(new_n1158));
  AOI22_X1  g0958(.A1(new_n863), .A2(new_n449), .B1(G50), .B2(new_n870), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT118), .ZN(new_n1160));
  OR2_X1    g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n436), .B1(new_n888), .B2(G87), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n202), .B2(new_n876), .C1(new_n846), .C2(new_n899), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G77), .B2(new_n867), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1155), .B1(new_n1158), .B2(new_n1166), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1145), .B(new_n1146), .C1(new_n1167), .C2(new_n839), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n1025), .B2(new_n1098), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1064), .A2(new_n811), .A3(new_n1068), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(new_n753), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1063), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1056), .A2(new_n1061), .A3(new_n743), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1173), .A2(KEYINPUT115), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT115), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1062), .B1(new_n1063), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1103), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1170), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT116), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1175), .A2(new_n1177), .A3(KEYINPUT116), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1182), .A2(new_n1183), .A3(new_n1045), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1179), .A2(new_n1184), .ZN(G390));
  NAND3_X1  g0985(.A1(new_n1049), .A2(new_n464), .A3(new_n1050), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n464), .A2(new_n810), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n695), .A3(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n944), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n951), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n810), .B2(new_n924), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n927), .A2(G330), .A3(new_n994), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n777), .A2(new_n786), .A3(new_n919), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n922), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1188), .B1(new_n1193), .B2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n922), .A3(new_n1190), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n985), .A2(new_n977), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n978), .B1(new_n985), .B2(KEYINPUT39), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n944), .A2(new_n951), .B1(new_n948), .B2(new_n734), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n810), .A2(KEYINPUT120), .A3(new_n994), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1206), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1201), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1198), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n1211), .A2(new_n919), .B1(new_n462), .B2(new_n921), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n789), .B(new_n923), .C1(new_n807), .C2(new_n809), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n924), .B1(new_n949), .B2(new_n950), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n1213), .A2(new_n1190), .B1(new_n928), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1193), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1216), .A2(new_n990), .A3(new_n1187), .ZN(new_n1217));
  AOI221_X4 g1017(.A(new_n1206), .B1(new_n1202), .B2(new_n1203), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1208), .B1(new_n1201), .B2(new_n1204), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1210), .A2(new_n1220), .A3(new_n753), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1202), .A2(new_n824), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n916), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n828), .B1(new_n378), .B2(new_n1224), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n866), .A2(new_n257), .B1(new_n857), .B2(new_n494), .ZN(new_n1226));
  XOR2_X1   g1026(.A(new_n1226), .B(KEYINPUT121), .Z(new_n1227));
  AOI22_X1  g1027(.A1(new_n863), .A2(G97), .B1(G294), .B2(new_n883), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n327), .B(new_n877), .C1(G68), .C2(new_n888), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n870), .A2(G107), .B1(new_n872), .B2(G283), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n903), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT53), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n876), .B2(new_n1156), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n883), .A2(G125), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(KEYINPUT54), .B(G143), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1235), .B1(new_n905), .B2(new_n857), .C1(new_n862), .C2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n327), .B1(new_n878), .B2(new_n207), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G137), .B2(new_n870), .ZN(new_n1239));
  INV_X1    g1039(.A(G128), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1239), .B1(new_n1240), .B2(new_n873), .C1(new_n866), .C2(new_n847), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n1227), .A2(new_n1231), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1225), .B1(new_n1242), .B2(new_n839), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1222), .A2(new_n1045), .B1(new_n1223), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1221), .A2(new_n1244), .ZN(G378));
  NOR2_X1   g1045(.A1(new_n365), .A2(new_n732), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n377), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1246), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n693), .A2(new_n361), .A3(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1250));
  AND3_X1   g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n999), .B2(G330), .ZN(new_n1255));
  AOI211_X1 g1055(.A(new_n789), .B(new_n1253), .C1(new_n996), .C2(new_n998), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n987), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1214), .B1(new_n809), .B2(new_n807), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n984), .A2(new_n972), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(new_n974), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n997), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n998), .ZN(new_n1262));
  OAI21_X1  g1062(.A(G330), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n1253), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n999), .A2(G330), .A3(new_n1254), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n988), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1046), .B1(new_n1257), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1253), .A2(new_n824), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n828), .B1(G50), .B2(new_n1224), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(G33), .A2(G41), .ZN(new_n1270));
  AOI211_X1 g1070(.A(G50), .B(new_n1270), .C1(new_n436), .C2(new_n296), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n858), .A2(G107), .B1(G283), .B2(new_n883), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n452), .A2(new_n859), .B1(new_n878), .B2(new_n201), .ZN(new_n1273));
  NOR4_X1   g1073(.A1(new_n1273), .A2(new_n1119), .A3(G41), .A4(new_n327), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n870), .A2(G97), .B1(new_n872), .B2(G116), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1073), .A2(new_n1272), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT58), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1271), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n871), .A2(new_n905), .ZN(new_n1279));
  INV_X1    g1079(.A(G137), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n876), .A2(new_n1236), .B1(new_n859), .B2(new_n1280), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1279), .B(new_n1281), .C1(G125), .C2(new_n872), .ZN(new_n1282));
  OAI221_X1 g1082(.A(new_n1282), .B1(new_n1240), .B2(new_n857), .C1(new_n1156), .C2(new_n866), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT59), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1270), .B1(new_n878), .B2(new_n847), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n883), .B2(G124), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1283), .A2(KEYINPUT59), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n1278), .B1(new_n1277), .B2(new_n1276), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1269), .B1(new_n1289), .B2(new_n839), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1268), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1267), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1257), .A2(new_n1266), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1295));
  OAI211_X1 g1095(.A(KEYINPUT57), .B(new_n1294), .C1(new_n1295), .C2(new_n1188), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n753), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1188), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1210), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(KEYINPUT57), .B1(new_n1299), .B2(new_n1294), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1293), .B1(new_n1297), .B2(new_n1300), .ZN(G375));
  INV_X1    g1101(.A(new_n1070), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1188), .A2(new_n1193), .A3(new_n1197), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1217), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n951), .A2(new_n824), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n828), .B1(G68), .B2(new_n1224), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n867), .A2(G50), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n858), .A2(G137), .B1(G128), .B2(new_n883), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n876), .A2(new_n847), .B1(new_n859), .B2(new_n1156), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n436), .B(new_n1309), .C1(G58), .C2(new_n888), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1236), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1311), .A2(new_n870), .B1(G132), .B2(new_n872), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1307), .A2(new_n1308), .A3(new_n1310), .A4(new_n1312), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n858), .A2(G283), .B1(new_n863), .B2(G107), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(new_n885), .B2(new_n846), .ZN(new_n1315));
  AOI211_X1 g1115(.A(new_n327), .B(new_n1078), .C1(G97), .C2(new_n903), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n870), .A2(G116), .B1(new_n872), .B2(G294), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1122), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1313), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1306), .B1(new_n1319), .B2(new_n839), .ZN(new_n1320));
  AOI22_X1  g1120(.A1(new_n1216), .A2(new_n1045), .B1(new_n1305), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1304), .A2(new_n1321), .ZN(G381));
  NOR2_X1   g1122(.A1(G375), .A2(G378), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1072), .A2(new_n1179), .A3(new_n1099), .A4(new_n1184), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1105), .A2(new_n896), .A3(new_n1142), .ZN(new_n1326));
  NOR3_X1   g1126(.A1(new_n1326), .A2(G381), .A3(G384), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1327), .ZN(G407));
  NAND2_X1  g1128(.A1(new_n733), .A2(G213), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1323), .A2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(G407), .A2(G213), .A3(new_n1331), .ZN(new_n1332));
  XOR2_X1   g1132(.A(new_n1332), .B(KEYINPUT122), .Z(G409));
  INV_X1    g1133(.A(KEYINPUT126), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G393), .A2(G396), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1335), .A2(new_n1326), .ZN(new_n1336));
  AOI22_X1  g1136(.A1(new_n1072), .A2(new_n1099), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1336), .B1(new_n1325), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(G387), .A2(G390), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1335), .A2(new_n1326), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1339), .A2(new_n1340), .A3(new_n1324), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1338), .A2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G375), .A2(G378), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1302), .B(new_n1294), .C1(new_n1295), .C2(new_n1188), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1345), .A2(new_n1221), .A3(new_n1244), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT123), .ZN(new_n1347));
  NOR3_X1   g1147(.A1(new_n1255), .A2(new_n1256), .A3(new_n987), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n988), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1045), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  AOI21_X1  g1150(.A(new_n1347), .B1(new_n1350), .B2(new_n1291), .ZN(new_n1351));
  NOR3_X1   g1151(.A1(new_n1267), .A2(KEYINPUT123), .A3(new_n1292), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1330), .B1(new_n1346), .B2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1217), .A2(KEYINPUT60), .ZN(new_n1355));
  AND2_X1   g1155(.A1(new_n1355), .A2(new_n1303), .ZN(new_n1356));
  NAND4_X1  g1156(.A1(new_n1188), .A2(new_n1197), .A3(KEYINPUT60), .A4(new_n1193), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n753), .ZN(new_n1358));
  OAI211_X1 g1158(.A(G384), .B(new_n1321), .C1(new_n1356), .C2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(G384), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1358), .B1(new_n1303), .B2(new_n1355), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1321), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1360), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  AND2_X1   g1163(.A1(new_n1359), .A2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1344), .A2(new_n1354), .A3(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT125), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT62), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1365), .A2(new_n1366), .A3(new_n1367), .ZN(new_n1368));
  INV_X1    g1168(.A(G378), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1352), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1350), .A2(new_n1291), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(KEYINPUT123), .ZN(new_n1372));
  NAND4_X1  g1172(.A1(new_n1369), .A2(new_n1370), .A3(new_n1372), .A4(new_n1345), .ZN(new_n1373));
  INV_X1    g1173(.A(new_n753), .ZN(new_n1374));
  AOI22_X1  g1174(.A1(new_n1210), .A2(new_n1298), .B1(new_n1266), .B2(new_n1257), .ZN(new_n1375));
  AOI21_X1  g1175(.A(new_n1374), .B1(new_n1375), .B2(KEYINPUT57), .ZN(new_n1376));
  NAND2_X1  g1176(.A1(new_n1299), .A2(new_n1294), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT57), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1377), .A2(new_n1378), .ZN(new_n1379));
  AOI21_X1  g1179(.A(new_n1371), .B1(new_n1376), .B2(new_n1379), .ZN(new_n1380));
  OAI211_X1 g1180(.A(new_n1373), .B(new_n1329), .C1(new_n1380), .C2(new_n1369), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1330), .A2(G2897), .ZN(new_n1382));
  AND3_X1   g1182(.A1(new_n1359), .A2(new_n1363), .A3(new_n1382), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1382), .B1(new_n1359), .B2(new_n1363), .ZN(new_n1384));
  NOR2_X1   g1184(.A1(new_n1383), .A2(new_n1384), .ZN(new_n1385));
  AOI21_X1  g1185(.A(KEYINPUT61), .B1(new_n1381), .B2(new_n1385), .ZN(new_n1386));
  AND2_X1   g1186(.A1(new_n1368), .A2(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1365), .A2(new_n1367), .ZN(new_n1388));
  NAND4_X1  g1188(.A1(new_n1344), .A2(new_n1354), .A3(new_n1364), .A4(KEYINPUT62), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1388), .A2(KEYINPUT125), .A3(new_n1389), .ZN(new_n1390));
  AOI21_X1  g1190(.A(new_n1343), .B1(new_n1387), .B2(new_n1390), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT61), .ZN(new_n1392));
  NAND3_X1  g1192(.A1(new_n1338), .A2(new_n1392), .A3(new_n1341), .ZN(new_n1393));
  INV_X1    g1193(.A(KEYINPUT124), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1381), .A2(new_n1385), .ZN(new_n1396));
  NAND4_X1  g1196(.A1(new_n1338), .A2(KEYINPUT124), .A3(new_n1392), .A4(new_n1341), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1395), .A2(new_n1396), .A3(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1365), .A2(KEYINPUT63), .ZN(new_n1399));
  OR2_X1    g1199(.A1(new_n1365), .A2(KEYINPUT63), .ZN(new_n1400));
  AOI21_X1  g1200(.A(new_n1398), .B1(new_n1399), .B2(new_n1400), .ZN(new_n1401));
  OAI21_X1  g1201(.A(new_n1334), .B1(new_n1391), .B2(new_n1401), .ZN(new_n1402));
  AND3_X1   g1202(.A1(new_n1388), .A2(KEYINPUT125), .A3(new_n1389), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1368), .A2(new_n1386), .ZN(new_n1404));
  OAI21_X1  g1204(.A(new_n1342), .B1(new_n1403), .B2(new_n1404), .ZN(new_n1405));
  NAND2_X1  g1205(.A1(new_n1400), .A2(new_n1399), .ZN(new_n1406));
  AND2_X1   g1206(.A1(new_n1395), .A2(new_n1396), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1406), .A2(new_n1407), .A3(new_n1397), .ZN(new_n1408));
  NAND3_X1  g1208(.A1(new_n1405), .A2(KEYINPUT126), .A3(new_n1408), .ZN(new_n1409));
  NAND2_X1  g1209(.A1(new_n1402), .A2(new_n1409), .ZN(G405));
  XNOR2_X1  g1210(.A(G375), .B(new_n1369), .ZN(new_n1411));
  XNOR2_X1  g1211(.A(new_n1411), .B(new_n1364), .ZN(new_n1412));
  OAI21_X1  g1212(.A(KEYINPUT127), .B1(new_n1412), .B2(new_n1343), .ZN(new_n1413));
  NAND2_X1  g1213(.A1(new_n1412), .A2(new_n1343), .ZN(new_n1414));
  NAND2_X1  g1214(.A1(new_n1413), .A2(new_n1414), .ZN(new_n1415));
  NOR3_X1   g1215(.A1(new_n1412), .A2(KEYINPUT127), .A3(new_n1343), .ZN(new_n1416));
  NOR2_X1   g1216(.A1(new_n1415), .A2(new_n1416), .ZN(G402));
endmodule


