//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  AND2_X1   g034(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n464), .B1(new_n469), .B2(KEYINPUT70), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n466), .A2(new_n468), .A3(new_n471), .A4(G125), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n462), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n465), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n462), .A2(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT71), .B1(new_n465), .B2(KEYINPUT3), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n478), .A2(new_n467), .A3(G2104), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(new_n479), .A3(new_n466), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n475), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n473), .A2(new_n481), .ZN(G160));
  NOR2_X1   g057(.A1(new_n480), .A2(new_n462), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OAI221_X1 g059(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  AND3_X1   g061(.A1(new_n477), .A2(new_n479), .A3(new_n466), .ZN(new_n487));
  INV_X1    g062(.A(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(new_n488), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n494), .A2(G138), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n466), .A2(new_n468), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n492), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT4), .A2(G138), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n462), .A2(new_n504), .B1(G126), .B2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n498), .B(new_n502), .C1(new_n505), .C2(new_n480), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT72), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n510), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n520), .A2(G88), .A3(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n524), .A2(KEYINPUT73), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT73), .B1(new_n524), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n513), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G166));
  NAND3_X1  g106(.A1(new_n510), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(G51), .B2(new_n526), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n520), .A2(G89), .A3(new_n523), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n516), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n542), .A2(G651), .B1(new_n526), .B2(G52), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT74), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n520), .A2(G90), .A3(new_n523), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n547), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(G68), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n516), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n553), .A2(G651), .B1(new_n526), .B2(G43), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n520), .A2(G81), .A3(new_n523), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT75), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n554), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(new_n521), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI22_X1  g144(.A1(new_n568), .A2(new_n569), .B1(KEYINPUT77), .B2(KEYINPUT9), .ZN(new_n570));
  XNOR2_X1  g145(.A(KEYINPUT77), .B(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n526), .A2(G53), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n510), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n512), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n520), .A2(G91), .A3(new_n523), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(G299));
  NAND2_X1  g152(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  OAI211_X1 g154(.A(new_n579), .B(new_n513), .C1(new_n528), .C2(new_n529), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G303));
  NAND3_X1  g156(.A1(new_n521), .A2(G49), .A3(G543), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n521), .A2(KEYINPUT79), .A3(G49), .A4(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n520), .A2(G87), .A3(new_n523), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n508), .B2(new_n509), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n592), .B2(KEYINPUT80), .ZN(new_n593));
  OAI211_X1 g168(.A(KEYINPUT80), .B(G61), .C1(new_n514), .C2(new_n515), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n520), .A2(G86), .A3(new_n523), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n526), .A2(G48), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n516), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n526), .B2(G47), .ZN(new_n603));
  XNOR2_X1  g178(.A(KEYINPUT81), .B(G85), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n520), .A2(new_n523), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(G290));
  NAND3_X1  g181(.A1(new_n520), .A2(G92), .A3(new_n523), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g184(.A1(new_n520), .A2(KEYINPUT10), .A3(G92), .A4(new_n523), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(G79), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n516), .B2(new_n613), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n614), .A2(G651), .B1(new_n526), .B2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  MUX2_X1   g191(.A(new_n616), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g192(.A(new_n616), .B(G301), .S(G868), .Z(G321));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G299), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G168), .B2(new_n619), .ZN(G280));
  XNOR2_X1  g196(.A(G280), .B(KEYINPUT82), .ZN(G297));
  INV_X1    g197(.A(new_n616), .ZN(new_n623));
  INV_X1    g198(.A(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n624), .B2(G860), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(G148));
  NAND2_X1  g201(.A1(new_n560), .A2(new_n619), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n616), .A2(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n619), .ZN(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g205(.A1(new_n488), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n483), .A2(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n489), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2096), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(G156));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n643), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n659), .A2(KEYINPUT85), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n655), .A2(new_n661), .A3(new_n657), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT17), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT87), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n666), .A2(new_n667), .ZN(new_n673));
  INV_X1    g248(.A(new_n665), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n669), .B1(new_n674), .B2(new_n668), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n669), .A2(new_n665), .A3(new_n667), .ZN(new_n677));
  XOR2_X1   g252(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n672), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(new_n634), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT88), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n684), .B(new_n685), .Z(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1981), .ZN(new_n699));
  INV_X1    g274(.A(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT89), .B(KEYINPUT90), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n701), .A2(new_n703), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n687), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n706), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n708), .A2(new_n686), .A3(new_n704), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(G229));
  INV_X1    g286(.A(G16), .ZN(new_n712));
  NOR2_X1   g287(.A1(G286), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(KEYINPUT97), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT97), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G16), .B2(G21), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1966), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n721), .B2(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G160), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT94), .B(G2067), .Z(new_n725));
  XOR2_X1   g300(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n720), .A2(G26), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n483), .A2(G128), .ZN(new_n729));
  OAI221_X1 g304(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n730));
  INV_X1    g305(.A(G140), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n489), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n728), .B1(new_n733), .B2(new_n720), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n719), .B1(G2084), .B2(new_n724), .C1(new_n725), .C2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n474), .A2(G105), .ZN(new_n736));
  INV_X1    g311(.A(G141), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n489), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT96), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  AOI211_X1 g316(.A(new_n738), .B(new_n741), .C1(G129), .C2(new_n483), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n720), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n720), .B2(G32), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n712), .A2(G20), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT23), .ZN(new_n748));
  INV_X1    g323(.A(G299), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(new_n712), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n746), .B1(G1956), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n734), .A2(new_n725), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n744), .B2(new_n745), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n720), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n720), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2090), .ZN(new_n757));
  NOR4_X1   g332(.A1(new_n735), .A2(new_n751), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT31), .B(G11), .Z(new_n759));
  INV_X1    g334(.A(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(KEYINPUT30), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(KEYINPUT30), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n639), .B2(new_n720), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n720), .A2(G33), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT25), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n494), .A2(new_n495), .ZN(new_n767));
  NAND2_X1  g342(.A1(G103), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n766), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n462), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n770));
  NAND2_X1  g345(.A1(G115), .A2(G2104), .ZN(new_n771));
  INV_X1    g346(.A(G127), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n497), .B2(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n769), .A2(new_n770), .B1(new_n773), .B2(new_n767), .ZN(new_n774));
  INV_X1    g349(.A(G139), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n489), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n765), .B1(new_n776), .B2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G164), .A2(new_n720), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G27), .B2(new_n720), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT98), .B(G2078), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n779), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g358(.A(new_n764), .B(new_n783), .C1(new_n781), .C2(new_n782), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n750), .A2(G1956), .B1(G2084), .B2(new_n724), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n777), .A2(new_n778), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n712), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n712), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(G1961), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n712), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n623), .B2(new_n712), .ZN(new_n793));
  INV_X1    g368(.A(G1348), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G1961), .B2(new_n789), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n791), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n712), .A2(G19), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(new_n561), .B2(new_n712), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT92), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(G1341), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n758), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(G166), .A2(G16), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G16), .B2(G22), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT32), .B(G1981), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n712), .A2(G23), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n712), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT33), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1976), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n804), .A2(new_n805), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n810), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(KEYINPUT34), .ZN(new_n819));
  NOR2_X1   g394(.A1(G25), .A2(G29), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n487), .A2(G131), .A3(new_n488), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT91), .Z(new_n822));
  OAI21_X1  g397(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n823));
  INV_X1    g398(.A(G107), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n767), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n483), .B2(G119), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n820), .B1(new_n827), .B2(G29), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT35), .B(G1991), .Z(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n712), .A2(G24), .ZN(new_n833));
  INV_X1    g408(.A(G290), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n712), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G1986), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n831), .A2(new_n832), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n818), .A2(new_n819), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT36), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n818), .A2(new_n840), .A3(new_n819), .A4(new_n837), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n802), .B1(new_n839), .B2(new_n841), .ZN(G311));
  INV_X1    g417(.A(G311), .ZN(G150));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n516), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT99), .B(G55), .Z(new_n847));
  AOI22_X1  g422(.A1(new_n846), .A2(G651), .B1(new_n526), .B2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT100), .B(G93), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n520), .A2(new_n523), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n560), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n556), .A2(new_n851), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT38), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n624), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(KEYINPUT39), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n859), .A2(new_n860), .A3(G860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n851), .A2(G860), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n861), .A2(new_n863), .ZN(G145));
  NAND2_X1  g439(.A1(new_n483), .A2(G130), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT101), .Z(new_n866));
  INV_X1    g441(.A(G142), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n462), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI221_X1 g444(.A(new_n866), .B1(new_n867), .B2(new_n489), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n732), .B(new_n506), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n827), .B(KEYINPUT102), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n632), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n742), .B(new_n776), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n822), .A2(new_n826), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT102), .ZN(new_n879));
  INV_X1    g454(.A(new_n632), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n875), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n877), .B1(new_n875), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n873), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n875), .A2(new_n881), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n876), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n875), .A2(new_n877), .A3(new_n881), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n886), .A2(new_n872), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n639), .B(G160), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G162), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  INV_X1    g468(.A(new_n891), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n884), .A2(new_n888), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n851), .A2(new_n619), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  XNOR2_X1  g474(.A(G305), .B(G288), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n530), .A2(new_n834), .ZN(new_n901));
  OAI211_X1 g476(.A(new_n513), .B(G290), .C1(new_n528), .C2(new_n529), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n900), .B1(new_n902), .B2(new_n901), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT104), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n904), .B2(new_n905), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n902), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n812), .B(G305), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT104), .A3(new_n903), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n906), .B1(new_n914), .B2(new_n899), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n616), .A2(new_n749), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n611), .A2(G299), .A3(new_n615), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(KEYINPUT41), .A3(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n916), .A2(KEYINPUT103), .A3(KEYINPUT41), .A4(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n916), .A2(new_n917), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n920), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n855), .B(new_n628), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n927), .B2(new_n922), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n915), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n898), .B1(new_n930), .B2(new_n619), .ZN(G295));
  OAI21_X1  g506(.A(new_n898), .B1(new_n930), .B2(new_n619), .ZN(G331));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  OAI21_X1  g508(.A(G168), .B1(new_n547), .B2(new_n548), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n543), .A2(new_n545), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT74), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n936), .A2(G286), .A3(new_n546), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n852), .A2(new_n934), .A3(new_n937), .A4(new_n854), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n936), .A2(G286), .A3(new_n546), .ZN(new_n939));
  AOI21_X1  g514(.A(G286), .B1(new_n936), .B2(new_n546), .ZN(new_n940));
  INV_X1    g515(.A(new_n851), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n941), .B1(new_n557), .B2(new_n559), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n939), .A2(new_n940), .B1(new_n942), .B2(new_n853), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(new_n943), .A3(new_n922), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n943), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n945), .B1(new_n925), .B2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(G37), .B1(new_n914), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n918), .A2(KEYINPUT105), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT105), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n916), .A2(new_n951), .A3(KEYINPUT41), .A4(new_n917), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n924), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n946), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n955), .A3(new_n946), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n913), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n948), .B(KEYINPUT107), .C1(new_n954), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n925), .A2(new_n946), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(new_n912), .A3(new_n908), .A4(new_n944), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n893), .B(new_n960), .C1(new_n957), .C2(new_n954), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n933), .B1(new_n958), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n959), .A2(new_n944), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n913), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT43), .B1(new_n948), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n948), .A2(new_n966), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT43), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n970), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(G397));
  XOR2_X1   g549(.A(new_n732), .B(G2067), .Z(new_n975));
  XNOR2_X1  g550(.A(new_n742), .B(G1996), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n878), .A2(new_n830), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n827), .A2(new_n829), .ZN(new_n978));
  AND4_X1   g553(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(G290), .B(new_n700), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(G40), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n473), .A2(new_n982), .A3(new_n481), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n506), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT108), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n506), .A2(new_n984), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(new_n983), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n586), .A2(new_n587), .A3(G1976), .A4(new_n588), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n992), .A2(KEYINPUT110), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(KEYINPUT110), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT52), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT52), .B1(G288), .B2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n597), .A2(new_n598), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(KEYINPUT111), .A3(new_n1002), .A4(new_n596), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n596), .A2(new_n1002), .A3(new_n597), .A4(new_n598), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(G305), .A2(G1981), .ZN(new_n1008));
  AND3_X1   g583(.A1(new_n1007), .A2(KEYINPUT49), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT49), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1000), .B1(new_n1011), .B2(new_n991), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n578), .A2(G8), .A3(new_n580), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n578), .A2(KEYINPUT55), .A3(G8), .A4(new_n580), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n506), .A2(new_n984), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1021), .A3(new_n983), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n805), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1024), .B1(new_n506), .B2(new_n984), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n469), .A2(KEYINPUT70), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(new_n472), .A3(new_n463), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n767), .ZN(new_n1028));
  INV_X1    g603(.A(new_n481), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(G40), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n506), .A2(new_n1024), .A3(new_n984), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT109), .B(G2090), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n989), .B1(new_n1023), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1012), .A2(new_n1017), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n997), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1037), .B(KEYINPUT112), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1007), .B1(new_n1011), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n991), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1017), .A2(new_n1035), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1044), .A2(KEYINPUT113), .A3(new_n983), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT113), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1025), .B2(new_n1030), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1045), .A2(new_n1047), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1023), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1012), .A2(new_n1043), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G286), .A2(new_n989), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1022), .A2(KEYINPUT114), .A3(new_n718), .ZN(new_n1054));
  INV_X1    g629(.A(G2084), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1031), .A2(new_n1055), .A3(new_n1032), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT114), .B1(new_n1022), .B2(new_n718), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1053), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1042), .B1(new_n1052), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1017), .A2(new_n1035), .ZN(new_n1061));
  OAI211_X1 g636(.A(KEYINPUT63), .B(new_n1053), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1061), .A2(new_n1043), .A3(new_n1012), .A4(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1041), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2078), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1020), .A2(new_n1066), .A3(new_n1021), .A4(new_n983), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1068));
  NAND3_X1  g643(.A1(new_n1044), .A2(new_n983), .A3(new_n1032), .ZN(new_n1069));
  INV_X1    g644(.A(G1961), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1067), .A2(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT122), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1073), .A2(new_n985), .A3(new_n1030), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1072), .B1(new_n1074), .B2(new_n1066), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT53), .B1(new_n1067), .B2(KEYINPUT122), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT124), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1080), .A3(G171), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1074), .A2(new_n1082), .A3(KEYINPUT53), .A4(new_n1066), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT125), .B1(new_n1067), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(G301), .A3(new_n1071), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT126), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT126), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n1089), .A3(G301), .A4(new_n1071), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1079), .A2(new_n1081), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1086), .B2(new_n1071), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1067), .A2(KEYINPUT122), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n985), .A2(new_n1030), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1096), .A2(new_n1072), .A3(new_n1066), .A4(new_n1021), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1097), .A3(KEYINPUT53), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1098), .A2(G301), .A3(new_n1071), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1094), .A2(new_n1099), .A3(new_n1092), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(new_n1052), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1074), .B2(G1966), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1103), .A2(G168), .A3(new_n1056), .A4(new_n1054), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(G8), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G286), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1108), .A2(new_n1104), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1093), .A2(new_n1101), .A3(new_n1111), .A4(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1045), .A2(new_n1047), .A3(new_n1032), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT115), .B(G1956), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1074), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n573), .B(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1120), .A2(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n575), .A2(new_n576), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT117), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1121), .A2(new_n1123), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT118), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1118), .A2(KEYINPUT118), .A3(new_n1124), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1069), .A2(new_n794), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1030), .A2(new_n1018), .A3(G2067), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n616), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT119), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1074), .A2(new_n1117), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1124), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1126), .A2(new_n1127), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1127), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(new_n1125), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1135), .A2(new_n1136), .A3(KEYINPUT120), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1139), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1139), .B1(new_n1118), .B2(new_n1124), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n1137), .ZN(new_n1148));
  AOI21_X1  g723(.A(G1348), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1149), .A2(new_n623), .A3(new_n1129), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT60), .B1(new_n1150), .B2(new_n1131), .ZN(new_n1151));
  OR4_X1    g726(.A1(KEYINPUT60), .A2(new_n1149), .A3(new_n616), .A4(new_n1129), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1030), .A2(new_n1018), .ZN(new_n1153));
  XNOR2_X1  g728(.A(KEYINPUT58), .B(G1341), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1022), .A2(G1996), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n561), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1156), .A2(KEYINPUT59), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1151), .B(new_n1152), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1148), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1138), .B1(new_n1146), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1065), .B1(new_n1114), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  AND3_X1   g738(.A1(new_n1107), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1112), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1111), .A2(KEYINPUT62), .A3(new_n1113), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1052), .B1(new_n1081), .B2(new_n1079), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n988), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(G290), .A2(G1986), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n987), .A2(KEYINPUT48), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n987), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1172), .B1(new_n979), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT48), .B1(new_n987), .B2(new_n1171), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(G1996), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n987), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g753(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(KEYINPUT46), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n975), .A2(new_n742), .ZN(new_n1181));
  OAI22_X1  g756(.A1(new_n1179), .A2(new_n1180), .B1(new_n1173), .B2(new_n1181), .ZN(new_n1182));
  XOR2_X1   g757(.A(new_n1182), .B(KEYINPUT47), .Z(new_n1183));
  NAND2_X1  g758(.A1(new_n976), .A2(new_n975), .ZN(new_n1184));
  OAI22_X1  g759(.A1(new_n1184), .A2(new_n978), .B1(G2067), .B2(new_n732), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1176), .B(new_n1183), .C1(new_n987), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1170), .A2(new_n1186), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g762(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1189));
  NAND4_X1  g763(.A1(new_n710), .A2(new_n971), .A3(new_n896), .A4(new_n1189), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


