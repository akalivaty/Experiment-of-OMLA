//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT26), .ZN(new_n203));
  NAND2_X1  g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(KEYINPUT26), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT68), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n214));
  XOR2_X1   g013(.A(new_n213), .B(new_n214), .Z(new_n215));
  NOR2_X1   g014(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT64), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n204), .B1(new_n202), .B2(KEYINPUT23), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  NOR3_X1   g020(.A1(new_n221), .A2(G169gat), .A3(G176gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n224));
  INV_X1    g023(.A(G183gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n212), .A2(G183gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n228), .B2(KEYINPUT24), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n202), .A2(KEYINPUT23), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n221), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n230), .A2(KEYINPUT64), .A3(new_n231), .A4(new_n204), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n223), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n237), .A3(new_n234), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n220), .A2(new_n222), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n229), .A2(new_n240), .A3(KEYINPUT25), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n218), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n233), .A2(new_n237), .A3(new_n234), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n237), .B1(new_n233), .B2(new_n234), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n218), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n217), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT70), .B(G120gat), .ZN(new_n248));
  INV_X1    g047(.A(G113gat), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  INV_X1    g050(.A(G120gat), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT1), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G127gat), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n255), .A2(KEYINPUT69), .A3(G134gat), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n251), .B2(KEYINPUT69), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n249), .B2(new_n252), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n250), .A2(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G227gat), .ZN(new_n261));
  INV_X1    g060(.A(G233gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT66), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n216), .B1(new_n265), .B2(new_n245), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n254), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n257), .A2(new_n258), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n260), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT32), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(G71gat), .B(G99gat), .Z(new_n275));
  XNOR2_X1  g074(.A(new_n275), .B(KEYINPUT72), .ZN(new_n276));
  XNOR2_X1  g075(.A(G15gat), .B(G43gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT71), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n276), .B(new_n278), .Z(new_n279));
  NAND3_X1  g078(.A1(new_n272), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n271), .B(KEYINPUT32), .C1(new_n273), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n263), .B1(new_n260), .B2(new_n270), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n285), .ZN(new_n287));
  AOI211_X1 g086(.A(new_n263), .B(new_n287), .C1(new_n260), .C2(new_n270), .ZN(new_n288));
  OR2_X1    g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(G155gat), .B2(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT78), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G155gat), .B(G162gat), .ZN(new_n295));
  XOR2_X1   g094(.A(G141gat), .B(G148gat), .Z(new_n296));
  AND3_X1   g095(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT2), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT78), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT77), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(KEYINPUT77), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n295), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n297), .A2(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(KEYINPUT22), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n307), .B1(new_n317), .B2(KEYINPUT29), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n305), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n294), .A2(new_n296), .A3(new_n295), .A4(new_n300), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n318), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G228gat), .A2(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(G228gat), .A3(G233gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n308), .A2(KEYINPUT84), .A3(new_n309), .ZN(new_n329));
  INV_X1    g128(.A(new_n317), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT84), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n310), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n328), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(G22gat), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G22gat), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n332), .A2(new_n329), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n326), .B(new_n335), .C1(new_n336), .C2(new_n328), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n338));
  INV_X1    g137(.A(G50gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G78gat), .B(G106gat), .Z(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  AND4_X1   g141(.A1(KEYINPUT85), .A2(new_n334), .A3(new_n337), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT85), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n337), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n345), .A2(new_n342), .B1(new_n334), .B2(new_n337), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n286), .A2(new_n288), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(new_n280), .A3(new_n282), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n290), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n320), .A2(new_n267), .A3(new_n321), .A4(new_n268), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n306), .A2(KEYINPUT79), .A3(new_n259), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n322), .A2(new_n357), .A3(new_n269), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n322), .B2(new_n269), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n355), .B(new_n356), .C1(new_n359), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n352), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n355), .A2(new_n356), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n308), .A2(new_n367), .A3(new_n269), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n306), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n366), .A2(new_n362), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n368), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n371), .A2(KEYINPUT5), .A3(new_n363), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT4), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n306), .A2(KEYINPUT81), .A3(new_n365), .A4(new_n259), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n353), .B2(KEYINPUT4), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n364), .A2(new_n370), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G1gat), .B(G29gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n378), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n378), .A2(new_n382), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(new_n378), .B2(new_n382), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n384), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n217), .A2(new_n264), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n309), .ZN(new_n395));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(new_n396), .B(KEYINPUT76), .Z(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n397), .B(new_n330), .C1(new_n266), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n266), .B2(KEYINPUT29), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n394), .A2(G226gat), .A3(G233gat), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n330), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n393), .B1(new_n401), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n403), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n317), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n400), .A3(new_n392), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n408), .A3(KEYINPUT30), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n407), .A2(new_n410), .A3(new_n400), .A4(new_n392), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT35), .B(new_n389), .C1(new_n409), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n351), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n283), .A2(KEYINPUT73), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT73), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n280), .A2(new_n415), .A3(new_n282), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n289), .A3(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n349), .A2(new_n347), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n389), .B1(new_n409), .B2(new_n411), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n413), .A2(KEYINPUT88), .B1(new_n420), .B2(KEYINPUT35), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT88), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n351), .A2(new_n422), .A3(new_n412), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n280), .A2(new_n415), .A3(new_n282), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n415), .B1(new_n280), .B2(new_n282), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n424), .A2(new_n425), .A3(new_n348), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n349), .A2(KEYINPUT36), .ZN(new_n427));
  OAI21_X1  g226(.A(KEYINPUT75), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT36), .ZN(new_n429));
  INV_X1    g228(.A(new_n290), .ZN(new_n430));
  INV_X1    g229(.A(new_n349), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n417), .A2(new_n433), .A3(KEYINPUT36), .A4(new_n349), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n419), .A2(new_n347), .ZN(new_n436));
  INV_X1    g235(.A(new_n347), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n409), .A2(new_n411), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n376), .A2(new_n374), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n371), .B1(new_n441), .B2(new_n373), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT86), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n442), .A2(new_n443), .A3(new_n362), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n377), .A2(new_n368), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT86), .B1(new_n445), .B2(new_n363), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n440), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n443), .B1(new_n442), .B2(new_n362), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(KEYINPUT86), .A3(new_n363), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n361), .A2(new_n363), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT39), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n451), .A3(new_n382), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT40), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n385), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n447), .A2(new_n451), .A3(KEYINPUT40), .A4(new_n382), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n437), .B1(new_n439), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n393), .A2(KEYINPUT37), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n406), .A2(new_n330), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT37), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n247), .A2(new_n398), .B1(new_n395), .B2(new_n396), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(new_n317), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n405), .A2(new_n458), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n407), .A2(new_n400), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n393), .B1(new_n465), .B2(KEYINPUT37), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n401), .B2(new_n404), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  OAI22_X1  g267(.A1(new_n463), .A2(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n389), .A3(new_n408), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n436), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n421), .A2(new_n423), .B1(new_n435), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT96), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT91), .B1(new_n339), .B2(G43gat), .ZN(new_n475));
  INV_X1    g274(.A(G43gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT90), .B1(new_n476), .B2(G50gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT91), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n476), .A3(G50gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n339), .A3(G43gat), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n475), .A2(new_n477), .A3(new_n479), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n339), .A2(G43gat), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n476), .A2(G50gat), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n486), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT89), .B(G29gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G36gat), .ZN(new_n492));
  NOR2_X1   g291(.A1(G29gat), .A2(G36gat), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n493), .A2(KEYINPUT14), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(KEYINPUT14), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n483), .B1(new_n482), .B2(new_n484), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n497), .A2(new_n496), .ZN(new_n498));
  OAI22_X1  g297(.A1(new_n490), .A2(new_n496), .B1(new_n498), .B2(new_n488), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n474), .B1(new_n499), .B2(KEYINPUT17), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n496), .B1(new_n485), .B2(new_n489), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n497), .A2(new_n496), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n502), .B2(new_n489), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT93), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT16), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n507), .B1(new_n508), .B2(G1gat), .ZN(new_n509));
  INV_X1    g308(.A(G8gat), .ZN(new_n510));
  OAI221_X1 g309(.A(new_n509), .B1(KEYINPUT94), .B2(new_n510), .C1(G1gat), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(KEYINPUT94), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n499), .B2(KEYINPUT17), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT95), .ZN(new_n516));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n513), .A2(new_n503), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT95), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n499), .A2(new_n474), .A3(KEYINPUT17), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT93), .B1(new_n503), .B2(new_n504), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n514), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT18), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G197gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT11), .B(G169gat), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n527), .B(new_n528), .Z(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT12), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n513), .B(new_n503), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n517), .B(KEYINPUT13), .Z(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n535), .B1(new_n523), .B2(new_n524), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n473), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n518), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n519), .B1(new_n506), .B2(new_n514), .ZN(new_n539));
  INV_X1    g338(.A(new_n517), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n541), .A2(KEYINPUT18), .B1(new_n533), .B2(new_n534), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n530), .B1(new_n523), .B2(new_n524), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT96), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n525), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n537), .A2(new_n544), .B1(new_n545), .B2(new_n530), .ZN(new_n546));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G71gat), .B(G78gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT97), .B(KEYINPUT21), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G231gat), .A2(G233gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(G127gat), .B(G155gat), .Z(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n556), .B(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(G183gat), .B(G211gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AND2_X1   g360(.A1(new_n551), .A2(KEYINPUT21), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n513), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT99), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n561), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G85gat), .A2(G92gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT7), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n577), .B(KEYINPUT100), .ZN(new_n582));
  INV_X1    g381(.A(new_n580), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n503), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(KEYINPUT17), .B2(new_n499), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n588), .B1(new_n589), .B2(new_n506), .ZN(new_n590));
  XOR2_X1   g389(.A(G190gat), .B(G218gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT101), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G134gat), .ZN(new_n595));
  INV_X1    g394(.A(G162gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n592), .A2(new_n598), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n585), .A2(new_n551), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n581), .A2(new_n584), .A3(new_n552), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(G230gat), .A2(G233gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n607), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n604), .A2(new_n611), .A3(new_n605), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n585), .A2(KEYINPUT10), .A3(new_n551), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  NAND3_X1  g417(.A1(new_n609), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n618), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n608), .B2(new_n614), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n570), .A2(new_n603), .A3(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n472), .A2(new_n546), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(new_n389), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g426(.A(KEYINPUT16), .B(G8gat), .Z(new_n628));
  AND3_X1   g427(.A1(new_n625), .A2(new_n439), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n510), .B1(new_n625), .B2(new_n439), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT42), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(KEYINPUT42), .B2(new_n629), .ZN(G1325gat));
  INV_X1    g431(.A(new_n435), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n625), .A2(G15gat), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n435), .A2(new_n471), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n420), .A2(KEYINPUT35), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT35), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n419), .A2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT88), .B1(new_n638), .B2(new_n350), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n636), .A2(new_n423), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n635), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n546), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n430), .A2(new_n431), .ZN(new_n643));
  INV_X1    g442(.A(new_n624), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(G15gat), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(KEYINPUT102), .B1(new_n645), .B2(new_n646), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n634), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT103), .ZN(G1326gat));
  NAND2_X1  g449(.A1(new_n625), .A2(new_n437), .ZN(new_n651));
  XNOR2_X1  g450(.A(KEYINPUT43), .B(G22gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(G1327gat));
  NAND3_X1  g452(.A1(new_n569), .A2(new_n602), .A3(new_n623), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT104), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n641), .A2(new_n642), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n389), .ZN(new_n657));
  OR2_X1    g456(.A1(new_n657), .A2(new_n491), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT45), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n641), .B2(new_n602), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(KEYINPUT44), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI211_X1 g466(.A(new_n603), .B(new_n667), .C1(new_n635), .C2(new_n640), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n569), .B(KEYINPUT105), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n671), .A2(new_n546), .A3(new_n622), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n389), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n491), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n661), .A2(new_n674), .ZN(G1328gat));
  INV_X1    g474(.A(G36gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n656), .A2(new_n676), .A3(new_n439), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT46), .Z(new_n678));
  AND3_X1   g477(.A1(new_n669), .A2(new_n439), .A3(new_n672), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n676), .B2(new_n679), .ZN(G1329gat));
  NAND3_X1  g479(.A1(new_n669), .A2(new_n633), .A3(new_n672), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(G43gat), .ZN(new_n682));
  INV_X1    g481(.A(new_n643), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(G43gat), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n641), .A2(new_n642), .A3(new_n655), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT107), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n682), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  NAND2_X1  g490(.A1(new_n641), .A2(new_n602), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n663), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n603), .B1(new_n635), .B2(new_n640), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n664), .A3(new_n666), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n693), .A2(new_n695), .A3(new_n437), .A4(new_n672), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(G50gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n656), .A2(new_n339), .A3(new_n437), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n697), .B2(new_n698), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(G1331gat));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n642), .A2(new_n569), .A3(new_n602), .A4(new_n623), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n472), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n641), .A2(KEYINPUT108), .A3(new_n704), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n657), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT109), .B(G57gat), .Z(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(G1332gat));
  AND2_X1   g510(.A1(new_n706), .A2(new_n707), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n438), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT110), .B1(new_n708), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OR2_X1    g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  NAND3_X1  g519(.A1(new_n706), .A2(new_n643), .A3(new_n707), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(G71gat), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n706), .A2(new_n707), .A3(KEYINPUT111), .A4(new_n643), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n712), .A2(G71gat), .A3(new_n633), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT50), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n726), .A2(new_n730), .A3(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n729), .A2(new_n731), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n712), .A2(new_n437), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g533(.A1(new_n642), .A2(new_n570), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n623), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n693), .A2(new_n695), .A3(new_n389), .A4(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT112), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n574), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(new_n739), .B2(new_n738), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n641), .A2(new_n742), .A3(new_n602), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n735), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n694), .A2(new_n742), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n692), .A2(KEYINPUT113), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n736), .B1(new_n694), .B2(new_n742), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT51), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n389), .A2(new_n574), .A3(new_n622), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n741), .B1(new_n751), .B2(new_n752), .ZN(G1336gat));
  NAND4_X1  g552(.A1(new_n693), .A2(new_n695), .A3(new_n439), .A4(new_n737), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n669), .A2(KEYINPUT114), .A3(new_n439), .A4(new_n737), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n756), .A2(new_n757), .A3(G92gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n438), .A2(G92gat), .A3(new_n623), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n747), .B2(new_n750), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n760), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n745), .B1(new_n744), .B2(new_n746), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n749), .A3(KEYINPUT51), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n754), .A2(G92gat), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT52), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n762), .A2(new_n768), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n669), .A2(new_n633), .A3(new_n737), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(G99gat), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n683), .A2(G99gat), .A3(new_n623), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n751), .B2(new_n772), .ZN(G1338gat));
  NOR3_X1   g572(.A1(new_n347), .A2(G106gat), .A3(new_n623), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT115), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n764), .B2(new_n765), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n693), .A2(new_n695), .A3(new_n437), .A4(new_n737), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT53), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT53), .B1(new_n777), .B2(G106gat), .ZN(new_n780));
  INV_X1    g579(.A(new_n774), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n751), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1339gat));
  NAND3_X1  g582(.A1(new_n612), .A2(new_n613), .A3(new_n610), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT116), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n612), .A2(new_n786), .A3(new_n613), .A4(new_n610), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n614), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n618), .B1(new_n614), .B2(new_n789), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(KEYINPUT55), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n619), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT117), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n793), .A2(new_n796), .A3(new_n619), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(new_n792), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n533), .A2(new_n534), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n516), .A2(new_n518), .A3(new_n522), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n540), .ZN(new_n804));
  INV_X1    g603(.A(new_n529), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n622), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n532), .A2(new_n536), .A3(new_n473), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT96), .B1(new_n542), .B2(new_n543), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n801), .A2(new_n546), .B1(new_n810), .B2(KEYINPUT118), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n810), .A2(KEYINPUT118), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n603), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI221_X1 g612(.A(new_n602), .B1(new_n805), .B2(new_n804), .C1(new_n808), .C2(new_n809), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n801), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n671), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n624), .A2(new_n642), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n439), .A2(new_n657), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n351), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n822), .A2(new_n249), .A3(new_n546), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n417), .A2(new_n418), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n642), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n249), .B2(new_n825), .ZN(G1340gat));
  OAI21_X1  g625(.A(G120gat), .B1(new_n822), .B2(new_n623), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n821), .A2(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n622), .A2(new_n248), .ZN(new_n829));
  XNOR2_X1  g628(.A(new_n829), .B(KEYINPUT119), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(G1341gat));
  OAI21_X1  g630(.A(new_n255), .B1(new_n828), .B2(new_n569), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n670), .A2(new_n255), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n822), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n821), .A2(KEYINPUT120), .A3(new_n351), .A4(new_n834), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n832), .A2(new_n836), .A3(new_n837), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n822), .B2(new_n603), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n603), .A2(G134gat), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT56), .B1(new_n828), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n821), .A2(new_n843), .A3(new_n824), .A4(new_n840), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n839), .A2(new_n842), .A3(new_n844), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n633), .A2(new_n347), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n546), .A2(G141gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n821), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n800), .A2(new_n619), .A3(new_n793), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n806), .B1(new_n537), .B2(new_n544), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n546), .A2(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n851), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n603), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n816), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n818), .B1(new_n856), .B2(new_n569), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT57), .B1(new_n857), .B2(new_n347), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(new_n437), .C1(new_n817), .C2(new_n818), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n435), .A2(new_n820), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n858), .A2(new_n642), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G141gat), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n863), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1344gat));
  NAND3_X1  g667(.A1(new_n819), .A2(new_n820), .A3(new_n846), .ZN(new_n869));
  OR3_X1    g668(.A1(new_n869), .A2(G148gat), .A3(new_n623), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871));
  INV_X1    g670(.A(new_n818), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n810), .A2(KEYINPUT121), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n873), .B(new_n853), .C1(new_n546), .C2(new_n849), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n815), .B1(new_n874), .B2(new_n603), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT122), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n569), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n855), .A2(new_n816), .A3(new_n876), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n347), .A2(KEYINPUT57), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n437), .B1(new_n817), .B2(new_n818), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT57), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n881), .A2(new_n622), .A3(new_n861), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n871), .B1(new_n884), .B2(G148gat), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n871), .A2(G148gat), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n858), .A2(new_n860), .A3(new_n861), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n622), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n870), .B1(new_n885), .B2(new_n888), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n569), .A2(G155gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n821), .A2(new_n846), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n858), .A2(new_n671), .A3(new_n860), .A4(new_n861), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G155gat), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT123), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(new_n596), .B1(new_n869), .B2(new_n603), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n603), .A2(new_n596), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n858), .A2(new_n860), .A3(new_n861), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT124), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n899), .A2(new_n904), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n438), .A2(new_n389), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n819), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n546), .A2(G169gat), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n824), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n351), .B(new_n907), .C1(new_n817), .C2(new_n818), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n546), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n910), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(G1348gat));
  INV_X1    g715(.A(G176gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n908), .A2(new_n824), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n623), .ZN(new_n919));
  INV_X1    g718(.A(new_n912), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(G176gat), .A3(new_n622), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT126), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n921), .A2(KEYINPUT126), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n919), .A2(new_n922), .A3(new_n923), .ZN(G1349gat));
  OAI21_X1  g723(.A(G183gat), .B1(new_n912), .B2(new_n670), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n570), .A2(new_n211), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n819), .A2(new_n824), .A3(new_n907), .A4(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n925), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  OR2_X1    g729(.A1(new_n928), .A2(KEYINPUT60), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n930), .B(new_n931), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n912), .B2(new_n603), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n933), .A2(KEYINPUT61), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n602), .A2(new_n212), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n934), .A2(new_n935), .B1(new_n918), .B2(new_n936), .ZN(G1351gat));
  NAND2_X1  g736(.A1(new_n435), .A2(new_n907), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n819), .A2(new_n437), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n642), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n881), .A2(new_n883), .A3(new_n939), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n642), .A2(G197gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  OAI21_X1  g745(.A(G204gat), .B1(new_n943), .B2(new_n623), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n623), .A2(G204gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT62), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  OR3_X1    g749(.A1(new_n940), .A2(KEYINPUT62), .A3(new_n949), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n947), .A2(new_n950), .A3(new_n951), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n941), .A2(new_n312), .A3(new_n570), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n881), .A2(new_n570), .A3(new_n883), .A4(new_n939), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  OAI21_X1  g756(.A(G218gat), .B1(new_n943), .B2(new_n603), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n941), .A2(new_n313), .A3(new_n602), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1355gat));
endmodule


