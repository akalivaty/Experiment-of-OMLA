//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1266, new_n1267,
    new_n1268, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  INV_X1    g0014(.A(new_n201), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT64), .Z(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(KEYINPUT70), .ZN(new_n246));
  INV_X1    g0046(.A(G200), .ZN(new_n247));
  INV_X1    g0047(.A(G1698), .ZN(new_n248));
  OR2_X1    g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n251), .A2(G223), .B1(new_n254), .B2(G77), .ZN(new_n255));
  INV_X1    g0055(.A(G222), .ZN(new_n256));
  AOI21_X1  g0056(.A(G1698), .B1(new_n249), .B2(new_n250), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(G33), .A2(G41), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G1), .A3(G13), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n264), .A2(new_n266), .A3(G274), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT66), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  INV_X1    g0069(.A(new_n218), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n269), .B1(new_n270), .B2(new_n265), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT66), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(new_n264), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n260), .A2(new_n264), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n268), .A2(new_n273), .B1(G226), .B2(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n247), .B1(new_n261), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT69), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n279), .A2(new_n218), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n209), .A2(G1), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n202), .ZN(new_n285));
  INV_X1    g0085(.A(new_n281), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n283), .A2(new_n285), .B1(new_n202), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n209), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(G150), .ZN(new_n290));
  NOR2_X1   g0090(.A1(G20), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI22_X1  g0092(.A1(new_n288), .A2(new_n289), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G20), .B2(new_n203), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n287), .B1(new_n294), .B2(new_n280), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n261), .A2(G190), .A3(new_n275), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n287), .B(KEYINPUT9), .C1(new_n294), .C2(new_n280), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n297), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n246), .B1(new_n278), .B2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n276), .B(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(new_n301), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(KEYINPUT70), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n276), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n306), .A2(new_n298), .A3(new_n297), .A4(new_n300), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n302), .A2(new_n305), .B1(KEYINPUT10), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n295), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n261), .A2(new_n275), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G179), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n261), .A2(new_n313), .A3(new_n275), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  INV_X1    g0117(.A(G232), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G1698), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(G226), .B2(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n317), .B1(new_n320), .B2(new_n254), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n260), .B1(new_n274), .B2(G238), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n268), .A2(new_n273), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n322), .B2(new_n324), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  INV_X1    g0128(.A(G190), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n280), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n291), .A2(G50), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT71), .ZN(new_n333));
  INV_X1    g0133(.A(G77), .ZN(new_n334));
  OAI22_X1  g0134(.A1(new_n289), .A2(new_n334), .B1(new_n209), .B2(G68), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n331), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT11), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(G68), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n282), .A2(new_n340), .A3(new_n284), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT12), .B1(new_n281), .B2(G68), .ZN(new_n342));
  OR3_X1    g0142(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(new_n339), .A3(new_n344), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n328), .A2(new_n330), .A3(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(G169), .C1(new_n325), .C2(new_n326), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n348), .B1(new_n327), .B2(new_n313), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n347), .B1(new_n327), .B2(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n288), .A2(new_n292), .B1(new_n209), .B2(new_n334), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT15), .B(G87), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n289), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n331), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(new_n356), .B(KEYINPUT67), .ZN(new_n357));
  OAI21_X1  g0157(.A(G77), .B1(new_n209), .B2(G1), .ZN(new_n358));
  OAI22_X1  g0158(.A1(new_n282), .A2(new_n358), .B1(G77), .B2(new_n281), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n251), .A2(G238), .ZN(new_n362));
  INV_X1    g0162(.A(G107), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT3), .B(G33), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n362), .B1(new_n363), .B2(new_n364), .C1(new_n258), .C2(new_n318), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n260), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n268), .A2(new_n273), .B1(G244), .B2(new_n274), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n313), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n311), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n361), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n368), .A2(G200), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n360), .A2(new_n373), .A3(KEYINPUT68), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(G190), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT68), .B1(new_n360), .B2(new_n373), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n372), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n352), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(KEYINPUT7), .B1(new_n254), .B2(new_n209), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NOR4_X1   g0181(.A1(new_n252), .A2(new_n253), .A3(new_n381), .A4(G20), .ZN(new_n382));
  OAI21_X1  g0182(.A(G68), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G58), .A2(G68), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n215), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G20), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT72), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n291), .A2(G159), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n209), .B1(new_n215), .B2(new_n384), .ZN(new_n390));
  INV_X1    g0190(.A(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT72), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n383), .A2(KEYINPUT16), .A3(new_n389), .A4(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n381), .B1(new_n364), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n340), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n386), .A2(new_n388), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n393), .A2(new_n399), .A3(new_n331), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n288), .A2(new_n284), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n282), .B1(KEYINPUT73), .B2(new_n401), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(KEYINPUT73), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n402), .A2(new_n403), .B1(new_n288), .B2(new_n286), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  NOR3_X1   g0205(.A1(new_n260), .A2(new_n264), .A3(new_n318), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n268), .B2(new_n273), .ZN(new_n407));
  OAI211_X1 g0207(.A(G223), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n408));
  OAI211_X1 g0208(.A(G226), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n409));
  INV_X1    g0209(.A(G33), .ZN(new_n410));
  INV_X1    g0210(.A(G87), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n408), .B(new_n409), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n260), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n407), .A2(G179), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n311), .B1(new_n407), .B2(new_n413), .ZN(new_n415));
  OAI21_X1  g0215(.A(KEYINPUT74), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n406), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n324), .A2(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n251), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n266), .B1(new_n419), .B2(new_n408), .ZN(new_n420));
  OAI21_X1  g0220(.A(G169), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n407), .A2(new_n413), .A3(G179), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n405), .A2(new_n416), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT18), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n247), .B1(new_n418), .B2(new_n420), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n407), .A2(new_n413), .A3(new_n329), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT75), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n400), .A4(new_n404), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n400), .A2(new_n404), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n434), .A2(new_n430), .A3(KEYINPUT17), .A4(new_n429), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n405), .A2(new_n416), .A3(new_n424), .A4(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n426), .A2(new_n433), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n316), .A2(new_n379), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT76), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n441), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n263), .A2(G1), .ZN(new_n446));
  XNOR2_X1  g0246(.A(KEYINPUT5), .B(G41), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n271), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(G264), .A3(new_n266), .ZN(new_n452));
  NOR2_X1   g0252(.A1(G250), .A2(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G257), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(new_n454), .B2(G1698), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n364), .B1(G33), .B2(G294), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n448), .B(new_n452), .C1(new_n456), .C2(new_n266), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(G1698), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G250), .B2(G1698), .ZN(new_n461));
  INV_X1    g0261(.A(G294), .ZN(new_n462));
  OAI22_X1  g0262(.A1(new_n461), .A2(new_n254), .B1(new_n410), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n260), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT83), .A3(new_n448), .A4(new_n452), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n459), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT84), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n451), .A2(new_n468), .A3(G264), .A4(new_n266), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n470), .A2(new_n448), .A3(new_n464), .ZN(new_n471));
  AOI22_X1  g0271(.A1(G169), .A2(new_n466), .B1(new_n471), .B2(G179), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n363), .A2(KEYINPUT23), .A3(G20), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT23), .B1(new_n363), .B2(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G116), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n473), .A2(new_n474), .B1(G20), .B2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n209), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT22), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT22), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n364), .A2(new_n479), .A3(new_n209), .A4(G87), .ZN(new_n480));
  AOI211_X1 g0280(.A(KEYINPUT24), .B(new_n476), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT24), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n478), .A2(new_n480), .ZN(new_n483));
  INV_X1    g0283(.A(new_n476), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n331), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT82), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(KEYINPUT82), .B(new_n331), .C1(new_n481), .C2(new_n485), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n286), .A2(KEYINPUT25), .A3(new_n363), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT25), .B1(new_n286), .B2(new_n363), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n280), .B(new_n281), .C1(G1), .C2(new_n410), .ZN(new_n494));
  OAI22_X1  g0294(.A1(new_n492), .A2(new_n493), .B1(new_n494), .B2(new_n363), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n472), .B1(new_n490), .B2(new_n496), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n266), .A2(G274), .A3(new_n446), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT77), .ZN(new_n499));
  OAI21_X1  g0299(.A(G250), .B1(new_n263), .B2(G1), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n260), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n208), .A2(G45), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n266), .A2(KEYINPUT77), .A3(G250), .A4(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(G244), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n505));
  OAI211_X1 g0305(.A(G238), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n475), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n260), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(KEYINPUT78), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT78), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n504), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n313), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n364), .A2(new_n209), .A3(G68), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT19), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n209), .B1(new_n317), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G87), .B2(new_n206), .ZN(new_n517));
  INV_X1    g0317(.A(G97), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n515), .B1(new_n289), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g0320(.A1(new_n520), .A2(new_n331), .B1(new_n286), .B2(new_n354), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n354), .B2(new_n494), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n504), .A2(new_n508), .A3(new_n511), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n511), .B1(new_n504), .B2(new_n508), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n513), .B(new_n522), .C1(new_n525), .C2(G169), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n523), .B2(new_n524), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n510), .A2(G190), .A3(new_n512), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n494), .A2(new_n411), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n497), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT81), .ZN(new_n534));
  AND2_X1   g0334(.A1(G264), .A2(G1698), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n252), .B2(new_n253), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(KEYINPUT79), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT79), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n538), .B(new_n535), .C1(new_n252), .C2(new_n253), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n257), .A2(G257), .B1(new_n254), .B2(G303), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT80), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n260), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n451), .A2(G270), .A3(new_n266), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n448), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(G190), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G116), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n286), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n494), .B2(new_n550), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n279), .A2(new_n218), .B1(G20), .B2(new_n550), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G283), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n554), .B(new_n209), .C1(G33), .C2(new_n518), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n553), .A2(KEYINPUT20), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(KEYINPUT20), .B1(new_n553), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n247), .B1(new_n545), .B2(new_n548), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n534), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n545), .A2(new_n548), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(G200), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n564), .A2(KEYINPUT81), .A3(new_n559), .A4(new_n549), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n559), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n448), .A2(new_n546), .A3(G179), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n545), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(G169), .B1(new_n552), .B2(new_n558), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n540), .A2(new_n541), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(KEYINPUT80), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n266), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n572), .B1(new_n576), .B2(new_n547), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT21), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT21), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n563), .A2(new_n579), .A3(new_n572), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n570), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  OAI211_X1 g0381(.A(G250), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n582));
  OAI211_X1 g0382(.A(G244), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n554), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(KEYINPUT4), .B1(new_n257), .B2(G244), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n260), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n260), .B1(new_n446), .B2(new_n447), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n447), .A2(new_n446), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n588), .A2(G257), .B1(new_n589), .B2(new_n271), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G200), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT6), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n593), .A2(new_n518), .A3(G107), .ZN(new_n594));
  XNOR2_X1  g0394(.A(G97), .B(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n594), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(new_n209), .B1(new_n334), .B2(new_n292), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n363), .B1(new_n395), .B2(new_n396), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n331), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  MUX2_X1   g0399(.A(new_n281), .B(new_n494), .S(G97), .Z(new_n600));
  NAND3_X1  g0400(.A1(new_n587), .A2(new_n590), .A3(G190), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n592), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n591), .A2(new_n311), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(new_n600), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n587), .A2(new_n590), .A3(new_n313), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n470), .A2(new_n448), .A3(new_n464), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n247), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(new_n466), .B2(G190), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n495), .B1(new_n488), .B2(new_n489), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n533), .A2(new_n566), .A3(new_n581), .A4(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n445), .A2(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n421), .A2(new_n423), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n405), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(KEYINPUT18), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n405), .A2(new_n615), .A3(new_n436), .ZN(new_n618));
  INV_X1    g0418(.A(new_n372), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n346), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n351), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n433), .A2(new_n435), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n617), .B(new_n618), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n302), .A2(new_n305), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n307), .A2(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n315), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n509), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n513), .B(new_n522), .C1(G169), .C2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n532), .A2(new_n606), .ZN(new_n631));
  XNOR2_X1  g0431(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n528), .B(new_n530), .C1(new_n247), .C2(new_n628), .ZN(new_n634));
  INV_X1    g0434(.A(new_n606), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n629), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n630), .B1(new_n633), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n579), .B1(new_n563), .B2(new_n572), .ZN(new_n640));
  AOI211_X1 g0440(.A(KEYINPUT21), .B(new_n571), .C1(new_n545), .C2(new_n548), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n569), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n497), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n476), .B1(new_n478), .B2(new_n480), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n644), .B(new_n482), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT82), .B1(new_n645), .B2(new_n331), .ZN(new_n646));
  INV_X1    g0446(.A(new_n489), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n610), .B(new_n496), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n602), .A2(new_n606), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n629), .A4(new_n634), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT85), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n643), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n648), .A2(new_n649), .A3(new_n629), .A4(new_n634), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n490), .A2(new_n496), .ZN(new_n654));
  INV_X1    g0454(.A(new_n472), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n581), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT85), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n639), .B1(new_n652), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n627), .B1(new_n445), .B2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G343), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OR3_X1    g0468(.A1(new_n611), .A2(KEYINPUT87), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT87), .B1(new_n611), .B2(new_n668), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n669), .A2(new_n648), .A3(new_n656), .A4(new_n670), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n671), .A2(new_n581), .A3(new_n667), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n667), .B(KEYINPUT88), .Z(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n497), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT89), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n672), .A2(KEYINPUT89), .A3(new_n675), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n566), .B(new_n581), .C1(new_n559), .C2(new_n668), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n642), .A2(new_n567), .A3(new_n667), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n671), .B1(new_n656), .B2(new_n668), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n680), .A2(new_n687), .ZN(G399));
  INV_X1    g0488(.A(new_n212), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(G41), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G1), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n216), .B2(new_n691), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT28), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT94), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n613), .B2(new_n673), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n648), .A2(new_n649), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n698), .A2(new_n497), .A3(new_n532), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n642), .B1(new_n562), .B2(new_n565), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT94), .A4(new_n674), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n470), .A2(new_n568), .A3(new_n464), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n587), .A2(KEYINPUT30), .A3(new_n590), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n525), .A2(new_n545), .A3(new_n704), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT92), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n576), .A2(new_n703), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(KEYINPUT92), .A3(new_n525), .A4(new_n705), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n591), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n525), .A2(new_n545), .A3(new_n704), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(KEYINPUT91), .B(KEYINPUT30), .Z(new_n714));
  AOI21_X1  g0514(.A(G179), .B1(new_n504), .B2(new_n508), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n608), .A2(new_n591), .A3(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n713), .A2(new_n714), .B1(new_n563), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(KEYINPUT90), .B(KEYINPUT31), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n718), .A2(new_n673), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n667), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n668), .B1(new_n711), .B2(new_n717), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT93), .B1(new_n725), .B2(KEYINPUT31), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n720), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n681), .B1(new_n702), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n651), .B1(new_n643), .B2(new_n650), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n653), .A2(new_n657), .A3(KEYINPUT85), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n673), .B1(new_n731), .B2(new_n639), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n653), .A2(new_n657), .ZN(new_n734));
  OAI22_X1  g0534(.A1(new_n631), .A2(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(new_n629), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(new_n668), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT29), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n728), .B1(new_n733), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n695), .B1(new_n740), .B2(G1), .ZN(G364));
  AND2_X1   g0541(.A1(new_n209), .A2(G13), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n208), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n690), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n212), .A2(new_n364), .ZN(new_n746));
  INV_X1    g0546(.A(G355), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n746), .A2(new_n747), .B1(G116), .B2(new_n212), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n689), .A2(new_n364), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n750), .B1(new_n263), .B2(new_n217), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n241), .A2(new_n263), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n218), .B1(G20), .B2(new_n311), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n745), .B1(new_n753), .B2(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n329), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n209), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n209), .A2(new_n313), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  AOI22_X1  g0566(.A1(G97), .A2(new_n763), .B1(new_n766), .B2(G68), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n768), .A2(KEYINPUT96), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n209), .A2(G179), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n770), .A2(new_n329), .A3(G200), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT95), .Z(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G107), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n768), .A2(KEYINPUT96), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n769), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n764), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G58), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n764), .A2(G190), .A3(new_n247), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n364), .B1(new_n777), .B2(new_n334), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n770), .A2(new_n776), .ZN(new_n781));
  INV_X1    g0581(.A(G159), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT32), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n765), .A2(new_n329), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n785), .B2(new_n202), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n411), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n782), .ZN(new_n789));
  OR4_X1    g0589(.A1(new_n780), .A2(new_n786), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  INV_X1    g0591(.A(new_n779), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n766), .A2(new_n791), .B1(new_n792), .B2(G322), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT97), .Z(new_n794));
  NAND2_X1  g0594(.A1(new_n772), .A2(G283), .ZN(new_n795));
  INV_X1    g0595(.A(G311), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n254), .B1(new_n777), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n781), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(G329), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n784), .A2(G326), .ZN(new_n800));
  INV_X1    g0600(.A(new_n787), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n763), .A2(G294), .B1(new_n801), .B2(G303), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n795), .A2(new_n799), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n775), .A2(new_n790), .B1(new_n794), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n760), .B1(new_n804), .B2(new_n757), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n682), .A2(new_n683), .ZN(new_n806));
  INV_X1    g0606(.A(new_n756), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n684), .A2(new_n745), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n806), .A2(G330), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(G396));
  INV_X1    g0611(.A(new_n777), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n792), .A2(G143), .B1(new_n812), .B2(G159), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n784), .A2(G137), .ZN(new_n814));
  INV_X1    g0614(.A(new_n766), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n814), .C1(new_n290), .C2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n772), .A2(G68), .ZN(new_n820));
  INV_X1    g0620(.A(G132), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n364), .B1(new_n781), .B2(new_n821), .C1(new_n762), .C2(new_n778), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G50), .B2(new_n801), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n818), .A2(new_n819), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n779), .A2(new_n462), .B1(new_n781), .B2(new_n796), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n364), .B(new_n825), .C1(G116), .C2(new_n812), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n772), .A2(G87), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n763), .A2(G97), .B1(new_n801), .B2(G107), .ZN(new_n828));
  AOI22_X1  g0628(.A1(G283), .A2(new_n766), .B1(new_n784), .B2(G303), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n826), .A2(new_n827), .A3(new_n828), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n757), .A2(new_n754), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n831), .A2(new_n757), .B1(new_n334), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n372), .A2(new_n667), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n376), .A2(new_n377), .B1(new_n360), .B2(new_n668), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n372), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n833), .B1(new_n836), .B2(new_n755), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n745), .ZN(new_n838));
  INV_X1    g0638(.A(new_n728), .ZN(new_n839));
  INV_X1    g0639(.A(new_n836), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n660), .B2(new_n673), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n659), .A2(new_n674), .A3(new_n836), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n690), .B2(new_n744), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n838), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT98), .Z(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(G384));
  INV_X1    g0648(.A(new_n596), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(G116), .A3(new_n219), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  NAND3_X1  g0653(.A1(new_n217), .A2(G77), .A3(new_n384), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n202), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n208), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n389), .A2(new_n392), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n394), .B1(new_n858), .B2(new_n397), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(new_n393), .A3(new_n331), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n665), .B1(new_n860), .B2(new_n404), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n438), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  INV_X1    g0663(.A(new_n665), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n405), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n429), .A2(new_n400), .A3(new_n404), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n425), .A2(new_n863), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n429), .A2(new_n400), .A3(new_n404), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n860), .A2(new_n404), .B1(new_n421), .B2(new_n423), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n868), .A2(new_n869), .A3(new_n861), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n867), .B1(new_n870), .B2(new_n863), .ZN(new_n871));
  AND3_X1   g0671(.A1(new_n862), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT38), .B1(new_n862), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n345), .A2(new_n667), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n346), .A2(new_n351), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n346), .B2(new_n351), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n834), .ZN(new_n880));
  AOI211_X1 g0680(.A(new_n874), .B(new_n879), .C1(new_n842), .C2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  INV_X1    g0682(.A(new_n865), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n617), .A2(new_n618), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n622), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n616), .A2(new_n865), .A3(new_n866), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n867), .B1(new_n886), .B2(new_n863), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n882), .B1(new_n872), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n862), .A2(new_n871), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n862), .A2(new_n871), .A3(KEYINPUT38), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n351), .A2(new_n667), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n884), .A2(new_n665), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR3_X1   g0699(.A1(new_n881), .A2(KEYINPUT99), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT99), .ZN(new_n901));
  AND2_X1   g0701(.A1(new_n897), .A2(new_n898), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n842), .A2(new_n880), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n892), .A2(new_n893), .ZN(new_n904));
  INV_X1    g0704(.A(new_n879), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n901), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n444), .A2(new_n733), .A3(new_n739), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n627), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n908), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n719), .A2(KEYINPUT101), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n718), .B2(new_n667), .ZN(new_n913));
  NAND2_X1  g0713(.A1(KEYINPUT90), .A2(KEYINPUT101), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n723), .ZN(new_n915));
  AOI211_X1 g0715(.A(new_n668), .B(new_n915), .C1(new_n711), .C2(new_n717), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n702), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n836), .B1(new_n877), .B2(new_n878), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n904), .A3(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n920), .B1(new_n702), .B2(new_n918), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT40), .ZN(new_n926));
  INV_X1    g0726(.A(new_n888), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n927), .B2(new_n893), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n922), .A2(new_n924), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n444), .A3(new_n919), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n917), .B1(new_n697), .B2(new_n701), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n923), .B1(new_n925), .B2(new_n904), .ZN(new_n932));
  OAI21_X1  g0732(.A(KEYINPUT40), .B1(new_n872), .B2(new_n888), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n931), .A2(new_n933), .A3(new_n920), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n445), .A2(new_n931), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n930), .A2(G330), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n911), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n208), .B2(new_n742), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n911), .A2(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n857), .B1(new_n938), .B2(new_n939), .ZN(G367));
  AOI21_X1  g0740(.A(new_n607), .B1(new_n604), .B2(new_n673), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT104), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n635), .A2(new_n673), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n686), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT106), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n629), .A2(new_n530), .A3(new_n668), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT102), .Z(new_n949));
  OAI211_X1 g0749(.A(new_n629), .B(new_n634), .C1(new_n530), .C2(new_n668), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT103), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n947), .B(new_n955), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n957));
  INV_X1    g0757(.A(new_n945), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n672), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT105), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n606), .B1(new_n943), .B2(new_n656), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n674), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n957), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n956), .B(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n690), .B(KEYINPUT41), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n581), .A2(new_n667), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n672), .B1(new_n685), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(new_n684), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n740), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT108), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n679), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT89), .B1(new_n672), .B2(new_n675), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n945), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT45), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(new_n680), .B2(new_n945), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n678), .A2(KEYINPUT44), .A3(new_n679), .A4(new_n958), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n979), .A2(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n687), .B1(new_n984), .B2(KEYINPUT107), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n979), .A2(new_n980), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n982), .A2(new_n983), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n687), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT107), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n974), .A2(new_n985), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n968), .B1(new_n991), .B2(new_n740), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n967), .B1(new_n992), .B2(new_n744), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n954), .A2(new_n807), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n758), .B1(new_n212), .B2(new_n354), .C1(new_n750), .C2(new_n237), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n745), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n792), .A2(G150), .B1(new_n798), .B2(G137), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n997), .B(new_n364), .C1(new_n202), .C2(new_n777), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n815), .A2(new_n782), .B1(new_n334), .B2(new_n771), .ZN(new_n999));
  INV_X1    g0799(.A(G143), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n785), .A2(new_n1000), .B1(new_n340), .B2(new_n762), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n787), .A2(new_n778), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT109), .Z(new_n1004));
  OAI22_X1  g0804(.A1(new_n785), .A2(new_n796), .B1(new_n363), .B2(new_n762), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n815), .A2(new_n462), .B1(new_n518), .B2(new_n771), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(G283), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n777), .A2(new_n1008), .B1(new_n781), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G303), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n254), .B1(new_n779), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT46), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n801), .A2(G116), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1010), .B(new_n1012), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1007), .B(new_n1015), .C1(new_n1013), .C2(new_n1014), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1004), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n996), .B1(new_n1018), .B2(new_n757), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n994), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n993), .A2(new_n1020), .ZN(G387));
  OR2_X1    g0821(.A1(new_n685), .A2(new_n807), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n746), .A2(new_n692), .B1(G107), .B2(new_n212), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n234), .A2(new_n263), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n692), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G45), .B(new_n1025), .C1(G68), .C2(G77), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n288), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n750), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1023), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n745), .B1(new_n1030), .B2(new_n759), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT110), .B(G150), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n779), .A2(new_n202), .B1(new_n781), .B2(new_n1032), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n254), .B(new_n1033), .C1(G68), .C2(new_n812), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n772), .A2(G97), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n354), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1036), .A2(new_n763), .B1(new_n784), .B2(G159), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n288), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n766), .A2(new_n1038), .B1(new_n801), .B2(G77), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1034), .A2(new_n1035), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n364), .B1(new_n798), .B2(G326), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n792), .A2(G317), .B1(new_n812), .B2(G303), .ZN(new_n1042));
  INV_X1    g0842(.A(G322), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1042), .B1(new_n815), .B2(new_n796), .C1(new_n1043), .C2(new_n785), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n763), .A2(G283), .B1(new_n801), .B2(G294), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT111), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(KEYINPUT111), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1041), .B1(new_n550), .B2(new_n771), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1040), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1031), .B1(new_n1056), .B2(new_n757), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n971), .A2(new_n744), .B1(new_n1022), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n690), .B1(new_n740), .B2(new_n971), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n974), .B2(new_n1059), .ZN(G393));
  AND2_X1   g0860(.A1(new_n991), .A2(new_n690), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n988), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n984), .A2(new_n687), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT114), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1064), .A2(new_n1065), .A3(new_n973), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n986), .A2(new_n987), .A3(new_n687), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n973), .B1(new_n1067), .B2(new_n988), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(KEYINPUT114), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1061), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n958), .A2(new_n756), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n749), .A2(new_n244), .ZN(new_n1073));
  OAI211_X1 g0873(.A(new_n1073), .B(new_n758), .C1(new_n518), .C2(new_n212), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT112), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT112), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1075), .A2(new_n745), .A3(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n254), .B1(new_n781), .B2(new_n1043), .C1(new_n1008), .C2(new_n787), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n772), .B2(G107), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT113), .Z(new_n1080));
  OAI22_X1  g0880(.A1(new_n785), .A2(new_n1009), .B1(new_n796), .B2(new_n779), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT52), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n766), .A2(G303), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n763), .A2(G116), .B1(new_n812), .B2(G294), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G150), .A2(new_n784), .B1(new_n792), .B2(G159), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT51), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n815), .A2(new_n202), .B1(new_n340), .B2(new_n787), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G77), .B2(new_n763), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n364), .B1(new_n781), .B2(new_n1000), .C1(new_n288), .C2(new_n777), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n827), .A3(new_n1091), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1080), .A2(new_n1085), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1077), .B1(new_n1093), .B2(new_n757), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1072), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1064), .B2(new_n743), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1071), .A2(new_n1097), .ZN(G390));
  AOI21_X1  g0898(.A(new_n681), .B1(new_n702), .B2(new_n918), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n444), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n909), .A2(new_n1100), .A3(new_n627), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n702), .A2(new_n727), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(G330), .A3(new_n921), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n835), .A2(new_n372), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n880), .B1(new_n737), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n905), .B1(new_n1099), .B2(new_n836), .ZN(new_n1109));
  OAI21_X1  g0909(.A(KEYINPUT115), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n919), .A2(G330), .A3(new_n836), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n879), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1106), .B1(new_n728), .B2(new_n921), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1099), .A2(new_n921), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n681), .B(new_n840), .C1(new_n702), .C2(new_n727), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n905), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n903), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1101), .B1(new_n1116), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n889), .A2(new_n894), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n879), .B1(new_n842), .B2(new_n880), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n896), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n896), .B1(new_n927), .B2(new_n893), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1107), .B2(new_n879), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1124), .A2(new_n1103), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1117), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT116), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n691), .B1(new_n1121), .B2(new_n1129), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n896), .B1(new_n903), .B2(new_n905), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1122), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1103), .B(new_n1126), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n834), .B1(new_n732), .B2(new_n836), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n895), .B1(new_n1135), .B2(new_n879), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1106), .A2(new_n905), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1136), .A2(new_n1122), .B1(new_n1137), .B2(new_n1125), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1134), .B1(new_n1138), .B2(new_n1117), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT116), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1110), .A2(new_n1115), .B1(new_n903), .B2(new_n1119), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1139), .B(new_n1140), .C1(new_n1141), .C2(new_n1101), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1130), .A2(new_n1131), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1122), .A2(new_n754), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n832), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n745), .B1(new_n1038), .B2(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n779), .A2(new_n550), .B1(new_n777), .B2(new_n518), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n364), .B(new_n1147), .C1(G294), .C2(new_n798), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n788), .B1(G77), .B2(new_n763), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G107), .A2(new_n766), .B1(new_n784), .B2(G283), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1148), .A2(new_n820), .A3(new_n1149), .A4(new_n1150), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n787), .A2(new_n1032), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT53), .Z(new_n1153));
  AOI22_X1  g0953(.A1(G159), .A2(new_n763), .B1(new_n784), .B2(G128), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n254), .B1(new_n792), .B2(G132), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n812), .A2(new_n1157), .B1(new_n798), .B2(G125), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n771), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n766), .A2(G137), .B1(new_n1159), .B2(G50), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1154), .A2(new_n1155), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1151), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1146), .B1(new_n1162), .B2(new_n757), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1129), .A2(new_n744), .B1(new_n1144), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1143), .A2(new_n1164), .ZN(G378));
  NAND3_X1  g0965(.A1(new_n902), .A2(new_n906), .A3(new_n901), .ZN(new_n1166));
  OAI21_X1  g0966(.A(KEYINPUT99), .B1(new_n881), .B2(new_n899), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n315), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n309), .A2(new_n665), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n626), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n308), .B2(new_n315), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1171), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n929), .B2(G330), .ZN(new_n1178));
  NOR4_X1   g0978(.A1(new_n932), .A2(new_n934), .A3(new_n681), .A4(new_n1176), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1166), .B(new_n1167), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n922), .A2(new_n924), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n919), .A2(new_n921), .A3(new_n928), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1181), .A2(G330), .A3(new_n1177), .A4(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n931), .A2(new_n874), .A3(new_n920), .ZN(new_n1184));
  OAI211_X1 g0984(.A(G330), .B(new_n1182), .C1(new_n1184), .C2(new_n923), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1176), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1183), .B(new_n1186), .C1(new_n900), .C2(new_n907), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1101), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1190), .A3(KEYINPUT57), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n691), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1186), .A2(KEYINPUT119), .A3(new_n1183), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(KEYINPUT120), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n908), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1186), .A2(new_n1183), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT120), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1167), .B2(new_n1166), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT119), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1196), .A2(new_n1190), .A3(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1188), .A2(new_n1190), .A3(KEYINPUT121), .A4(KEYINPUT57), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1193), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n784), .A2(G125), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n815), .B2(new_n821), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n792), .A2(G128), .B1(new_n812), .B2(G137), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n787), .B2(new_n1156), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1208), .B(new_n1210), .C1(G150), .C2(new_n763), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1159), .A2(G159), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n254), .A2(new_n262), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(new_n801), .B2(G77), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT117), .Z(new_n1220));
  AOI22_X1  g1020(.A1(new_n792), .A2(G107), .B1(new_n798), .B2(G283), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n354), .B2(new_n777), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n763), .A2(G68), .B1(new_n1159), .B2(G58), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n1223), .B1(new_n518), .B2(new_n815), .C1(new_n550), .C2(new_n785), .ZN(new_n1224));
  NOR3_X1   g1024(.A1(new_n1220), .A2(new_n1222), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1218), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1225), .A2(KEYINPUT58), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1217), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n757), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT118), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1231), .B(new_n745), .C1(G50), .C2(new_n1145), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(new_n1176), .B2(new_n754), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1196), .A2(new_n1201), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n744), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1206), .A2(new_n1235), .ZN(G375));
  NOR2_X1   g1036(.A1(new_n1141), .A2(new_n743), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n879), .A2(new_n754), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n745), .B1(G68), .B2(new_n1145), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n777), .A2(new_n363), .B1(new_n781), .B2(new_n1011), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n364), .B(new_n1240), .C1(G283), .C2(new_n792), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n772), .A2(G77), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n763), .A2(new_n1036), .B1(new_n801), .B2(G97), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G116), .A2(new_n766), .B1(new_n784), .B2(G294), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n364), .B1(new_n771), .B2(new_n778), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1246), .B(KEYINPUT122), .Z(new_n1247));
  AOI22_X1  g1047(.A1(G132), .A2(new_n784), .B1(new_n766), .B2(new_n1157), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n792), .A2(G137), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G150), .A2(new_n812), .B1(new_n798), .B2(G128), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n763), .A2(G50), .B1(new_n801), .B2(G159), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .A4(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1245), .B1(new_n1247), .B2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1239), .B1(new_n1253), .B2(new_n757), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1237), .B1(new_n1238), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1121), .A2(new_n968), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1141), .A2(new_n1101), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(G381));
  OR2_X1    g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NOR4_X1   g1061(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1143), .A2(new_n1164), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1262), .A2(new_n993), .A3(new_n1020), .A4(new_n1263), .ZN(new_n1264));
  OR2_X1    g1064(.A1(new_n1264), .A2(G375), .ZN(G407));
  NAND2_X1  g1065(.A1(new_n666), .A2(G213), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1263), .A2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(G407), .B(G213), .C1(G375), .C2(new_n1268), .ZN(G409));
  AOI21_X1  g1069(.A(new_n1096), .B1(new_n1061), .B2(new_n1070), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G390), .A2(new_n993), .A3(new_n1020), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1261), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT125), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1273), .A2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1261), .A2(KEYINPUT125), .A3(new_n1274), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1277), .A2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(new_n1280), .A3(new_n1272), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT123), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n968), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1196), .A2(new_n1190), .A3(new_n1284), .A4(new_n1201), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1233), .B1(new_n1188), .B2(new_n744), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1283), .B1(new_n1263), .B2(new_n1287), .ZN(new_n1288));
  AND4_X1   g1088(.A1(new_n1283), .A2(new_n1287), .A3(new_n1143), .A4(new_n1164), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1206), .A2(G378), .A3(new_n1235), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1267), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT60), .B1(new_n1141), .B2(new_n1101), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1293), .A2(new_n1258), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1101), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n690), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1255), .B1(new_n1294), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G384), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n847), .B(new_n1255), .C1(new_n1294), .C2(new_n1296), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1267), .A2(G2897), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1302), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1298), .A2(G2897), .A3(new_n1267), .A4(new_n1299), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT124), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1307), .A3(new_n1304), .ZN(new_n1308));
  AND3_X1   g1108(.A1(new_n1206), .A2(G378), .A3(new_n1235), .ZN(new_n1309));
  AND2_X1   g1109(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT123), .B1(new_n1310), .B2(G378), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1287), .A2(new_n1283), .A3(new_n1143), .A4(new_n1164), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1266), .B1(new_n1309), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1306), .A2(new_n1308), .A3(new_n1314), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1266), .B(new_n1300), .C1(new_n1309), .C2(new_n1313), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1282), .A2(new_n1301), .A3(new_n1315), .A4(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT61), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1320), .B1(new_n1292), .B2(new_n1305), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1322));
  OR2_X1    g1122(.A1(new_n1316), .A2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(new_n1316), .B2(new_n1322), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1321), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1278), .A2(new_n1281), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1319), .B1(new_n1326), .B2(new_n1327), .ZN(G405));
  AOI21_X1  g1128(.A(G378), .B1(new_n1206), .B2(new_n1235), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1330), .A2(new_n1299), .A3(new_n1298), .A4(new_n1291), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1300), .B1(new_n1309), .B2(new_n1329), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(KEYINPUT127), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT127), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1331), .A2(new_n1335), .A3(new_n1332), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1334), .A2(new_n1281), .A3(new_n1278), .A4(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1327), .A2(new_n1335), .A3(new_n1332), .A4(new_n1331), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(G402));
endmodule


