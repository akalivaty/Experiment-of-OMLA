//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT86), .B(G22gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  AOI211_X1 g007(.A(KEYINPUT72), .B(KEYINPUT22), .C1(G211gat), .C2(G218gat), .ZN(new_n209));
  AOI21_X1  g008(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n208), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  XOR2_X1   g012(.A(G211gat), .B(G218gat), .Z(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n213), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT73), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT29), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT73), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n219), .A3(new_n214), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(G155gat), .B(G162gat), .Z(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G141gat), .B(G148gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(new_n229), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n224), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G155gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT80), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G155gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G162gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT2), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g041(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(KEYINPUT79), .A2(G148gat), .ZN(new_n244));
  OAI21_X1  g043(.A(G141gat), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n226), .ZN(new_n246));
  INV_X1    g045(.A(new_n224), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n242), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n235), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n220), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n248), .A3(new_n222), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n218), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G228gat), .ZN(new_n257));
  INV_X1    g056(.A(G233gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n217), .A2(new_n220), .B1(new_n218), .B2(new_n252), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT87), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n250), .A2(new_n256), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT31), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n233), .A2(new_n229), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT2), .B1(new_n233), .B2(new_n229), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n224), .B1(new_n226), .B2(new_n245), .ZN(new_n267));
  AOI22_X1  g066(.A1(new_n266), .A2(new_n224), .B1(new_n267), .B2(new_n242), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n216), .A2(KEYINPUT29), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(new_n222), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n270), .A2(new_n260), .B1(new_n257), .B2(new_n258), .ZN(new_n271));
  AND3_X1   g070(.A1(new_n262), .A2(new_n263), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n263), .B1(new_n262), .B2(new_n271), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n207), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n262), .A2(new_n271), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT31), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n262), .A2(new_n263), .A3(new_n271), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n206), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT74), .ZN(new_n280));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OR3_X1    g085(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n282), .A2(new_n283), .A3(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n286), .A2(new_n290), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n288), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  INV_X1    g096(.A(G169gat), .ZN(new_n298));
  INV_X1    g097(.A(G176gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n296), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n283), .ZN(new_n304));
  NAND3_X1  g103(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n304), .B(new_n305), .C1(new_n306), .C2(KEYINPUT65), .ZN(new_n307));
  AND2_X1   g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT65), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT24), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n302), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(KEYINPUT68), .A2(KEYINPUT24), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n291), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(KEYINPUT68), .B2(KEYINPUT24), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT69), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n304), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n303), .B2(new_n283), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n315), .B(new_n316), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n300), .A2(new_n301), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n296), .A2(KEYINPUT67), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT67), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n312), .B1(new_n288), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g123(.A1(new_n321), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n313), .A2(KEYINPUT66), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n309), .B1(new_n308), .B2(KEYINPUT24), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n306), .A2(KEYINPUT65), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n304), .A4(new_n305), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT25), .B1(new_n329), .B2(new_n302), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT66), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n295), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n281), .B1(new_n333), .B2(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(new_n320), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n335), .B1(new_n330), .B2(new_n331), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n313), .A2(KEYINPUT66), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n294), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n281), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n280), .B1(new_n334), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n339), .B1(new_n338), .B2(new_n218), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(KEYINPUT74), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n251), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n251), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n333), .A2(new_n281), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n344), .A2(KEYINPUT75), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n349), .B(new_n251), .C1(new_n341), .C2(new_n343), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT76), .ZN(new_n352));
  XNOR2_X1  g151(.A(G8gat), .B(G36gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n348), .A2(KEYINPUT30), .A3(new_n350), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n347), .A2(new_n345), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT74), .B1(new_n342), .B2(new_n346), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n334), .A2(new_n280), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n345), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n357), .B1(new_n360), .B2(new_n349), .ZN(new_n361));
  INV_X1    g160(.A(new_n350), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n344), .A2(KEYINPUT75), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n365), .A2(new_n350), .A3(new_n357), .A4(new_n355), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT77), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n348), .A2(new_n368), .A3(new_n350), .A4(new_n355), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT30), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G134gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G127gat), .ZN(new_n374));
  INV_X1    g173(.A(G127gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G134gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(KEYINPUT1), .ZN(new_n379));
  INV_X1    g178(.A(G120gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G113gat), .ZN(new_n381));
  INV_X1    g180(.A(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(G127gat), .B(G134gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(new_n235), .A3(new_n248), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n388), .A2(new_n235), .A3(new_n248), .A4(KEYINPUT82), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(KEYINPUT4), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g193(.A(new_n388), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n252), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n389), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G225gat), .A2(G233gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT81), .Z(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n393), .A2(new_n396), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n252), .A2(new_n395), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n405), .A2(new_n394), .B1(new_n397), .B2(new_n389), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n406), .A2(KEYINPUT83), .A3(new_n393), .A4(new_n401), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT5), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n388), .A2(new_n235), .A3(new_n248), .A4(KEYINPUT4), .ZN(new_n410));
  INV_X1    g209(.A(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n405), .B2(new_n394), .ZN(new_n413));
  AOI21_X1  g212(.A(KEYINPUT82), .B1(new_n268), .B2(new_n388), .ZN(new_n414));
  INV_X1    g213(.A(new_n392), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n397), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n409), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  OAI22_X1  g216(.A1(new_n414), .A2(new_n415), .B1(new_n268), .B2(new_n388), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n400), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(G1gat), .B(G29gat), .ZN(new_n421));
  INV_X1    g220(.A(G85gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n421), .B(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT0), .B(G57gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n423), .B(new_n424), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n420), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n420), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n425), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n408), .A2(new_n420), .A3(new_n432), .A4(new_n426), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n428), .A2(new_n430), .A3(new_n431), .A4(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n429), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n425), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n430), .B2(new_n431), .ZN(new_n437));
  AND3_X1   g236(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n279), .B1(new_n372), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  XNOR2_X1  g240(.A(G15gat), .B(G43gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(G71gat), .B(G99gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  XOR2_X1   g244(.A(new_n445), .B(KEYINPUT64), .Z(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n338), .A2(new_n395), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n388), .B(new_n294), .C1(new_n336), .C2(new_n337), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n444), .B1(new_n450), .B2(KEYINPUT33), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT32), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n447), .A3(new_n449), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(KEYINPUT34), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n449), .ZN(new_n457));
  AOI221_X4 g256(.A(new_n452), .B1(KEYINPUT33), .B2(new_n444), .C1(new_n457), .C2(new_n446), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n454), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT34), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n455), .B(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n326), .A2(new_n332), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n388), .B1(new_n462), .B2(new_n294), .ZN(new_n463));
  INV_X1    g262(.A(new_n449), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n446), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n468), .A3(new_n444), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n453), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n461), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n441), .B1(new_n459), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n456), .B1(new_n454), .B2(new_n458), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n471), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n473), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n202), .B1(new_n440), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n477), .A2(new_n473), .ZN(new_n480));
  INV_X1    g279(.A(new_n475), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n469), .A2(new_n470), .A3(new_n461), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT71), .B1(new_n474), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n484), .B2(new_n473), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT30), .B1(new_n367), .B2(new_n369), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n486), .A2(new_n438), .A3(new_n364), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n485), .B(KEYINPUT88), .C1(new_n487), .C2(new_n279), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n418), .A2(new_n400), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(KEYINPUT89), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n411), .B1(new_n406), .B2(new_n393), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n491), .B1(new_n494), .B2(new_n490), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n425), .B1(new_n492), .B2(new_n489), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT40), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT92), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n495), .A2(new_n500), .A3(KEYINPUT40), .A4(new_n496), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n499), .A2(new_n501), .B1(new_n498), .B2(new_n497), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n404), .A2(new_n407), .B1(new_n417), .B2(new_n419), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n425), .B1(new_n503), .B2(KEYINPUT90), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n408), .A2(new_n420), .A3(KEYINPUT90), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT91), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n426), .B1(new_n429), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(KEYINPUT90), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n502), .B(new_n512), .C1(new_n486), .C2(new_n364), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n428), .A2(new_n431), .A3(new_n433), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n506), .B2(new_n511), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n437), .A2(new_n435), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT94), .B(KEYINPUT37), .Z(new_n519));
  NAND4_X1  g318(.A1(new_n365), .A2(new_n350), .A3(new_n357), .A4(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(KEYINPUT95), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT93), .B(KEYINPUT38), .Z(new_n522));
  OAI21_X1  g321(.A(new_n345), .B1(new_n341), .B2(new_n343), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(new_n347), .B2(new_n251), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n348), .A2(new_n527), .A3(new_n350), .A4(new_n519), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n521), .A2(new_n526), .A3(new_n354), .A4(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n516), .A2(new_n518), .A3(new_n529), .A4(new_n370), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT37), .B1(new_n361), .B2(new_n362), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n521), .A2(new_n354), .A3(new_n528), .A4(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n279), .B(new_n513), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n479), .A2(new_n488), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT35), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n515), .B2(new_n517), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n472), .A2(new_n279), .A3(new_n475), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n372), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n279), .A2(new_n477), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n372), .A2(new_n439), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n543), .B2(new_n536), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n535), .A2(KEYINPUT96), .A3(new_n544), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT99), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT99), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(G29gat), .B2(G36gat), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT14), .ZN(new_n554));
  OR3_X1    g353(.A1(new_n550), .A2(KEYINPUT99), .A3(KEYINPUT14), .ZN(new_n555));
  NAND2_X1  g354(.A1(G29gat), .A2(G36gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G43gat), .B(G50gat), .Z(new_n558));
  AOI21_X1  g357(.A(new_n557), .B1(KEYINPUT100), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n558), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(KEYINPUT15), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n561), .B1(KEYINPUT15), .B2(new_n559), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G22gat), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT16), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(G1gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G1gat), .B2(new_n563), .ZN(new_n566));
  INV_X1    g365(.A(G8gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT101), .Z(new_n571));
  XNOR2_X1  g370(.A(new_n562), .B(KEYINPUT17), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(new_n568), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT102), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n577), .A2(KEYINPUT18), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(KEYINPUT18), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n569), .B2(new_n562), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n575), .B(KEYINPUT13), .Z(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT97), .B(KEYINPUT11), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G169gat), .B(G197gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(KEYINPUT98), .B(KEYINPUT12), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n583), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n583), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT8), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT105), .B(G92gat), .Z(new_n597));
  OAI21_X1  g396(.A(new_n596), .B1(new_n597), .B2(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT106), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G85gat), .A2(G92gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT7), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(G99gat), .B(G106gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n572), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  INV_X1    g406(.A(KEYINPUT107), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT41), .ZN(new_n609));
  NAND2_X1  g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  OAI22_X1  g409(.A1(new_n607), .A2(new_n608), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n605), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n611), .B1(new_n612), .B2(new_n562), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n606), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n608), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n609), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n620), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(G57gat), .B(G64gat), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G71gat), .B(G78gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n568), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n569), .B1(KEYINPUT21), .B2(new_n628), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G127gat), .B(G155gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n303), .ZN(new_n638));
  INV_X1    g437(.A(G211gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n636), .B(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n623), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(G230gat), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n258), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT108), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n605), .B(new_n628), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT10), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n612), .A2(KEYINPUT10), .A3(new_n628), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n648), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n647), .B2(new_n649), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n659), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AND4_X1   g462(.A1(new_n549), .A2(new_n594), .A3(new_n644), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n438), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n372), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT42), .B1(new_n668), .B2(new_n567), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  MUX2_X1   g470(.A(KEYINPUT42), .B(new_n669), .S(new_n671), .Z(G1325gat));
  AOI21_X1  g471(.A(G15gat), .B1(new_n664), .B2(new_n484), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n478), .A2(G15gat), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(new_n664), .B2(new_n674), .ZN(G1326gat));
  INV_X1    g474(.A(new_n279), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n664), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT43), .B(G22gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1327gat));
  NAND3_X1  g478(.A1(new_n594), .A2(new_n643), .A3(new_n663), .ZN(new_n680));
  INV_X1    g479(.A(new_n623), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n547), .A2(new_n548), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(G29gat), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n438), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT45), .Z(new_n687));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n547), .A2(new_n548), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n536), .B1(new_n487), .B2(new_n542), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n537), .A2(new_n486), .A3(new_n364), .A4(new_n539), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n691), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n541), .B(KEYINPUT109), .C1(new_n536), .C2(new_n543), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n440), .A2(new_n478), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n534), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n623), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(new_n688), .ZN(new_n700));
  INV_X1    g499(.A(new_n680), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n690), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT110), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n690), .A2(new_n700), .A3(KEYINPUT110), .A4(new_n701), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n439), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n685), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT111), .ZN(new_n708));
  OR3_X1    g507(.A1(new_n687), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n687), .B2(new_n707), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(G1328gat));
  NOR3_X1   g510(.A1(new_n683), .A2(G36gat), .A3(new_n372), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT46), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n704), .A2(new_n705), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT112), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n667), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G36gat), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(new_n714), .B2(new_n667), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n713), .B1(new_n717), .B2(new_n718), .ZN(G1329gat));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n684), .A2(new_n721), .A3(new_n484), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n721), .B1(new_n714), .B2(new_n478), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI211_X1 g524(.A(KEYINPUT113), .B(new_n721), .C1(new_n714), .C2(new_n478), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n720), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G43gat), .B1(new_n702), .B2(new_n485), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(KEYINPUT47), .A3(new_n722), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1330gat));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n676), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n731), .A2(new_n732), .A3(G50gat), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n279), .B1(new_n704), .B2(new_n705), .ZN(new_n734));
  INV_X1    g533(.A(G50gat), .ZN(new_n735));
  OAI21_X1  g534(.A(KEYINPUT115), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n279), .A2(G50gat), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n683), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n683), .A2(new_n738), .ZN(new_n741));
  AOI21_X1  g540(.A(KEYINPUT117), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n741), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n743), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n733), .A2(new_n736), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G50gat), .B1(new_n702), .B2(new_n279), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n750), .B(KEYINPUT48), .C1(new_n743), .C2(new_n739), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1331gat));
  NOR4_X1   g551(.A1(new_n594), .A2(new_n663), .A3(new_n643), .A4(new_n623), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n698), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n438), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g556(.A1(new_n754), .A2(new_n372), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n755), .A2(new_n763), .A3(new_n484), .ZN(new_n764));
  OAI21_X1  g563(.A(G71gat), .B1(new_n754), .B2(new_n485), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g566(.A1(new_n755), .A2(new_n676), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  INV_X1    g568(.A(new_n643), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n594), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n690), .A2(new_n700), .A3(new_n662), .A4(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n772), .A2(new_n422), .A3(new_n439), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n698), .A2(new_n623), .A3(new_n771), .ZN(new_n774));
  XOR2_X1   g573(.A(new_n774), .B(KEYINPUT51), .Z(new_n775));
  AND2_X1   g574(.A1(new_n775), .A2(new_n662), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n438), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n773), .B1(new_n777), .B2(new_n422), .ZN(G1336gat));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT118), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n372), .A2(G92gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n776), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(KEYINPUT118), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n597), .B1(new_n772), .B2(new_n372), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n783), .B1(new_n782), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(G1337gat));
  XNOR2_X1  g586(.A(KEYINPUT119), .B(G99gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n776), .A2(new_n484), .A3(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n788), .B1(new_n772), .B2(new_n485), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(G1338gat));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  OAI21_X1  g592(.A(G106gat), .B1(new_n772), .B2(new_n279), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT121), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n279), .A2(G106gat), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n776), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n795), .B1(new_n776), .B2(new_n796), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n793), .B(new_n794), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n662), .A2(new_n796), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT120), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n775), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n802), .A2(new_n794), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n799), .B1(new_n793), .B2(new_n803), .ZN(G1339gat));
  NOR4_X1   g603(.A1(new_n594), .A2(new_n643), .A3(new_n662), .A4(new_n623), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n653), .A2(new_n647), .A3(new_n654), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n806), .A2(KEYINPUT54), .A3(new_n655), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n655), .A2(KEYINPUT54), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n808), .A3(new_n659), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n580), .A2(new_n581), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n574), .A2(new_n576), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n588), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n583), .B2(new_n591), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n811), .A2(new_n660), .A3(new_n812), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n770), .B1(new_n817), .B2(new_n623), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n623), .B1(new_n816), .B2(new_n662), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n811), .A2(new_n660), .A3(new_n812), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n592), .A2(new_n593), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n805), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n439), .A3(new_n667), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(new_n542), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(new_n382), .A3(new_n594), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n540), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n821), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1340gat));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n380), .A3(new_n662), .ZN(new_n830));
  OAI21_X1  g629(.A(G120gat), .B1(new_n827), .B2(new_n663), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1341gat));
  AOI21_X1  g631(.A(G127gat), .B1(new_n825), .B2(new_n770), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n827), .A2(new_n375), .A3(new_n643), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n833), .A2(new_n834), .ZN(G1342gat));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n373), .A3(new_n623), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n836), .A2(KEYINPUT56), .ZN(new_n837));
  OAI21_X1  g636(.A(G134gat), .B1(new_n827), .B2(new_n681), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(KEYINPUT56), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(G1343gat));
  NOR2_X1   g639(.A1(new_n667), .A2(new_n439), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n485), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n823), .A2(new_n279), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n225), .A3(new_n594), .ZN(new_n844));
  NAND2_X1  g643(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n823), .A2(new_n279), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n823), .B2(new_n279), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n842), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n851), .A2(new_n594), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n846), .B1(new_n853), .B2(G141gat), .ZN(new_n854));
  NOR2_X1   g653(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1344gat));
  OAI211_X1 g655(.A(new_n843), .B(new_n662), .C1(new_n244), .C2(new_n243), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT123), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n663), .B(new_n842), .C1(new_n848), .C2(new_n850), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n858), .B(KEYINPUT59), .C1(new_n859), .C2(new_n227), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n851), .A2(new_n662), .A3(new_n852), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n243), .A2(new_n244), .A3(KEYINPUT59), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(G148gat), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n858), .B1(new_n865), .B2(KEYINPUT59), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n857), .B1(new_n864), .B2(new_n866), .ZN(G1345gat));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n868), .A2(new_n240), .A3(new_n643), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n843), .A2(new_n770), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n240), .B2(new_n870), .ZN(G1346gat));
  OAI21_X1  g670(.A(G162gat), .B1(new_n868), .B2(new_n681), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n843), .A2(new_n241), .A3(new_n623), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1347gat));
  NOR3_X1   g673(.A1(new_n823), .A2(new_n438), .A3(new_n372), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n542), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n298), .A3(new_n594), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n875), .A2(new_n540), .ZN(new_n878));
  OAI21_X1  g677(.A(G169gat), .B1(new_n878), .B2(new_n821), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g679(.A(new_n880), .B(KEYINPUT124), .Z(G1348gat));
  NAND2_X1  g680(.A1(new_n876), .A2(new_n662), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(KEYINPUT125), .A3(new_n299), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT125), .B1(new_n882), .B2(new_n299), .ZN(new_n884));
  NOR3_X1   g683(.A1(new_n878), .A2(new_n299), .A3(new_n663), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1349gat));
  NAND3_X1  g685(.A1(new_n876), .A2(new_n282), .A3(new_n770), .ZN(new_n887));
  OAI21_X1  g686(.A(G183gat), .B1(new_n878), .B2(new_n643), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n889), .B(new_n890), .Z(G1350gat));
  NAND3_X1  g690(.A1(new_n876), .A2(new_n283), .A3(new_n623), .ZN(new_n892));
  OAI21_X1  g691(.A(G190gat), .B1(new_n878), .B2(new_n681), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(KEYINPUT61), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1351gat));
  NOR3_X1   g695(.A1(new_n478), .A2(new_n372), .A3(new_n438), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT127), .Z(new_n898));
  NAND2_X1  g697(.A1(new_n851), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(G197gat), .B1(new_n899), .B2(new_n821), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n847), .A2(new_n897), .ZN(new_n901));
  INV_X1    g700(.A(G197gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n594), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(G1352gat));
  INV_X1    g703(.A(G204gat), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n905), .A3(new_n662), .ZN(new_n906));
  XOR2_X1   g705(.A(new_n906), .B(KEYINPUT62), .Z(new_n907));
  OAI21_X1  g706(.A(G204gat), .B1(new_n899), .B2(new_n663), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(G1353gat));
  NAND3_X1  g708(.A1(new_n901), .A2(new_n639), .A3(new_n770), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n851), .A2(new_n770), .A3(new_n898), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n911), .B2(G211gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  INV_X1    g713(.A(G218gat), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n915), .A3(new_n681), .ZN(new_n916));
  AOI21_X1  g715(.A(G218gat), .B1(new_n901), .B2(new_n623), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1355gat));
endmodule


