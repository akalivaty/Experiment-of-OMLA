

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U549 ( .A(n725), .ZN(n700) );
  BUF_X1 U550 ( .A(n604), .Z(n605) );
  NAND2_X1 U551 ( .A1(n762), .A2(n764), .ZN(n725) );
  XOR2_X1 U552 ( .A(n760), .B(KEYINPUT97), .Z(n517) );
  NOR2_X1 U553 ( .A1(n682), .A2(G168), .ZN(n683) );
  INV_X1 U554 ( .A(KEYINPUT94), .ZN(n717) );
  NOR2_X1 U555 ( .A1(G651), .A2(G543), .ZN(n623) );
  NAND2_X1 U556 ( .A1(n623), .A2(G89), .ZN(n518) );
  XNOR2_X1 U557 ( .A(n518), .B(KEYINPUT4), .ZN(n520) );
  XOR2_X1 U558 ( .A(KEYINPUT0), .B(G543), .Z(n635) );
  INV_X1 U559 ( .A(G651), .ZN(n522) );
  NOR2_X1 U560 ( .A1(n635), .A2(n522), .ZN(n626) );
  NAND2_X1 U561 ( .A1(G76), .A2(n626), .ZN(n519) );
  NAND2_X1 U562 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U563 ( .A(n521), .B(KEYINPUT5), .ZN(n529) );
  XNOR2_X1 U564 ( .A(KEYINPUT71), .B(KEYINPUT6), .ZN(n527) );
  NOR2_X1 U565 ( .A1(G543), .A2(n522), .ZN(n523) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n523), .Z(n639) );
  NAND2_X1 U567 ( .A1(G63), .A2(n639), .ZN(n525) );
  NOR2_X1 U568 ( .A1(G651), .A2(n635), .ZN(n633) );
  NAND2_X1 U569 ( .A1(G51), .A2(n633), .ZN(n524) );
  NAND2_X1 U570 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U571 ( .A(n527), .B(n526), .ZN(n528) );
  NAND2_X1 U572 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U573 ( .A(KEYINPUT7), .B(n530), .ZN(G168) );
  XNOR2_X1 U574 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n532) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XNOR2_X2 U576 ( .A(n532), .B(n531), .ZN(n895) );
  NAND2_X1 U577 ( .A1(n895), .A2(G137), .ZN(n542) );
  INV_X1 U578 ( .A(G2104), .ZN(n537) );
  NAND2_X1 U579 ( .A1(n537), .A2(G2105), .ZN(n533) );
  XNOR2_X1 U580 ( .A(n533), .B(KEYINPUT65), .ZN(n670) );
  NAND2_X1 U581 ( .A1(G125), .A2(n670), .ZN(n536) );
  NAND2_X1 U582 ( .A1(G2105), .A2(G2104), .ZN(n534) );
  XOR2_X1 U583 ( .A(KEYINPUT66), .B(n534), .Z(n671) );
  NAND2_X1 U584 ( .A1(G113), .A2(n671), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n540) );
  NOR2_X1 U586 ( .A1(G2105), .A2(n537), .ZN(n604) );
  NAND2_X1 U587 ( .A1(G101), .A2(n604), .ZN(n538) );
  XNOR2_X1 U588 ( .A(KEYINPUT23), .B(n538), .ZN(n539) );
  NOR2_X1 U589 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U590 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X2 U591 ( .A(KEYINPUT64), .B(n543), .Z(G160) );
  NAND2_X1 U592 ( .A1(G72), .A2(n626), .ZN(n545) );
  NAND2_X1 U593 ( .A1(G85), .A2(n623), .ZN(n544) );
  NAND2_X1 U594 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U595 ( .A1(G60), .A2(n639), .ZN(n547) );
  NAND2_X1 U596 ( .A1(G47), .A2(n633), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n547), .A2(n546), .ZN(n548) );
  OR2_X1 U598 ( .A1(n549), .A2(n548), .ZN(G290) );
  AND2_X1 U599 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U600 ( .A(G57), .ZN(G237) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  NAND2_X1 U603 ( .A1(G64), .A2(n639), .ZN(n551) );
  NAND2_X1 U604 ( .A1(G52), .A2(n633), .ZN(n550) );
  NAND2_X1 U605 ( .A1(n551), .A2(n550), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G77), .A2(n626), .ZN(n553) );
  NAND2_X1 U607 ( .A1(G90), .A2(n623), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U609 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  NOR2_X1 U610 ( .A1(n556), .A2(n555), .ZN(G171) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G88), .A2(n623), .ZN(n557) );
  XNOR2_X1 U613 ( .A(n557), .B(KEYINPUT78), .ZN(n564) );
  NAND2_X1 U614 ( .A1(G62), .A2(n639), .ZN(n559) );
  NAND2_X1 U615 ( .A1(G50), .A2(n633), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n559), .A2(n558), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G75), .A2(n626), .ZN(n560) );
  XNOR2_X1 U618 ( .A(KEYINPUT79), .B(n560), .ZN(n561) );
  NOR2_X1 U619 ( .A1(n562), .A2(n561), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n564), .A2(n563), .ZN(G303) );
  INV_X1 U621 ( .A(G303), .ZN(G166) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U623 ( .A(n565), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U624 ( .A(G223), .B(KEYINPUT68), .Z(n815) );
  NAND2_X1 U625 ( .A1(n815), .A2(G567), .ZN(n566) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  XNOR2_X1 U627 ( .A(KEYINPUT69), .B(KEYINPUT13), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n623), .A2(G81), .ZN(n567) );
  XNOR2_X1 U629 ( .A(n567), .B(KEYINPUT12), .ZN(n569) );
  NAND2_X1 U630 ( .A1(G68), .A2(n626), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U632 ( .A(n571), .B(n570), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n639), .A2(G56), .ZN(n572) );
  XOR2_X1 U634 ( .A(KEYINPUT14), .B(n572), .Z(n573) );
  NOR2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U636 ( .A1(n633), .A2(G43), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n1005) );
  INV_X1 U638 ( .A(G860), .ZN(n596) );
  OR2_X1 U639 ( .A1(n1005), .A2(n596), .ZN(G153) );
  INV_X1 U640 ( .A(G171), .ZN(G301) );
  NAND2_X1 U641 ( .A1(G868), .A2(G301), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(KEYINPUT70), .ZN(n586) );
  NAND2_X1 U643 ( .A1(G79), .A2(n626), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G92), .A2(n623), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G66), .A2(n639), .ZN(n581) );
  NAND2_X1 U647 ( .A1(G54), .A2(n633), .ZN(n580) );
  NAND2_X1 U648 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U649 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U650 ( .A(KEYINPUT15), .B(n584), .Z(n1004) );
  OR2_X1 U651 ( .A1(G868), .A2(n1004), .ZN(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G65), .A2(n639), .ZN(n588) );
  NAND2_X1 U654 ( .A1(G53), .A2(n633), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G78), .A2(n626), .ZN(n590) );
  NAND2_X1 U657 ( .A1(G91), .A2(n623), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U659 ( .A1(n592), .A2(n591), .ZN(n993) );
  INV_X1 U660 ( .A(n993), .ZN(G299) );
  XOR2_X1 U661 ( .A(G868), .B(KEYINPUT72), .Z(n593) );
  NOR2_X1 U662 ( .A1(G286), .A2(n593), .ZN(n595) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n597), .A2(n1004), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT73), .ZN(n599) );
  XOR2_X1 U668 ( .A(KEYINPUT16), .B(n599), .Z(G148) );
  NOR2_X1 U669 ( .A1(G868), .A2(n1005), .ZN(n602) );
  NAND2_X1 U670 ( .A1(n1004), .A2(G868), .ZN(n600) );
  NOR2_X1 U671 ( .A1(G559), .A2(n600), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(G282) );
  BUF_X1 U673 ( .A(n670), .Z(n891) );
  NAND2_X1 U674 ( .A1(G123), .A2(n891), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n603), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U676 ( .A1(G99), .A2(n605), .ZN(n607) );
  BUF_X1 U677 ( .A(n671), .Z(n892) );
  NAND2_X1 U678 ( .A1(G111), .A2(n892), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U680 ( .A1(n895), .A2(G135), .ZN(n608) );
  XOR2_X1 U681 ( .A(KEYINPUT74), .B(n608), .Z(n609) );
  NOR2_X1 U682 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n922) );
  XOR2_X1 U684 ( .A(n922), .B(G2096), .Z(n614) );
  XNOR2_X1 U685 ( .A(G2100), .B(KEYINPUT75), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n1004), .A2(G559), .ZN(n651) );
  XNOR2_X1 U688 ( .A(n1005), .B(n651), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n615), .A2(G860), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G67), .A2(n639), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G55), .A2(n633), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G80), .A2(n626), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G93), .A2(n623), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n621), .A2(n620), .ZN(n649) );
  XNOR2_X1 U697 ( .A(n622), .B(n649), .ZN(G145) );
  NAND2_X1 U698 ( .A1(G86), .A2(n623), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G48), .A2(n633), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT2), .B(KEYINPUT77), .Z(n628) );
  NAND2_X1 U702 ( .A1(n626), .A2(G73), .ZN(n627) );
  XOR2_X1 U703 ( .A(n628), .B(n627), .Z(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n639), .A2(G61), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U707 ( .A1(G49), .A2(n633), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT76), .ZN(n641) );
  NAND2_X1 U709 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(G288) );
  NOR2_X1 U714 ( .A1(G868), .A2(n649), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(KEYINPUT81), .ZN(n654) );
  XOR2_X1 U716 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n643) );
  XNOR2_X1 U717 ( .A(G290), .B(n643), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n644), .B(G305), .ZN(n645) );
  XNOR2_X1 U719 ( .A(n645), .B(n1005), .ZN(n646) );
  XNOR2_X1 U720 ( .A(G166), .B(n646), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n647), .B(G288), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n993), .B(n648), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(n649), .ZN(n859) );
  XOR2_X1 U724 ( .A(n859), .B(n651), .Z(n652) );
  NAND2_X1 U725 ( .A1(G868), .A2(n652), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U727 ( .A1(G2084), .A2(G2078), .ZN(n655) );
  XOR2_X1 U728 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U729 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U730 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U732 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U733 ( .A1(G220), .A2(G219), .ZN(n659) );
  XOR2_X1 U734 ( .A(KEYINPUT22), .B(n659), .Z(n660) );
  NOR2_X1 U735 ( .A1(G218), .A2(n660), .ZN(n661) );
  NAND2_X1 U736 ( .A1(G96), .A2(n661), .ZN(n820) );
  NAND2_X1 U737 ( .A1(n820), .A2(G2106), .ZN(n665) );
  NAND2_X1 U738 ( .A1(G69), .A2(G120), .ZN(n662) );
  NOR2_X1 U739 ( .A1(G237), .A2(n662), .ZN(n663) );
  NAND2_X1 U740 ( .A1(G108), .A2(n663), .ZN(n821) );
  NAND2_X1 U741 ( .A1(n821), .A2(G567), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n915) );
  NAND2_X1 U743 ( .A1(G483), .A2(G661), .ZN(n666) );
  NOR2_X1 U744 ( .A1(n915), .A2(n666), .ZN(n819) );
  NAND2_X1 U745 ( .A1(n819), .A2(G36), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT82), .B(n667), .ZN(G176) );
  NAND2_X1 U747 ( .A1(G102), .A2(n605), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G138), .A2(n895), .ZN(n668) );
  NAND2_X1 U749 ( .A1(n669), .A2(n668), .ZN(n675) );
  NAND2_X1 U750 ( .A1(G126), .A2(n670), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G114), .A2(n671), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U753 ( .A1(n675), .A2(n674), .ZN(G164) );
  NOR2_X1 U754 ( .A1(G1981), .A2(G305), .ZN(n676) );
  XNOR2_X1 U755 ( .A(KEYINPUT24), .B(n676), .ZN(n679) );
  NAND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n677) );
  XNOR2_X1 U757 ( .A(n677), .B(KEYINPUT83), .ZN(n762) );
  NOR2_X1 U758 ( .A1(G164), .A2(G1384), .ZN(n764) );
  NAND2_X1 U759 ( .A1(G8), .A2(n725), .ZN(n678) );
  XNOR2_X2 U760 ( .A(n678), .B(KEYINPUT90), .ZN(n745) );
  INV_X1 U761 ( .A(n745), .ZN(n747) );
  NAND2_X1 U762 ( .A1(n679), .A2(n747), .ZN(n741) );
  NOR2_X1 U763 ( .A1(n745), .A2(G1966), .ZN(n719) );
  NOR2_X1 U764 ( .A1(G2084), .A2(n725), .ZN(n720) );
  NOR2_X1 U765 ( .A1(n719), .A2(n720), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n680), .A2(G8), .ZN(n681) );
  XNOR2_X1 U767 ( .A(KEYINPUT30), .B(n681), .ZN(n682) );
  XNOR2_X1 U768 ( .A(n683), .B(KEYINPUT93), .ZN(n687) );
  XOR2_X1 U769 ( .A(G2078), .B(KEYINPUT25), .Z(n942) );
  NOR2_X1 U770 ( .A1(n942), .A2(n725), .ZN(n685) );
  NOR2_X1 U771 ( .A1(n700), .A2(G1961), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n685), .A2(n684), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n689), .A2(G301), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U775 ( .A(n688), .B(KEYINPUT31), .ZN(n716) );
  OR2_X1 U776 ( .A1(n689), .A2(G301), .ZN(n714) );
  NAND2_X1 U777 ( .A1(n700), .A2(G2072), .ZN(n690) );
  XNOR2_X1 U778 ( .A(n690), .B(KEYINPUT27), .ZN(n692) );
  XNOR2_X1 U779 ( .A(KEYINPUT91), .B(G1956), .ZN(n970) );
  NOR2_X1 U780 ( .A1(n970), .A2(n700), .ZN(n691) );
  NOR2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n694) );
  NOR2_X1 U782 ( .A1(n993), .A2(n694), .ZN(n693) );
  XOR2_X1 U783 ( .A(n693), .B(KEYINPUT28), .Z(n711) );
  NAND2_X1 U784 ( .A1(n993), .A2(n694), .ZN(n709) );
  AND2_X1 U785 ( .A1(n700), .A2(G1996), .ZN(n695) );
  XOR2_X1 U786 ( .A(n695), .B(KEYINPUT26), .Z(n698) );
  AND2_X1 U787 ( .A1(n725), .A2(G1341), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n696), .A2(n1005), .ZN(n697) );
  AND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n1004), .A2(n705), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n725), .A2(G1348), .ZN(n699) );
  XNOR2_X1 U792 ( .A(n699), .B(KEYINPUT92), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n700), .A2(G2067), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U795 ( .A1(n704), .A2(n703), .ZN(n707) );
  OR2_X1 U796 ( .A1(n1004), .A2(n705), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U798 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U800 ( .A(n712), .B(KEYINPUT29), .Z(n713) );
  NAND2_X1 U801 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n724) );
  XNOR2_X1 U803 ( .A(n724), .B(n717), .ZN(n718) );
  NOR2_X1 U804 ( .A1(n719), .A2(n718), .ZN(n722) );
  NAND2_X1 U805 ( .A1(G8), .A2(n720), .ZN(n721) );
  NAND2_X1 U806 ( .A1(n722), .A2(n721), .ZN(n736) );
  AND2_X1 U807 ( .A1(G286), .A2(G8), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n724), .A2(n723), .ZN(n732) );
  INV_X1 U809 ( .A(G8), .ZN(n730) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n725), .ZN(n727) );
  NOR2_X1 U811 ( .A1(n745), .A2(G1971), .ZN(n726) );
  NOR2_X1 U812 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U813 ( .A1(n728), .A2(G303), .ZN(n729) );
  OR2_X1 U814 ( .A1(n730), .A2(n729), .ZN(n731) );
  AND2_X1 U815 ( .A1(n732), .A2(n731), .ZN(n734) );
  XOR2_X1 U816 ( .A(KEYINPUT32), .B(KEYINPUT95), .Z(n733) );
  XNOR2_X1 U817 ( .A(n734), .B(n733), .ZN(n735) );
  NAND2_X1 U818 ( .A1(n736), .A2(n735), .ZN(n744) );
  NOR2_X1 U819 ( .A1(G2090), .A2(G303), .ZN(n737) );
  NAND2_X1 U820 ( .A1(G8), .A2(n737), .ZN(n738) );
  NAND2_X1 U821 ( .A1(n744), .A2(n738), .ZN(n739) );
  NAND2_X1 U822 ( .A1(n739), .A2(n745), .ZN(n740) );
  NAND2_X1 U823 ( .A1(n741), .A2(n740), .ZN(n761) );
  INV_X1 U824 ( .A(G1971), .ZN(n963) );
  AND2_X1 U825 ( .A1(G166), .A2(n963), .ZN(n742) );
  NOR2_X1 U826 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NOR2_X1 U827 ( .A1(n742), .A2(n990), .ZN(n743) );
  AND2_X1 U828 ( .A1(n744), .A2(n743), .ZN(n746) );
  NOR2_X1 U829 ( .A1(n746), .A2(n745), .ZN(n753) );
  NAND2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n994) );
  INV_X1 U831 ( .A(KEYINPUT33), .ZN(n755) );
  NAND2_X1 U832 ( .A1(n990), .A2(n747), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n755), .A2(n748), .ZN(n749) );
  XOR2_X1 U834 ( .A(n749), .B(KEYINPUT96), .Z(n754) );
  AND2_X1 U835 ( .A1(n994), .A2(n754), .ZN(n751) );
  XNOR2_X1 U836 ( .A(G1981), .B(G305), .ZN(n1002) );
  INV_X1 U837 ( .A(n1002), .ZN(n750) );
  AND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n759) );
  INV_X1 U840 ( .A(n754), .ZN(n756) );
  OR2_X1 U841 ( .A1(n756), .A2(n755), .ZN(n757) );
  OR2_X1 U842 ( .A1(n1002), .A2(n757), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U844 ( .A1(n761), .A2(n517), .ZN(n788) );
  XNOR2_X1 U845 ( .A(G1986), .B(G290), .ZN(n997) );
  INV_X1 U846 ( .A(n762), .ZN(n763) );
  NOR2_X1 U847 ( .A1(n764), .A2(n763), .ZN(n810) );
  NAND2_X1 U848 ( .A1(n997), .A2(n810), .ZN(n765) );
  XNOR2_X1 U849 ( .A(n765), .B(KEYINPUT84), .ZN(n786) );
  NAND2_X1 U850 ( .A1(G95), .A2(n605), .ZN(n767) );
  NAND2_X1 U851 ( .A1(G131), .A2(n895), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U853 ( .A(KEYINPUT86), .B(n768), .Z(n772) );
  NAND2_X1 U854 ( .A1(n892), .A2(G107), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G119), .A2(n891), .ZN(n769) );
  AND2_X1 U856 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n870) );
  NAND2_X1 U858 ( .A1(n870), .A2(G1991), .ZN(n782) );
  NAND2_X1 U859 ( .A1(G129), .A2(n891), .ZN(n774) );
  NAND2_X1 U860 ( .A1(G117), .A2(n892), .ZN(n773) );
  NAND2_X1 U861 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U862 ( .A1(n605), .A2(G105), .ZN(n775) );
  XOR2_X1 U863 ( .A(KEYINPUT38), .B(n775), .Z(n776) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U865 ( .A(KEYINPUT87), .B(n778), .Z(n780) );
  NAND2_X1 U866 ( .A1(n895), .A2(G141), .ZN(n779) );
  NAND2_X1 U867 ( .A1(n780), .A2(n779), .ZN(n873) );
  NAND2_X1 U868 ( .A1(G1996), .A2(n873), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT88), .ZN(n918) );
  NAND2_X1 U871 ( .A1(n918), .A2(n810), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT89), .ZN(n803) );
  INV_X1 U873 ( .A(n803), .ZN(n785) );
  NAND2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U875 ( .A1(n788), .A2(n787), .ZN(n799) );
  NAND2_X1 U876 ( .A1(n895), .A2(G140), .ZN(n789) );
  XOR2_X1 U877 ( .A(KEYINPUT85), .B(n789), .Z(n791) );
  NAND2_X1 U878 ( .A1(n605), .A2(G104), .ZN(n790) );
  NAND2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U880 ( .A(KEYINPUT34), .B(n792), .ZN(n797) );
  NAND2_X1 U881 ( .A1(G128), .A2(n891), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G116), .A2(n892), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  XOR2_X1 U884 ( .A(KEYINPUT35), .B(n795), .Z(n796) );
  NOR2_X1 U885 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U886 ( .A(KEYINPUT36), .B(n798), .ZN(n871) );
  XNOR2_X1 U887 ( .A(G2067), .B(KEYINPUT37), .ZN(n800) );
  NOR2_X1 U888 ( .A1(n871), .A2(n800), .ZN(n937) );
  NAND2_X1 U889 ( .A1(n937), .A2(n810), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n799), .A2(n806), .ZN(n813) );
  NAND2_X1 U891 ( .A1(n871), .A2(n800), .ZN(n916) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n873), .ZN(n920) );
  NOR2_X1 U893 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U894 ( .A1(G1991), .A2(n870), .ZN(n925) );
  NOR2_X1 U895 ( .A1(n801), .A2(n925), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U897 ( .A1(n920), .A2(n804), .ZN(n805) );
  XNOR2_X1 U898 ( .A(KEYINPUT39), .B(n805), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n807), .A2(n806), .ZN(n808) );
  NAND2_X1 U900 ( .A1(n916), .A2(n808), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U902 ( .A(n811), .B(KEYINPUT98), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U904 ( .A(n814), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n815), .ZN(G217) );
  NAND2_X1 U906 ( .A1(G15), .A2(G2), .ZN(n816) );
  XOR2_X1 U907 ( .A(KEYINPUT102), .B(n816), .Z(n817) );
  NAND2_X1 U908 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U910 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U912 ( .A(G120), .ZN(G236) );
  INV_X1 U913 ( .A(G96), .ZN(G221) );
  INV_X1 U914 ( .A(G69), .ZN(G235) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U917 ( .A(G2443), .B(G2438), .ZN(n831) );
  XOR2_X1 U918 ( .A(G2454), .B(G2430), .Z(n823) );
  XNOR2_X1 U919 ( .A(G2446), .B(KEYINPUT99), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n827) );
  XOR2_X1 U921 ( .A(G2451), .B(G2427), .Z(n825) );
  XNOR2_X1 U922 ( .A(G1341), .B(G1348), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n826) );
  XOR2_X1 U924 ( .A(n827), .B(n826), .Z(n829) );
  XNOR2_X1 U925 ( .A(G2435), .B(KEYINPUT100), .ZN(n828) );
  XNOR2_X1 U926 ( .A(n829), .B(n828), .ZN(n830) );
  XNOR2_X1 U927 ( .A(n831), .B(n830), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n832), .A2(G14), .ZN(n833) );
  XNOR2_X1 U929 ( .A(KEYINPUT101), .B(n833), .ZN(G401) );
  XOR2_X1 U930 ( .A(G2096), .B(G2090), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2072), .B(G2067), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n845) );
  XOR2_X1 U933 ( .A(KEYINPUT106), .B(G2678), .Z(n837) );
  XNOR2_X1 U934 ( .A(KEYINPUT104), .B(KEYINPUT103), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U936 ( .A(G2100), .B(KEYINPUT43), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U940 ( .A(G2084), .B(G2078), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(n845), .B(n844), .Z(G227) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G1986), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1971), .B(G1976), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n848), .B(KEYINPUT108), .Z(n850) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U949 ( .A(G1956), .B(G1961), .Z(n852) );
  XNOR2_X1 U950 ( .A(G1981), .B(G1966), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2474), .B(KEYINPUT107), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U955 ( .A(KEYINPUT119), .B(G286), .Z(n858) );
  XNOR2_X1 U956 ( .A(G171), .B(n1004), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  NOR2_X1 U959 ( .A1(G37), .A2(n861), .ZN(G397) );
  NAND2_X1 U960 ( .A1(G100), .A2(n605), .ZN(n863) );
  NAND2_X1 U961 ( .A1(G136), .A2(n895), .ZN(n862) );
  NAND2_X1 U962 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U963 ( .A1(G124), .A2(n891), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n864), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U965 ( .A1(n892), .A2(G112), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT109), .B(n865), .Z(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(G162) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U971 ( .A(n922), .B(n874), .ZN(n884) );
  NAND2_X1 U972 ( .A1(G103), .A2(n605), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G139), .A2(n895), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n881) );
  NAND2_X1 U975 ( .A1(G127), .A2(n891), .ZN(n878) );
  NAND2_X1 U976 ( .A1(G115), .A2(n892), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT112), .B(n882), .Z(n928) );
  XNOR2_X1 U981 ( .A(n928), .B(G162), .ZN(n883) );
  XNOR2_X1 U982 ( .A(n884), .B(n883), .ZN(n907) );
  XOR2_X1 U983 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n886) );
  XNOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT116), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n890) );
  XOR2_X1 U986 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n888) );
  XNOR2_X1 U987 ( .A(KEYINPUT113), .B(KEYINPUT111), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U989 ( .A(n890), .B(n889), .Z(n904) );
  NAND2_X1 U990 ( .A1(G130), .A2(n891), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G118), .A2(n892), .ZN(n893) );
  NAND2_X1 U992 ( .A1(n894), .A2(n893), .ZN(n901) );
  NAND2_X1 U993 ( .A1(n895), .A2(G142), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n896), .B(KEYINPUT110), .ZN(n898) );
  NAND2_X1 U995 ( .A1(G106), .A2(n605), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT45), .B(n899), .Z(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(G164), .B(n902), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(G160), .B(n905), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1004 ( .A(KEYINPUT118), .B(n909), .ZN(G395) );
  OR2_X1 U1005 ( .A1(n915), .A2(G401), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G397), .A2(G395), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1011 ( .A(G225), .ZN(G308) );
  INV_X1 U1012 ( .A(n915), .ZN(G319) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  INV_X1 U1014 ( .A(n916), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n935) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n921), .Z(n927) );
  XNOR2_X1 U1019 ( .A(G160), .B(G2084), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n930) );
  XNOR2_X1 U1024 ( .A(G2072), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1026 ( .A(KEYINPUT50), .B(n931), .Z(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1028 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1031 ( .A(KEYINPUT55), .ZN(n959) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n959), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1034 ( .A(G2090), .B(G35), .ZN(n954) );
  XOR2_X1 U1035 ( .A(G1991), .B(G25), .Z(n941) );
  NAND2_X1 U1036 ( .A1(n941), .A2(G28), .ZN(n951) );
  XNOR2_X1 U1037 ( .A(n942), .B(G27), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G32), .B(G1996), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(KEYINPUT120), .B(n945), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(G2072), .B(G33), .ZN(n947) );
  XNOR2_X1 U1042 ( .A(G2067), .B(G26), .ZN(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(KEYINPUT53), .B(n952), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1048 ( .A(G2084), .B(KEYINPUT54), .Z(n955) );
  XNOR2_X1 U1049 ( .A(G34), .B(n955), .ZN(n956) );
  NAND2_X1 U1050 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(n959), .B(n958), .ZN(n961) );
  INV_X1 U1052 ( .A(G29), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1054 ( .A1(G11), .A2(n962), .ZN(n1020) );
  XOR2_X1 U1055 ( .A(KEYINPUT124), .B(G16), .Z(n989) );
  XNOR2_X1 U1056 ( .A(G22), .B(n963), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G1976), .B(G23), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(G1986), .B(G24), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n968) );
  XNOR2_X1 U1062 ( .A(n969), .B(n968), .ZN(n985) );
  XNOR2_X1 U1063 ( .A(G20), .B(n970), .ZN(n974) );
  XNOR2_X1 U1064 ( .A(G1981), .B(G6), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(G19), .B(G1341), .ZN(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1068 ( .A(KEYINPUT59), .B(G1348), .Z(n975) );
  XNOR2_X1 U1069 ( .A(G4), .B(n975), .ZN(n976) );
  NOR2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(KEYINPUT60), .B(n978), .ZN(n982) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G21), .ZN(n980) );
  XNOR2_X1 U1073 ( .A(G1961), .B(G5), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1076 ( .A(KEYINPUT125), .B(n983), .ZN(n984) );
  NAND2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(n986), .B(KEYINPUT127), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT61), .B(n987), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n1018) );
  XOR2_X1 U1081 ( .A(n990), .B(KEYINPUT121), .Z(n992) );
  XOR2_X1 U1082 ( .A(G166), .B(G1971), .Z(n991) );
  NOR2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(n993), .B(G1956), .ZN(n995) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(KEYINPUT122), .B(n1000), .ZN(n1013) );
  XOR2_X1 U1089 ( .A(G168), .B(G1966), .Z(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(KEYINPUT57), .B(n1003), .Z(n1011) );
  XNOR2_X1 U1092 ( .A(n1004), .B(G1348), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(G1341), .B(n1005), .Z(n1006) );
  NAND2_X1 U1094 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G1961), .B(G301), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1098 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1099 ( .A(n1014), .B(KEYINPUT123), .ZN(n1016) );
  XNOR2_X1 U1100 ( .A(G16), .B(KEYINPUT56), .ZN(n1015) );
  NAND2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

