//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT67), .Z(G261));
  AND2_X1   g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n457), .A2(new_n458), .ZN(new_n460));
  AOI211_X1 g035(.A(new_n459), .B(new_n460), .C1(G567), .C2(new_n454), .ZN(G319));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(KEYINPUT69), .B(G2105), .C1(new_n467), .C2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  AOI21_X1  g053(.A(KEYINPUT69), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n474), .A2(new_n479), .ZN(G160));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(new_n465), .B2(new_n466), .ZN(new_n482));
  MUX2_X1   g057(.A(G100), .B(G112), .S(G2105), .Z(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n482), .B1(new_n483), .B2(G2104), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n471), .A2(G136), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT70), .ZN(G162));
  NAND2_X1  g062(.A1(G114), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G102), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2104), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n481), .C1(new_n475), .C2(new_n476), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  XNOR2_X1  g070(.A(KEYINPUT3), .B(G2104), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n496), .A2(new_n497), .A3(G138), .A4(new_n481), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n495), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT72), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(new_n501), .A3(G543), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  INV_X1    g086(.A(G50), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G543), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n505), .A2(G62), .A3(new_n506), .A4(new_n508), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  XOR2_X1   g092(.A(new_n517), .B(KEYINPUT73), .Z(new_n518));
  AOI21_X1  g093(.A(new_n515), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n514), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  INV_X1    g097(.A(G51), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n522), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  AND4_X1   g099(.A1(new_n505), .A2(new_n506), .A3(new_n508), .A4(new_n509), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n524), .B1(G89), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n502), .A2(new_n504), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n506), .A2(new_n508), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n505), .A2(KEYINPUT74), .A3(new_n506), .A4(new_n508), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(G63), .A2(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n526), .B1(new_n532), .B2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND3_X1  g110(.A1(new_n530), .A2(G64), .A3(new_n531), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n515), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n510), .A2(new_n539), .B1(new_n540), .B2(new_n513), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  INV_X1    g117(.A(new_n513), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n530), .A2(G56), .A3(new_n531), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g122(.A(KEYINPUT75), .B(new_n544), .C1(new_n547), .C2(new_n515), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT75), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n515), .B1(new_n545), .B2(new_n546), .ZN(new_n550));
  INV_X1    g125(.A(new_n544), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND4_X1  g135(.A1(new_n505), .A2(G65), .A3(new_n506), .A4(new_n508), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n525), .A2(new_n567), .A3(G91), .ZN(new_n568));
  INV_X1    g143(.A(G91), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT76), .B1(new_n510), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n564), .A2(new_n566), .A3(new_n568), .A4(new_n570), .ZN(G299));
  INV_X1    g146(.A(G171), .ZN(G301));
  INV_X1    g147(.A(G166), .ZN(G303));
  AOI22_X1  g148(.A1(new_n525), .A2(G87), .B1(G49), .B2(new_n543), .ZN(new_n574));
  AOI21_X1  g149(.A(G74), .B1(new_n530), .B2(new_n531), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n515), .ZN(G288));
  NAND2_X1  g151(.A1(new_n525), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n543), .A2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n505), .A2(G61), .A3(new_n506), .A4(new_n508), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  XOR2_X1   g157(.A(new_n582), .B(KEYINPUT77), .Z(new_n583));
  AOI21_X1  g158(.A(new_n515), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI211_X1 g162(.A(new_n586), .B(new_n515), .C1(new_n581), .C2(new_n583), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n580), .A2(new_n587), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(G72), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G60), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n532), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G54), .B2(new_n543), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n525), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n510), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g184(.A(new_n608), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  XNOR2_X1  g186(.A(G299), .B(KEYINPUT79), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G297));
  OAI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G280));
  AND2_X1   g189(.A1(new_n601), .A2(new_n606), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G860), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT80), .Z(G148));
  NAND2_X1  g193(.A1(new_n615), .A2(new_n616), .ZN(new_n619));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g196(.A(new_n621), .B1(new_n554), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g198(.A(new_n471), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT12), .B1(new_n624), .B2(new_n464), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n471), .A2(new_n626), .A3(G2104), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT81), .B(G2100), .Z(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  MUX2_X1   g207(.A(G99), .B(G111), .S(G2105), .Z(new_n633));
  AOI22_X1  g208(.A1(G123), .A2(new_n482), .B1(new_n633), .B2(G2104), .ZN(new_n634));
  INV_X1    g209(.A(G135), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n624), .ZN(new_n636));
  INV_X1    g211(.A(G2096), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G1341), .B(G1348), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT14), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT15), .B(G2435), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2438), .ZN(new_n648));
  XOR2_X1   g223(.A(G2427), .B(G2430), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT82), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n648), .B2(new_n650), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n645), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(G14), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  INV_X1    g236(.A(new_n657), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(new_n659), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n665), .B1(new_n662), .B2(new_n663), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n657), .A2(new_n659), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n658), .B1(new_n667), .B2(KEYINPUT17), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n661), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(new_n637), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(G2100), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT84), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n683));
  NOR2_X1   g258(.A1(new_n678), .A2(new_n681), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n682), .A2(new_n683), .B1(new_n684), .B2(new_n674), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n680), .B(new_n685), .C1(new_n682), .C2(new_n683), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n688), .B(new_n691), .Z(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  MUX2_X1   g268(.A(G6), .B(G305), .S(G16), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT90), .B(G1971), .Z(new_n701));
  XOR2_X1   g276(.A(new_n700), .B(new_n701), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n697), .A2(G23), .ZN(new_n703));
  INV_X1    g278(.A(G288), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n697), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT33), .B(G1976), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n705), .B(new_n706), .Z(new_n707));
  NOR3_X1   g282(.A1(new_n696), .A2(new_n702), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G290), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT86), .B(G1986), .Z(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT87), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G95), .B(G107), .S(G2105), .Z(new_n718));
  AOI22_X1  g293(.A1(G119), .A2(new_n482), .B1(new_n718), .B2(G2104), .ZN(new_n719));
  INV_X1    g294(.A(G131), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n624), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT85), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n710), .A2(new_n711), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n730), .ZN(new_n732));
  NAND4_X1  g307(.A1(new_n710), .A2(new_n711), .A3(new_n727), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n729), .A2(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n697), .A2(G19), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n554), .B2(new_n697), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1341), .Z(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT29), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(G299), .A2(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n697), .A2(G20), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT23), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G1956), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  MUX2_X1   g326(.A(G104), .B(G116), .S(G2105), .Z(new_n752));
  AOI22_X1  g327(.A1(G128), .A2(new_n482), .B1(new_n752), .B2(G2104), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n471), .A2(G140), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT93), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT94), .B(G2067), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n615), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G4), .B2(G16), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT92), .B(G1348), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n759), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AND4_X1   g340(.A1(new_n738), .A2(new_n742), .A3(new_n748), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G34), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(new_n749), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT95), .Z(new_n769));
  INV_X1    g344(.A(G160), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(new_n749), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g348(.A1(G168), .A2(new_n697), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n697), .B2(G21), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT98), .B(G1966), .Z(new_n776));
  AOI21_X1  g351(.A(new_n773), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT27), .B(G1996), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT26), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G105), .B2(new_n472), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n471), .A2(G141), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n482), .A2(G129), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT96), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n785), .A2(G29), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G29), .B2(G32), .ZN(new_n787));
  OAI221_X1 g362(.A(new_n777), .B1(new_n775), .B2(new_n776), .C1(new_n778), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n749), .A2(G33), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n496), .A2(G127), .ZN(new_n790));
  NAND2_X1  g365(.A1(G115), .A2(G2104), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n481), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n472), .A2(G103), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT25), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n792), .B(new_n794), .C1(G139), .C2(new_n471), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n789), .B1(new_n795), .B2(new_n749), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G2072), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n771), .A2(new_n772), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n636), .A2(new_n749), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT31), .B(G11), .Z(new_n800));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n749), .B1(new_n801), .B2(G28), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n801), .B2(G28), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n788), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n697), .A2(G5), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G171), .B2(new_n697), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(G1961), .Z(new_n811));
  NOR2_X1   g386(.A1(G27), .A2(G29), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G164), .B2(G29), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT101), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT100), .B(G2078), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n787), .A2(new_n778), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT97), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n787), .A2(new_n819), .A3(new_n778), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n816), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n808), .A2(KEYINPUT102), .A3(new_n811), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n766), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n818), .A2(new_n820), .ZN(new_n824));
  INV_X1    g399(.A(new_n816), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n826), .A2(new_n788), .A3(new_n807), .ZN(new_n827));
  AOI21_X1  g402(.A(KEYINPUT102), .B1(new_n827), .B2(new_n811), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT103), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n808), .A2(new_n811), .A3(new_n821), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT103), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n832), .A2(new_n833), .A3(new_n822), .A4(new_n766), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n734), .A2(new_n735), .B1(new_n829), .B2(new_n834), .ZN(G311));
  NAND2_X1  g410(.A1(new_n734), .A2(new_n735), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n829), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(G150));
  XNOR2_X1  g413(.A(KEYINPUT105), .B(G860), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n532), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G651), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n525), .A2(G93), .B1(G55), .B2(new_n543), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n615), .A2(G559), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT104), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n843), .A2(new_n844), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n548), .A2(new_n850), .A3(new_n552), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n843), .B(new_n844), .C1(new_n550), .C2(new_n551), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n849), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(KEYINPUT106), .Z(new_n857));
  OAI21_X1  g432(.A(new_n839), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n846), .B1(new_n857), .B2(new_n858), .ZN(G145));
  INV_X1    g434(.A(KEYINPUT107), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n493), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n495), .A2(new_n498), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n491), .A2(new_n492), .A3(KEYINPUT107), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n756), .B(new_n864), .Z(new_n865));
  MUX2_X1   g440(.A(G106), .B(G118), .S(G2105), .Z(new_n866));
  AOI22_X1  g441(.A1(G130), .A2(new_n482), .B1(new_n866), .B2(G2104), .ZN(new_n867));
  INV_X1    g442(.A(G142), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n868), .B2(new_n624), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT108), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n721), .B(new_n628), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n865), .B(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n795), .A2(new_n784), .ZN(new_n874));
  INV_X1    g449(.A(new_n785), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n875), .B2(new_n795), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n873), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G162), .B(new_n770), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n636), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g458(.A1(new_n850), .A2(G868), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n619), .B(KEYINPUT109), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(new_n853), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n607), .A2(G299), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n607), .A2(G299), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OR2_X1    g469(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n889), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT42), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT42), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(G305), .B(G303), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n713), .A2(new_n704), .ZN(new_n904));
  NOR2_X1   g479(.A1(G290), .A2(G288), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n902), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n899), .A2(new_n910), .A3(new_n901), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n884), .B1(new_n912), .B2(G868), .ZN(G295));
  AOI21_X1  g488(.A(new_n884), .B1(new_n912), .B2(G868), .ZN(G331));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  NAND2_X1  g490(.A1(G171), .A2(G168), .ZN(new_n916));
  OAI21_X1  g491(.A(G286), .B1(new_n538), .B2(new_n541), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n853), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(new_n851), .A3(new_n852), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n893), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n896), .A3(new_n921), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n910), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n908), .A2(new_n923), .A3(new_n924), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n926), .A2(KEYINPUT43), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n892), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n887), .A2(KEYINPUT110), .A3(new_n891), .A4(new_n888), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n890), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n922), .A2(KEYINPUT111), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT111), .B1(new_n922), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n924), .B(KEYINPUT112), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n908), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n928), .A2(new_n927), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n915), .B(new_n929), .C1(new_n940), .C2(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n926), .A2(new_n942), .A3(new_n927), .A4(new_n928), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(KEYINPUT44), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT43), .B1(new_n938), .B2(new_n939), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT113), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n944), .B2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n941), .B1(new_n946), .B2(new_n947), .ZN(G397));
  INV_X1    g523(.A(G1384), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n864), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G40), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n474), .A2(new_n479), .A3(new_n951), .ZN(new_n952));
  XOR2_X1   g527(.A(KEYINPUT114), .B(KEYINPUT45), .Z(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G2067), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n756), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n784), .A2(G1996), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n957), .B(new_n958), .C1(G1996), .C2(new_n875), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n721), .B(new_n725), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(G290), .B(G1986), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n955), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n864), .A2(new_n965), .A3(new_n949), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n952), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT121), .B(G1961), .Z(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n864), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n953), .B1(G164), .B2(G1384), .ZN(new_n972));
  INV_X1    g547(.A(G2078), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n971), .A2(new_n972), .A3(new_n952), .A4(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT53), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n974), .A2(KEYINPUT122), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT122), .B1(new_n974), .B2(new_n975), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n975), .A2(new_n951), .A3(G2078), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n469), .B1(new_n496), .B2(G125), .ZN(new_n980));
  OAI211_X1 g555(.A(new_n473), .B(new_n979), .C1(new_n481), .C2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n950), .B2(new_n953), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n982), .A2(KEYINPUT123), .A3(new_n971), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT123), .B1(new_n982), .B2(new_n971), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(G171), .B1(new_n978), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n974), .A2(new_n975), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT122), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n974), .A2(KEYINPUT122), .A3(new_n975), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT69), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(new_n980), .B2(new_n481), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n994), .A2(G40), .A3(new_n473), .A4(new_n470), .ZN(new_n995));
  INV_X1    g570(.A(new_n953), .ZN(new_n996));
  AND2_X1   g571(.A1(new_n491), .A2(new_n492), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n862), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n995), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n950), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1001), .A3(new_n973), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n999), .A2(new_n1001), .A3(KEYINPUT120), .A4(new_n973), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n992), .A2(new_n1006), .A3(G301), .A4(new_n970), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n987), .A2(new_n1007), .A3(KEYINPUT54), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT124), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n987), .A2(new_n1007), .A3(KEYINPUT124), .A4(KEYINPUT54), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1996), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n971), .A2(new_n972), .A3(new_n952), .A4(new_n1013), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT58), .B(G1341), .Z(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n950), .B2(new_n995), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT119), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1017), .A2(new_n1018), .A3(new_n552), .A4(new_n548), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT59), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1017), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT119), .B1(new_n1021), .B2(new_n553), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(KEYINPUT119), .B(KEYINPUT59), .C1(new_n1021), .C2(new_n553), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT61), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n998), .A2(KEYINPUT116), .A3(new_n965), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT116), .B1(new_n998), .B2(new_n965), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n997), .A2(KEYINPUT107), .B1(new_n495), .B2(new_n498), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1384), .B1(new_n1030), .B2(new_n861), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n952), .B1(new_n1031), .B2(new_n965), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n747), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  XOR2_X1   g608(.A(KEYINPUT56), .B(G2072), .Z(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  AND4_X1   g610(.A1(new_n952), .A2(new_n971), .A3(new_n972), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n564), .A2(new_n568), .A3(new_n570), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1038), .B(new_n566), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n564), .A2(new_n568), .A3(KEYINPUT117), .A4(new_n570), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n1041));
  NAND3_X1  g616(.A1(G299), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1033), .A2(new_n1037), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1026), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n995), .B1(new_n950), .B2(KEYINPUT50), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1036), .B1(new_n1048), .B2(new_n747), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1026), .B1(new_n1049), .B2(new_n1043), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n1039), .A2(new_n1042), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1028), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n998), .A2(KEYINPUT116), .A3(new_n965), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1956), .B1(new_n1056), .B2(new_n1047), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1052), .A2(new_n1053), .B1(new_n1057), .B2(new_n1036), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n762), .ZN(new_n1060));
  INV_X1    g635(.A(new_n998), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n995), .B1(new_n1061), .B2(KEYINPUT50), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1062), .B2(new_n966), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n950), .A2(new_n995), .A3(G2067), .ZN(new_n1064));
  NOR4_X1   g639(.A1(new_n1063), .A2(KEYINPUT60), .A3(new_n607), .A4(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n615), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n968), .A2(new_n762), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1064), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n607), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1070), .B2(KEYINPUT60), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1025), .A2(new_n1046), .A3(new_n1059), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1049), .A2(new_n1043), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1066), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1075), .A2(new_n1058), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1005), .ZN(new_n1078));
  OAI21_X1  g653(.A(G171), .B1(new_n1078), .B2(new_n978), .ZN(new_n1079));
  INV_X1    g654(.A(new_n985), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(new_n983), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n992), .A2(new_n1081), .A3(G301), .A4(new_n970), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT54), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n862), .A2(new_n997), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n949), .A3(new_n996), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n952), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT45), .B1(new_n864), .B2(new_n949), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n776), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n966), .A2(new_n967), .A3(new_n952), .A4(new_n772), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(G168), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT51), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  OAI211_X1 g669(.A(G8), .B(new_n1090), .C1(new_n1093), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1976), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(G288), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G8), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1031), .B2(new_n952), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n574), .B(G1976), .C1(new_n575), .C2(new_n515), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1101), .ZN(new_n1103));
  OAI21_X1  g678(.A(G8), .B1(new_n950), .B2(new_n995), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT52), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND2_X1   g680(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n514), .B2(new_n519), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT55), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1107), .B(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n995), .B1(new_n1061), .B2(new_n953), .ZN(new_n1110));
  AOI21_X1  g685(.A(G1971), .B1(new_n1110), .B2(new_n971), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n968), .A2(G2090), .ZN(new_n1112));
  OAI211_X1 g687(.A(G8), .B(new_n1109), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n577), .B(new_n578), .C1(new_n584), .C2(KEYINPUT78), .ZN(new_n1115));
  NOR3_X1   g690(.A1(new_n1115), .A2(G1981), .A3(new_n588), .ZN(new_n1116));
  OAI21_X1  g691(.A(G1981), .B1(new_n579), .B2(new_n584), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1114), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(KEYINPUT49), .B(new_n1117), .C1(G305), .C2(G1981), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1100), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1106), .A2(new_n1113), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1048), .A2(G2090), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1123), .B2(new_n1111), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1109), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1096), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1083), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1012), .A2(new_n1077), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n704), .A2(new_n1097), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1116), .B1(new_n1121), .B2(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1100), .B(KEYINPUT115), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1106), .A2(new_n1121), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n1133), .A2(new_n1134), .B1(new_n1135), .B2(new_n1113), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1139), .A2(G8), .A3(G168), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1137), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(G8), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1137), .B(new_n1140), .C1(new_n1125), .C2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1122), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1136), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1129), .A2(new_n1130), .A3(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1138), .A2(new_n1079), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT62), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1092), .A2(new_n1095), .A3(KEYINPUT62), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1146), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1130), .B1(new_n1129), .B2(new_n1145), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n964), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n784), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n954), .B1(new_n957), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT126), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n955), .A2(new_n1013), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT46), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT47), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n721), .A2(new_n725), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n959), .A2(new_n1161), .B1(G2067), .B2(new_n756), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(new_n955), .ZN(new_n1163));
  NOR2_X1   g738(.A1(G290), .A2(G1986), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1164), .A2(KEYINPUT48), .A3(new_n955), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT48), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1164), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1166), .B1(new_n1167), .B2(new_n954), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(new_n1168), .C1(new_n961), .C2(new_n954), .ZN(new_n1169));
  AND3_X1   g744(.A1(new_n1160), .A2(new_n1163), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1153), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g746(.A1(G319), .A2(new_n655), .ZN(new_n1173));
  AND3_X1   g747(.A1(new_n1173), .A2(KEYINPUT127), .A3(new_n671), .ZN(new_n1174));
  AOI21_X1  g748(.A(KEYINPUT127), .B1(new_n1173), .B2(new_n671), .ZN(new_n1175));
  OAI21_X1  g749(.A(new_n692), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g750(.A(new_n1176), .B1(new_n880), .B2(new_n881), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n1177), .B(new_n929), .C1(KEYINPUT43), .C2(new_n940), .ZN(G225));
  INV_X1    g752(.A(G225), .ZN(G308));
endmodule


