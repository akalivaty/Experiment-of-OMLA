//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:49 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325;
  XOR2_X1   g0000(.A(KEYINPUT65), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(KEYINPUT64), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND3_X1  g0004(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G77), .ZN(new_n208));
  AND3_X1   g0008(.A1(new_n201), .A2(new_n207), .A3(new_n208), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n212), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G107), .ZN(new_n226));
  INV_X1    g0026(.A(G264), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n208), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n214), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n217), .B1(new_n220), .B2(new_n223), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT2), .B(G226), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G264), .B(G270), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT67), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NAND2_X1  g0051(.A1(new_n236), .A2(G1698), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n252), .B1(G226), .B2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G97), .ZN(new_n259));
  OAI22_X1  g0059(.A1(new_n253), .A2(new_n258), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n260), .A2(new_n263), .B1(G238), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(G274), .B1(new_n269), .B2(new_n218), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n270), .B2(new_n264), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  AND2_X1   g0072(.A1(G1), .A2(G13), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n272), .B1(new_n273), .B2(new_n261), .ZN(new_n274));
  INV_X1    g0074(.A(new_n264), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(KEYINPUT68), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT13), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n267), .A2(new_n280), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(G169), .ZN(new_n284));
  INV_X1    g0084(.A(G179), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(new_n282), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n283), .B1(new_n282), .B2(G169), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G20), .A2(G33), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n288), .A2(G50), .B1(G20), .B2(new_n204), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n212), .A2(G33), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n289), .B1(new_n208), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n218), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT11), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G13), .ZN(new_n295));
  NOR3_X1   g0095(.A1(new_n295), .A2(new_n212), .A3(G1), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n204), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT12), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n291), .A2(KEYINPUT11), .A3(new_n293), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n296), .A2(new_n293), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n211), .A2(G20), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n300), .A2(G68), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n298), .A2(new_n299), .A3(new_n302), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n286), .A2(new_n287), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n221), .B1(new_n211), .B2(G20), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n300), .A2(new_n305), .B1(new_n221), .B2(new_n296), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT71), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n306), .B(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n212), .B1(new_n201), .B2(new_n207), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n288), .A2(G150), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT8), .B(G58), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n311), .B2(new_n290), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n293), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n308), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT3), .B(G33), .ZN(new_n317));
  INV_X1    g0117(.A(G1698), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n317), .A2(G222), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT69), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n319), .B(new_n320), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n258), .A2(new_n318), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G223), .B1(G77), .B2(new_n258), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n262), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G226), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n277), .B1(new_n325), .B2(new_n265), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n328), .A2(KEYINPUT72), .A3(G179), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT72), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n327), .B2(new_n285), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n316), .B(new_n330), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n282), .A2(G200), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n303), .A2(new_n294), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n282), .ZN(new_n338));
  INV_X1    g0138(.A(new_n293), .ZN(new_n339));
  INV_X1    g0139(.A(new_n311), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n340), .A2(new_n288), .B1(G20), .B2(G77), .ZN(new_n341));
  XOR2_X1   g0141(.A(KEYINPUT15), .B(G87), .Z(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n212), .A3(G33), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n339), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n300), .A2(G77), .A3(new_n301), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n295), .A2(G1), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G20), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n345), .B1(G77), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n266), .A2(G244), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n317), .A2(G232), .A3(new_n318), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n226), .B2(new_n317), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G238), .B2(new_n322), .ZN(new_n353));
  OAI211_X1 g0153(.A(new_n277), .B(new_n350), .C1(new_n353), .C2(new_n262), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n354), .B2(new_n329), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(G179), .B2(new_n354), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n354), .A2(G200), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n349), .C1(new_n337), .C2(new_n354), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n304), .A2(new_n334), .A3(new_n338), .A4(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n316), .B(KEYINPUT9), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT10), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n327), .A2(G190), .ZN(new_n363));
  OAI21_X1  g0163(.A(G200), .B1(new_n324), .B2(new_n326), .ZN(new_n364));
  AND2_X1   g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n361), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT16), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT7), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n317), .B2(G20), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n258), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n204), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G58), .A2(G68), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n205), .A2(new_n206), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n288), .A2(G159), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n370), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT74), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n376), .A2(G20), .B1(G159), .B2(new_n288), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT73), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n256), .B2(KEYINPUT3), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n254), .A2(KEYINPUT73), .A3(G33), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(new_n257), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(new_n371), .A3(new_n212), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G68), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n371), .B1(new_n387), .B2(new_n212), .ZN(new_n390));
  OAI211_X1 g0190(.A(KEYINPUT16), .B(new_n383), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  OAI211_X1 g0191(.A(KEYINPUT74), .B(new_n370), .C1(new_n374), .C2(new_n379), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n382), .A2(new_n293), .A3(new_n391), .A4(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n300), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n340), .A2(new_n301), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n394), .A2(new_n395), .B1(new_n347), .B2(new_n340), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT75), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n270), .A2(new_n268), .A3(new_n264), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT68), .B1(new_n274), .B2(new_n275), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n401), .A2(new_n402), .B1(new_n236), .B2(new_n265), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G223), .A2(G1698), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n325), .B2(G1698), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(new_n385), .A3(new_n386), .A4(new_n257), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n262), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n400), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n262), .A2(G232), .A3(new_n264), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n271), .B2(new_n276), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n325), .A2(G1698), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(G223), .B2(G1698), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n407), .B1(new_n387), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n263), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT75), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n403), .A2(new_n408), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n417), .A2(new_n329), .B1(new_n285), .B2(new_n418), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n398), .A2(new_n399), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n399), .B1(new_n398), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT77), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT7), .B1(new_n258), .B2(new_n212), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n371), .B(G20), .C1(new_n255), .C2(new_n257), .ZN(new_n425));
  OAI21_X1  g0225(.A(G68), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n383), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT74), .B1(new_n427), .B2(new_n370), .ZN(new_n428));
  INV_X1    g0228(.A(new_n392), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n391), .A2(new_n293), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n396), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(G200), .B1(new_n409), .B2(new_n416), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT76), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n403), .A2(new_n408), .A3(G190), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G200), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n411), .A2(new_n415), .A3(KEYINPUT75), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT75), .B1(new_n411), .B2(new_n415), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n435), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT76), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n432), .B(KEYINPUT17), .C1(new_n436), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n434), .B1(new_n433), .B2(new_n435), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n440), .A2(KEYINPUT76), .A3(new_n441), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(KEYINPUT17), .B1(new_n447), .B2(new_n432), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n423), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n432), .B1(new_n436), .B2(new_n442), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT17), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(KEYINPUT77), .A3(new_n443), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n369), .A2(new_n422), .A3(new_n449), .A4(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n385), .A2(new_n386), .A3(new_n257), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT89), .A3(G250), .A4(new_n318), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT89), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n385), .A2(new_n386), .A3(new_n318), .A4(new_n257), .ZN(new_n458));
  INV_X1    g0258(.A(G250), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g0260(.A1(G257), .A2(G1698), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n385), .A2(new_n386), .A3(new_n257), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G294), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n456), .A2(new_n460), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT90), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n262), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n456), .A2(new_n464), .A3(new_n460), .A4(KEYINPUT90), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n211), .A2(G45), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT5), .B(G41), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n274), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n471), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G264), .A3(new_n262), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n469), .A2(G190), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n211), .A2(G33), .ZN(new_n477));
  AND3_X1   g0277(.A1(new_n339), .A2(new_n347), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(KEYINPUT25), .B1(new_n296), .B2(new_n226), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n226), .ZN(new_n481));
  AOI22_X1  g0281(.A1(G107), .A2(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT80), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT80), .A2(G116), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n212), .A3(G33), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT88), .A2(KEYINPUT23), .ZN(new_n491));
  OAI211_X1 g0291(.A(G20), .B(new_n226), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  OAI22_X1  g0292(.A1(new_n212), .A2(G107), .B1(KEYINPUT88), .B2(KEYINPUT23), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(G87), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G20), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT22), .B1(new_n317), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT24), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n385), .A2(new_n386), .A3(new_n212), .A4(new_n257), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  NOR3_X1   g0301(.A1(new_n500), .A2(new_n501), .A3(new_n495), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n317), .A2(new_n496), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n501), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n506), .A2(new_n489), .A3(new_n493), .A4(new_n492), .ZN(new_n507));
  OAI21_X1  g0307(.A(KEYINPUT24), .B1(new_n507), .B2(new_n502), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n483), .B1(new_n509), .B2(new_n293), .ZN(new_n510));
  INV_X1    g0310(.A(new_n473), .ZN(new_n511));
  INV_X1    g0311(.A(new_n475), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n467), .C2(new_n468), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n476), .B(new_n510), .C1(new_n513), .C2(new_n437), .ZN(new_n514));
  OR2_X1    g0314(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g0315(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n259), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(KEYINPUT79), .A3(new_n516), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g0320(.A(G97), .B(G107), .Z(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n519), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n522), .A2(G20), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n372), .A2(new_n373), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(G107), .B1(G77), .B2(new_n288), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n293), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n317), .A2(G250), .A3(G1698), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n225), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n532), .A2(new_n318), .A3(new_n255), .A4(new_n257), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n531), .B1(new_n458), .B2(new_n225), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n262), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n474), .A2(G257), .A3(new_n262), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n473), .ZN(new_n539));
  OAI21_X1  g0339(.A(G200), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n539), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n455), .A2(G244), .A3(new_n318), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(new_n531), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G190), .B(new_n541), .C1(new_n544), .C2(new_n262), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n347), .A2(G97), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n546), .B1(new_n478), .B2(G97), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n529), .A2(new_n540), .A3(new_n545), .A4(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n329), .B1(new_n537), .B2(new_n539), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n285), .B(new_n541), .C1(new_n544), .C2(new_n262), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n339), .B1(new_n525), .B2(new_n527), .ZN(new_n551));
  INV_X1    g0351(.A(new_n547), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  AND2_X1   g0353(.A1(new_n548), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n486), .A2(new_n487), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n478), .A2(G116), .B1(new_n296), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n486), .A2(G20), .A3(new_n487), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n534), .B(new_n212), .C1(G33), .C2(new_n259), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n293), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT20), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n558), .A4(new_n293), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n474), .A2(G270), .A3(new_n262), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n565), .A2(new_n473), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n254), .A2(G33), .ZN(new_n568));
  OAI21_X1  g0368(.A(G303), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n227), .A2(G1698), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(G257), .B2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n569), .B1(new_n387), .B2(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n572), .A2(KEYINPUT86), .A3(new_n263), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT86), .B1(new_n572), .B2(new_n263), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n566), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n564), .B1(new_n575), .B2(G200), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n337), .B2(new_n575), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n514), .A2(new_n554), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n329), .B1(new_n556), .B2(new_n563), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n575), .A2(new_n579), .A3(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n572), .A2(new_n263), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT86), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n572), .A2(KEYINPUT86), .A3(new_n263), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n565), .A2(G179), .A3(new_n473), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n564), .A3(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n580), .A2(KEYINPUT87), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT87), .B1(new_n580), .B2(new_n587), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT21), .B1(new_n575), .B2(new_n579), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n469), .A2(new_n285), .A3(new_n473), .A4(new_n475), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n499), .B1(new_n498), .B2(new_n503), .ZN(new_n593));
  NOR3_X1   g0393(.A1(new_n507), .A2(KEYINPUT24), .A3(new_n502), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n293), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n482), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n592), .B(new_n596), .C1(new_n513), .C2(G169), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n274), .A2(new_n471), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n262), .A2(G250), .A3(new_n470), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n225), .A2(G1698), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(G238), .B2(G1698), .ZN(new_n602));
  OAI22_X1  g0402(.A1(new_n387), .A2(new_n602), .B1(new_n555), .B2(new_n256), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n603), .B2(new_n263), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n285), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n605), .B(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n478), .A2(new_n342), .ZN(new_n607));
  INV_X1    g0407(.A(new_n342), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n296), .ZN(new_n609));
  NAND3_X1  g0409(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n610), .A2(KEYINPUT82), .A3(new_n212), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n495), .A2(new_n259), .A3(new_n226), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT82), .B1(new_n610), .B2(new_n212), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n290), .A2(new_n259), .ZN(new_n615));
  OAI22_X1  g0415(.A1(new_n613), .A2(new_n614), .B1(KEYINPUT19), .B2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n455), .A2(KEYINPUT83), .A3(new_n212), .A4(G68), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT83), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n500), .B2(new_n204), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n293), .B1(new_n620), .B2(KEYINPUT84), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT84), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n622), .B(new_n616), .C1(new_n619), .C2(new_n617), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n607), .B(new_n609), .C1(new_n621), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n603), .A2(new_n263), .ZN(new_n625));
  INV_X1    g0425(.A(new_n600), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n329), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n606), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n478), .A2(G87), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n627), .B2(G200), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n631), .B(new_n609), .C1(new_n621), .C2(new_n623), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT85), .ZN(new_n633));
  AND2_X1   g0433(.A1(new_n617), .A2(new_n619), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n622), .B1(new_n634), .B2(new_n616), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n620), .A2(KEYINPUT84), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n293), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT85), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n637), .A2(new_n638), .A3(new_n609), .A4(new_n631), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n604), .A2(G190), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n591), .A2(new_n597), .A3(new_n629), .A4(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n454), .A2(new_n578), .A3(new_n642), .ZN(G372));
  INV_X1    g0443(.A(KEYINPUT92), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n368), .B(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n356), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n338), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n304), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n449), .A2(new_n648), .A3(new_n453), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n422), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n651), .A2(new_n334), .ZN(new_n652));
  INV_X1    g0452(.A(new_n454), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n632), .A2(KEYINPUT85), .B1(G190), .B2(new_n604), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n624), .A2(new_n628), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n639), .A2(new_n654), .B1(new_n655), .B2(new_n606), .ZN(new_n656));
  INV_X1    g0456(.A(new_n553), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(KEYINPUT91), .A3(KEYINPUT26), .A4(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n624), .A2(new_n605), .A3(new_n628), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n637), .A2(new_n609), .A3(new_n631), .A4(new_n640), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n657), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT91), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n641), .A2(new_n629), .A3(KEYINPUT26), .A4(new_n657), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n580), .A2(new_n587), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n590), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n597), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n659), .A2(new_n660), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n554), .A4(new_n514), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n658), .A2(new_n665), .A3(new_n659), .A4(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n653), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n652), .A2(new_n672), .ZN(G369));
  NAND2_X1  g0473(.A1(new_n346), .A2(new_n212), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  XOR2_X1   g0475(.A(new_n675), .B(KEYINPUT93), .Z(new_n676));
  INV_X1    g0476(.A(G213), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G343), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n514), .B1(new_n510), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n597), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n680), .A2(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n597), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n577), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n564), .ZN(new_n689));
  NOR3_X1   g0489(.A1(new_n689), .A2(new_n666), .A3(new_n590), .ZN(new_n690));
  INV_X1    g0490(.A(new_n591), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n688), .B(new_n690), .C1(new_n691), .C2(new_n689), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G330), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n682), .A2(new_n597), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n591), .A2(new_n684), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n685), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n215), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n612), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n223), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n671), .A2(new_n707), .A3(new_n681), .ZN(new_n708));
  INV_X1    g0508(.A(new_n659), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n709), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n641), .A2(new_n629), .A3(new_n662), .A4(new_n657), .ZN(new_n711));
  INV_X1    g0511(.A(new_n588), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT87), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n590), .B1(new_n666), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n597), .A2(new_n712), .A3(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n514), .A2(new_n554), .A3(new_n659), .A4(new_n660), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n710), .B(new_n711), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT29), .B1(new_n718), .B2(new_n684), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n708), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n469), .A2(new_n475), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n537), .A2(new_n539), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n585), .A3(new_n586), .A4(new_n604), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n604), .B(new_n586), .C1(new_n573), .C2(new_n574), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n541), .B1(new_n544), .B2(new_n262), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT30), .A3(new_n475), .A4(new_n469), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n469), .A2(new_n473), .A3(new_n475), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n604), .A2(G179), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n728), .A2(new_n575), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n726), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT31), .B1(new_n735), .B2(new_n684), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n578), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(new_n715), .A3(new_n656), .A4(new_n681), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n721), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n720), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n706), .B1(new_n742), .B2(G1), .ZN(G364));
  XOR2_X1   g0543(.A(new_n693), .B(KEYINPUT94), .Z(new_n744));
  NOR2_X1   g0544(.A1(new_n295), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n211), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR3_X1    g0547(.A1(new_n701), .A2(KEYINPUT95), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT95), .B1(new_n701), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n744), .B(new_n750), .C1(G330), .C2(new_n692), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n215), .A2(G355), .A3(new_n317), .ZN(new_n752));
  INV_X1    g0552(.A(G45), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n247), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n700), .A2(new_n455), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n223), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n752), .B1(G116), .B2(new_n215), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n218), .B1(G20), .B2(new_n329), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n750), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n761), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT97), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(G190), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT98), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(KEYINPUT98), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G159), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT32), .Z(new_n774));
  AND2_X1   g0574(.A1(new_n766), .A2(G190), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n212), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n259), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n285), .A2(G200), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n778), .A2(G20), .A3(G190), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n767), .A2(new_n778), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n203), .B1(new_n780), .B2(new_n208), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT96), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n212), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n337), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n258), .B1(new_n787), .B2(G107), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n783), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n495), .ZN(new_n791));
  NAND3_X1  g0591(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n792), .A2(new_n337), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n794), .A2(new_n204), .B1(new_n796), .B2(new_n221), .ZN(new_n797));
  NOR4_X1   g0597(.A1(new_n777), .A2(new_n789), .A3(new_n791), .A4(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n779), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT33), .B(G317), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n799), .A2(G322), .B1(new_n793), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(KEYINPUT100), .ZN(new_n802));
  INV_X1    g0602(.A(G294), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  INV_X1    g0604(.A(new_n790), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n317), .B1(new_n805), .B2(G303), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n776), .A2(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n802), .B(new_n807), .C1(new_n804), .C2(new_n806), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n801), .A2(KEYINPUT100), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n795), .A2(G326), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n780), .B2(new_n811), .C1(new_n812), .C2(new_n786), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n809), .B(new_n813), .C1(new_n772), .C2(G329), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n774), .A2(new_n798), .B1(new_n808), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n760), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n763), .B1(new_n764), .B2(new_n815), .C1(new_n692), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n751), .A2(new_n817), .ZN(G396));
  INV_X1    g0618(.A(new_n750), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n359), .A2(new_n681), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n671), .A2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n671), .A2(new_n681), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n356), .A2(new_n684), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n358), .B1(new_n349), .B2(new_n681), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n356), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n821), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n741), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n819), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n761), .A2(new_n758), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n819), .B1(G77), .B2(new_n831), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n258), .B1(new_n779), .B2(new_n803), .C1(new_n555), .C2(new_n780), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n787), .A2(G87), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(new_n794), .B2(new_n812), .ZN(new_n835));
  INV_X1    g0635(.A(G303), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n796), .A2(new_n836), .B1(new_n790), .B2(new_n226), .ZN(new_n837));
  NOR4_X1   g0637(.A1(new_n777), .A2(new_n833), .A3(new_n835), .A4(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n772), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n838), .B1(new_n811), .B2(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n793), .A2(G150), .B1(new_n795), .B2(G137), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT101), .Z(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  INV_X1    g0643(.A(G159), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n779), .C1(new_n844), .C2(new_n780), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT34), .Z(new_n846));
  NOR2_X1   g0646(.A1(new_n786), .A2(new_n204), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n387), .B(new_n847), .C1(G50), .C2(new_n805), .ZN(new_n848));
  INV_X1    g0648(.A(G132), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n203), .B2(new_n776), .C1(new_n839), .C2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n840), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n832), .B1(new_n851), .B2(new_n761), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n759), .B2(new_n825), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n829), .A2(new_n853), .ZN(G384));
  NOR2_X1   g0654(.A1(new_n745), .A2(new_n211), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n304), .A2(new_n338), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n681), .A2(new_n336), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n738), .A2(new_n740), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n858), .A2(new_n859), .A3(new_n825), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n398), .A2(new_n680), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT103), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n398), .A2(new_n419), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n864), .A2(new_n865), .A3(new_n450), .A4(new_n862), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n679), .B1(new_n393), .B2(new_n397), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n867), .B2(KEYINPUT103), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n865), .A2(new_n862), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n398), .B1(new_n445), .B2(new_n446), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n422), .A2(new_n452), .A3(new_n443), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n867), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n872), .B1(new_n874), .B2(KEYINPUT104), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT104), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n873), .A2(new_n876), .A3(new_n867), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n417), .A2(new_n329), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n418), .A2(new_n285), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n383), .B1(new_n389), .B2(new_n390), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n370), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n431), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n882), .A2(new_n679), .B1(new_n397), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(KEYINPUT37), .B1(new_n886), .B2(new_n870), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n450), .A2(new_n861), .A3(new_n865), .A4(new_n862), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n449), .A2(new_n422), .A3(new_n453), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n679), .B1(new_n885), .B2(new_n397), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n879), .B(new_n889), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n860), .B1(new_n878), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n890), .A2(new_n891), .ZN(new_n894));
  INV_X1    g0694(.A(new_n889), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n879), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n858), .A2(new_n859), .A3(new_n825), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n900), .A2(KEYINPUT40), .ZN(new_n901));
  AOI22_X1  g0701(.A1(KEYINPUT40), .A2(new_n893), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n454), .B1(new_n740), .B2(new_n738), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n721), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n903), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT39), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n878), .B2(new_n892), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n304), .A2(new_n684), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n908), .B(new_n910), .C1(new_n899), .C2(new_n907), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n422), .A2(new_n680), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n823), .B1(new_n671), .B2(new_n820), .ZN(new_n913));
  INV_X1    g0713(.A(new_n858), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n899), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n720), .A2(new_n653), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n652), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n917), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n855), .B1(new_n906), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n920), .B2(new_n906), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n522), .A2(new_n524), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n485), .B(new_n220), .C1(new_n923), .C2(KEYINPUT35), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(KEYINPUT35), .B2(new_n923), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT36), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n222), .A2(G77), .A3(new_n375), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(KEYINPUT102), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n201), .A2(G68), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n927), .B2(KEYINPUT102), .ZN(new_n930));
  OAI211_X1 g0730(.A(G1), .B(new_n295), .C1(new_n928), .C2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n926), .A3(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n637), .A2(new_n609), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n684), .B1(new_n933), .B2(new_n630), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n669), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n659), .B2(new_n934), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT107), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n553), .A2(new_n681), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT105), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n684), .B1(new_n551), .B2(new_n552), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n554), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n686), .A2(new_n697), .A3(new_n944), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n945), .A2(KEYINPUT42), .B1(new_n657), .B2(new_n681), .ZN(new_n946));
  INV_X1    g0746(.A(new_n685), .ZN(new_n947));
  INV_X1    g0747(.A(new_n697), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n947), .B1(new_n683), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(KEYINPUT42), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n944), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n946), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n937), .A2(new_n938), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n939), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n938), .B(new_n937), .C1(new_n952), .C2(new_n954), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n944), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n695), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n959), .B(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n701), .B(KEYINPUT41), .Z(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT109), .B1(new_n686), .B2(new_n697), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n686), .A2(new_n697), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n964), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n744), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n693), .B2(new_n966), .ZN(new_n968));
  INV_X1    g0768(.A(new_n742), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n698), .A2(new_n944), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT44), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n698), .B2(new_n944), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n949), .A2(KEYINPUT44), .A3(new_n960), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(KEYINPUT108), .A3(new_n974), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n979), .A2(new_n694), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n694), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n970), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n963), .B1(new_n983), .B2(new_n742), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n962), .B1(new_n984), .B2(new_n747), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n936), .A2(new_n816), .ZN(new_n986));
  INV_X1    g0786(.A(new_n755), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n762), .B1(new_n215), .B2(new_n608), .C1(new_n987), .C2(new_n242), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n819), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n772), .A2(G137), .ZN(new_n990));
  INV_X1    g0790(.A(G150), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n317), .B1(new_n779), .B2(new_n991), .C1(new_n201), .C2(new_n780), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n796), .A2(new_n843), .B1(new_n786), .B2(new_n208), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n794), .A2(new_n844), .B1(new_n790), .B2(new_n203), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n990), .B(new_n995), .C1(new_n204), .C2(new_n776), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n776), .A2(new_n226), .B1(new_n812), .B2(new_n780), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT110), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n772), .A2(G317), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n259), .B2(new_n786), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT46), .B1(new_n805), .B2(new_n488), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n387), .B1(new_n794), .B2(new_n803), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n799), .A2(G303), .B1(G311), .B2(new_n795), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT111), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n999), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n996), .B1(new_n998), .B2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n989), .B1(new_n1010), .B2(new_n761), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n986), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n985), .A2(new_n1012), .ZN(G387));
  AND2_X1   g0813(.A1(new_n968), .A2(new_n969), .ZN(new_n1014));
  OR3_X1    g0814(.A1(new_n1014), .A2(new_n970), .A3(new_n702), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n762), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n703), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(new_n215), .A3(new_n317), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(G107), .B2(new_n215), .ZN(new_n1019));
  OR2_X1    g0819(.A1(new_n239), .A2(new_n753), .ZN(new_n1020));
  AOI211_X1 g0820(.A(G45), .B(new_n1017), .C1(G68), .C2(G77), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n311), .A2(G50), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT50), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n987), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1019), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n776), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n342), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n780), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n799), .A2(G50), .B1(new_n1028), .B2(G68), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n805), .A2(G77), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n794), .B2(new_n311), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n796), .A2(new_n844), .B1(new_n786), .B2(new_n259), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1027), .A2(new_n455), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G150), .B2(new_n772), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n799), .A2(G317), .B1(new_n1028), .B2(G303), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(KEYINPUT114), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n793), .A2(G311), .B1(new_n795), .B2(G322), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT48), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1026), .A2(G283), .B1(G294), .B2(new_n805), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT49), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n387), .B1(new_n555), .B2(new_n786), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n772), .B2(G326), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1035), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n819), .B1(new_n1016), .B2(new_n1025), .C1(new_n1049), .C2(new_n764), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n687), .B2(new_n760), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT113), .ZN(new_n1052));
  OR3_X1    g0852(.A1(new_n968), .A2(new_n1052), .A3(new_n746), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n968), .B2(new_n746), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1015), .A2(new_n1055), .ZN(G393));
  INV_X1    g0856(.A(new_n982), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1057), .A2(new_n746), .A3(new_n980), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n960), .A2(new_n760), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n834), .B1(new_n204), .B2(new_n790), .C1(new_n794), .C2(new_n201), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n387), .B(new_n1060), .C1(new_n340), .C2(new_n1028), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n796), .A2(new_n991), .B1(new_n779), .B2(new_n844), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT51), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1026), .A2(G77), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n772), .A2(G143), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n772), .A2(G322), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n799), .A2(G311), .B1(G317), .B2(new_n795), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n1026), .A2(new_n488), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n258), .B1(new_n780), .B2(new_n803), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n794), .A2(new_n836), .B1(new_n790), .B2(new_n812), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G107), .C2(new_n787), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n764), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n987), .A2(new_n250), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1016), .B(new_n1077), .C1(G97), .C2(new_n700), .ZN(new_n1078));
  NOR3_X1   g0878(.A1(new_n1076), .A2(new_n750), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1058), .B1(new_n1059), .B2(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n980), .A2(new_n1057), .B1(new_n969), .B2(new_n968), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n983), .A3(new_n701), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(G390));
  INV_X1    g0883(.A(KEYINPUT115), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1084), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n909), .B1(new_n913), .B2(new_n914), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(KEYINPUT115), .ZN(new_n1087));
  AOI21_X1  g0887(.A(KEYINPUT38), .B1(new_n894), .B2(new_n895), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1088), .A2(new_n892), .A3(new_n907), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n874), .A2(KEYINPUT104), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n872), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1090), .A2(new_n877), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n879), .ZN(new_n1093));
  AOI21_X1  g0893(.A(KEYINPUT39), .B1(new_n1093), .B2(new_n898), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1085), .B(new_n1087), .C1(new_n1089), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n824), .A2(new_n356), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n717), .A2(new_n681), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n823), .ZN(new_n1098));
  AND2_X1   g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n909), .B1(new_n1099), .B2(new_n914), .C1(new_n892), .C2(new_n878), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1095), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n741), .A2(new_n825), .A3(new_n858), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1095), .A2(new_n1102), .A3(new_n1100), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(new_n746), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1108), .A2(new_n759), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n258), .B1(new_n780), .B2(new_n259), .C1(new_n485), .C2(new_n779), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n791), .A2(new_n847), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n794), .B2(new_n226), .C1(new_n812), .C2(new_n796), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1110), .B(new_n1112), .C1(G77), .C2(new_n1026), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n772), .A2(G294), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n790), .A2(new_n991), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n776), .B2(new_n844), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(KEYINPUT54), .B(G143), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n317), .B1(new_n780), .B2(new_n1118), .C1(new_n849), .C2(new_n779), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n793), .A2(G137), .B1(new_n795), .B2(G128), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1120), .B1(new_n201), .B2(new_n786), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n772), .A2(G125), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1113), .A2(new_n1114), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n819), .B1(new_n340), .B2(new_n831), .C1(new_n1124), .C2(new_n764), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1109), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1107), .A2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n642), .A2(new_n578), .A3(new_n684), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n735), .A2(new_n684), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT31), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n684), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g0933(.A(G330), .B(new_n825), .C1(new_n1128), .C2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n914), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1135), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n913), .B1(new_n1135), .B2(new_n1102), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n827), .A2(new_n454), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n918), .A2(new_n1140), .A3(new_n652), .ZN(new_n1141));
  OAI21_X1  g0941(.A(KEYINPUT116), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1135), .A2(new_n1102), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n913), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1135), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n454), .B1(new_n708), .B2(new_n719), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n651), .A2(new_n334), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1139), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT116), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1142), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1104), .A2(new_n1105), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n701), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT117), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1105), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1102), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1158));
  OAI21_X1  g0958(.A(KEYINPUT118), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT118), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1104), .A2(new_n1160), .A3(new_n1105), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1153), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1161), .A3(KEYINPUT119), .A4(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT117), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1154), .A2(new_n1164), .A3(new_n701), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1156), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1153), .B1(new_n1106), .B2(KEYINPUT118), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT119), .B1(new_n1167), .B2(new_n1161), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1127), .B1(new_n1166), .B2(new_n1168), .ZN(G378));
  OAI221_X1 g0969(.A(new_n1030), .B1(new_n226), .B2(new_n779), .C1(new_n608), .C2(new_n780), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n794), .A2(new_n259), .B1(new_n796), .B2(new_n485), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n786), .A2(new_n203), .ZN(new_n1172));
  INV_X1    g0972(.A(G41), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n387), .A2(new_n1173), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1174), .ZN(new_n1175));
  OAI221_X1 g0975(.A(new_n1175), .B1(new_n204), .B2(new_n776), .C1(new_n812), .C2(new_n839), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT58), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G50), .B1(new_n256), .B2(new_n1173), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1176), .A2(new_n1177), .B1(new_n1174), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1118), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n805), .A2(new_n1180), .B1(G125), .B2(new_n795), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n799), .A2(G128), .B1(new_n1028), .B2(G137), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n849), .C2(new_n794), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n1026), .B2(G150), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n256), .B(new_n1173), .C1(new_n786), .C2(new_n844), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n772), .B2(G124), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT59), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1188), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n1179), .B1(new_n1177), .B2(new_n1176), .C1(new_n1186), .C2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n761), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n750), .B1(new_n201), .B2(new_n830), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n645), .A2(new_n334), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n316), .A2(new_n680), .ZN(new_n1196));
  XOR2_X1   g0996(.A(new_n1196), .B(KEYINPUT55), .Z(new_n1197));
  XNOR2_X1  g0997(.A(new_n1195), .B(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n1199));
  XNOR2_X1  g0999(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1194), .B1(new_n1201), .B2(new_n758), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n911), .B(new_n916), .C1(new_n902), .C2(new_n721), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n893), .A2(KEYINPUT40), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n899), .A2(new_n901), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n721), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n917), .A2(new_n1207), .ZN(new_n1208));
  AND3_X1   g1008(.A1(new_n1204), .A2(new_n1208), .A3(new_n1200), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1200), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1203), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1204), .A2(new_n1208), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1201), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1204), .A2(new_n1208), .A3(new_n1200), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(KEYINPUT121), .A3(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1202), .B1(new_n1216), .B2(new_n747), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1154), .A2(new_n1150), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT122), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1154), .A2(KEYINPUT122), .A3(new_n1150), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1213), .A2(KEYINPUT57), .A3(new_n1214), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1154), .A2(KEYINPUT122), .A3(new_n1150), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT122), .B1(new_n1154), .B2(new_n1150), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n701), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1217), .B1(new_n1223), .B2(new_n1228), .ZN(G375));
  NAND2_X1  g1029(.A1(new_n914), .A2(new_n758), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n819), .B1(G68), .B2(new_n831), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n839), .A2(new_n836), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n258), .B1(new_n780), .B2(new_n226), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(G283), .B2(new_n799), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n805), .A2(G97), .B1(new_n787), .B2(G77), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n488), .A2(new_n793), .B1(new_n795), .B2(G294), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1027), .A2(new_n1234), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1026), .A2(G50), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n849), .A2(new_n796), .B1(new_n794), .B2(new_n1118), .ZN(new_n1239));
  AOI211_X1 g1039(.A(new_n1172), .B(new_n1239), .C1(G159), .C2(new_n805), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n799), .A2(G137), .B1(new_n1028), .B2(G150), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1238), .A2(new_n1240), .A3(new_n455), .A4(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(new_n772), .A2(G128), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n1232), .A2(new_n1237), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1231), .B1(new_n1244), .B2(new_n761), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1147), .A2(new_n747), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1153), .B1(new_n1141), .B2(new_n1138), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n963), .B(KEYINPUT123), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1248), .B2(new_n1249), .ZN(G381));
  OR4_X1    g1050(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1251), .A2(G387), .A3(G381), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1127), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1156), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1168), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(G375), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1252), .A2(new_n1256), .A3(new_n1257), .ZN(G407));
  NOR2_X1   g1058(.A1(new_n677), .A2(G343), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1260), .A2(KEYINPUT124), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(KEYINPUT124), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G213), .B(G407), .C1(new_n1261), .C2(new_n1262), .ZN(G409));
  INV_X1    g1063(.A(G390), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(G396), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(G393), .B(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n985), .A2(new_n1012), .A3(G390), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1267), .A2(new_n1269), .B1(new_n1265), .B2(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1265), .A2(KEYINPUT126), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1217), .C1(new_n1223), .C2(new_n1228), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1202), .B1(new_n1277), .B2(new_n747), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1215), .B(new_n1211), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1278), .B1(new_n1279), .B2(new_n1249), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1256), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1259), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT60), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n702), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1287), .B1(new_n1247), .B2(new_n1286), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1246), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  AND2_X1   g1091(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1289), .B1(new_n1292), .B2(new_n1290), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1259), .A2(G2897), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1294), .B(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1284), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1294), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1282), .A2(new_n1283), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT62), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1259), .B1(new_n1276), .B2(new_n1281), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT62), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(new_n1300), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1275), .B1(new_n1299), .B2(new_n1306), .ZN(new_n1307));
  AND3_X1   g1107(.A1(new_n1303), .A2(KEYINPUT63), .A3(new_n1300), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT63), .B1(new_n1303), .B2(new_n1300), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1274), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT127), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1295), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1294), .B(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(new_n1312), .B(new_n1298), .C1(new_n1303), .C2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1307), .A2(new_n1317), .ZN(G405));
  NAND2_X1  g1118(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1294), .B1(new_n1321), .B2(new_n1272), .ZN(new_n1322));
  NOR3_X1   g1122(.A1(new_n1271), .A2(new_n1273), .A3(new_n1300), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(G375), .B(G378), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(new_n1324), .B(new_n1325), .ZN(G402));
endmodule


