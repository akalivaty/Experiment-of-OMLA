//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1276, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT0), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT65), .Z(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G58), .ZN(new_n215));
  INV_X1    g0015(.A(G232), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT67), .B(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n221), .A2(G77), .B1(G68), .B2(G238), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n219), .B2(KEYINPUT68), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n204), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n207), .B1(new_n211), .B2(new_n213), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n216), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n231), .B(new_n232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT69), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n233), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G58), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT70), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT71), .ZN(new_n241));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G351));
  NOR2_X1   g0048(.A1(KEYINPUT78), .A2(KEYINPUT10), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT8), .B(G58), .Z(new_n250));
  INV_X1    g0050(.A(KEYINPUT74), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n251), .B1(new_n252), .B2(G20), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n209), .A2(KEYINPUT74), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  NOR3_X1   g0056(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n257));
  INV_X1    g0057(.A(G150), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n256), .B1(new_n209), .B2(new_n257), .C1(new_n258), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n208), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  INV_X1    g0068(.A(G50), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n265), .B2(G20), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n268), .A2(new_n270), .B1(new_n269), .B2(new_n267), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  AND2_X1   g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n275), .A2(KEYINPUT73), .A3(new_n208), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT73), .ZN(new_n277));
  AND2_X1   g0077(.A1(G1), .A2(G13), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G41), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G222), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G223), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n281), .B(new_n288), .C1(G77), .C2(new_n284), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n265), .A2(new_n292), .B1(new_n278), .B2(new_n279), .ZN(new_n293));
  OR2_X1    g0093(.A1(KEYINPUT72), .A2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(KEYINPUT72), .A2(G45), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G274), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G1), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n293), .A2(G226), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G190), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n300), .A2(G200), .B1(KEYINPUT78), .B2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n249), .B1(new_n274), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n272), .B(KEYINPUT9), .ZN(new_n306));
  INV_X1    g0106(.A(new_n249), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n306), .A2(new_n307), .A3(new_n302), .A4(new_n303), .ZN(new_n308));
  INV_X1    g0108(.A(new_n272), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n310), .B2(new_n300), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(G179), .B2(new_n300), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n305), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n284), .A2(G232), .A3(new_n286), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n284), .A2(G238), .A3(G1698), .ZN(new_n315));
  AND2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G107), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n315), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(new_n281), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n293), .A2(new_n221), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n296), .A2(new_n298), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n310), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n324), .B1(new_n281), .B2(new_n320), .ZN(new_n328));
  INV_X1    g0128(.A(G179), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT76), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n266), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n265), .A2(KEYINPUT76), .A3(G13), .A4(G20), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G77), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n263), .B1(new_n332), .B2(new_n333), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n265), .B2(G20), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n335), .A2(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(KEYINPUT8), .B(G58), .ZN(new_n340));
  OAI22_X1  g0140(.A1(new_n340), .A2(new_n260), .B1(new_n209), .B2(new_n336), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT15), .B(G87), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT75), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n341), .B1(new_n344), .B2(new_n255), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n262), .A2(new_n208), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n327), .A2(new_n330), .A3(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n313), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(G68), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT7), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(new_n284), .B2(G20), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n318), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n215), .A2(new_n351), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G58), .A2(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(G20), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n259), .A2(G159), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n350), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(KEYINPUT7), .B1(new_n318), .B2(new_n209), .ZN(new_n362));
  NOR4_X1   g0162(.A1(new_n316), .A2(new_n317), .A3(new_n352), .A4(G20), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(new_n360), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(KEYINPUT16), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n361), .A2(new_n263), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n265), .A2(G20), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n250), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n346), .A2(new_n266), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n369), .A2(new_n370), .B1(new_n266), .B2(new_n250), .ZN(new_n371));
  XNOR2_X1  g0171(.A(new_n371), .B(KEYINPUT80), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  OR2_X1    g0173(.A1(G223), .A2(G1698), .ZN(new_n374));
  INV_X1    g0174(.A(G226), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G1698), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n376), .C1(new_n316), .C2(new_n317), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n281), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n293), .A2(G232), .B1(new_n296), .B2(new_n298), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(KEYINPUT81), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT81), .B1(new_n380), .B2(new_n381), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n310), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n381), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n329), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n373), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT18), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT81), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n382), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(new_n310), .B1(new_n329), .B2(new_n387), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT18), .A3(new_n373), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(KEYINPUT82), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(G200), .B1(new_n393), .B2(new_n382), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n386), .A2(G190), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n367), .B(new_n372), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n383), .B2(new_n384), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(G190), .B2(new_n386), .ZN(new_n405));
  INV_X1    g0205(.A(new_n373), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT17), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT82), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n395), .A2(new_n408), .A3(KEYINPUT18), .A4(new_n373), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n402), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n326), .A2(G200), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT77), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT15), .B(G87), .Z(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n343), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n342), .A2(KEYINPUT75), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(new_n255), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n341), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n263), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n411), .A2(new_n412), .A3(new_n419), .A4(new_n339), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n403), .B1(new_n321), .B2(new_n325), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT77), .B1(new_n347), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n328), .A2(G190), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n349), .A2(new_n397), .A3(new_n410), .A4(new_n424), .ZN(new_n425));
  OAI211_X1 g0225(.A(G226), .B(new_n286), .C1(new_n316), .C2(new_n317), .ZN(new_n426));
  OAI211_X1 g0226(.A(G232), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n427));
  INV_X1    g0227(.A(G97), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n426), .B(new_n427), .C1(new_n252), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n281), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n293), .A2(G238), .B1(new_n296), .B2(new_n298), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n430), .A2(new_n434), .A3(new_n431), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(KEYINPUT79), .A3(new_n435), .ZN(new_n436));
  OR3_X1    g0236(.A1(new_n432), .A2(KEYINPUT79), .A3(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(G169), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT14), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n436), .A2(new_n437), .A3(new_n440), .A4(G169), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n433), .A2(G179), .A3(new_n435), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n255), .A2(G77), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n259), .A2(G50), .B1(G20), .B2(new_n351), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n346), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n337), .A2(G68), .A3(new_n368), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT12), .B1(new_n334), .B2(G68), .ZN(new_n450));
  INV_X1    g0250(.A(G13), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT12), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(G20), .A4(new_n351), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n447), .A2(new_n448), .A3(new_n449), .A4(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n443), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n436), .A2(new_n437), .A3(G200), .ZN(new_n458));
  INV_X1    g0258(.A(G190), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n432), .B2(KEYINPUT13), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n456), .B1(new_n460), .B2(new_n435), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n425), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT85), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT21), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n291), .A2(G1), .ZN(new_n467));
  AND2_X1   g0267(.A1(KEYINPUT5), .A2(G41), .ZN(new_n468));
  NOR2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n278), .A2(new_n279), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(G270), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n297), .B1(new_n278), .B2(new_n279), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(new_n467), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(G257), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n286), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n218), .A2(G1698), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n478), .B(new_n479), .C1(new_n316), .C2(new_n317), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n281), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT84), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT84), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n281), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n476), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n265), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n334), .A2(G116), .A3(new_n346), .A4(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G116), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n332), .A2(new_n490), .A3(new_n333), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n262), .A2(new_n208), .B1(G20), .B2(new_n490), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n494), .B(new_n209), .C1(G33), .C2(new_n428), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n493), .A2(KEYINPUT20), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(KEYINPUT20), .B1(new_n493), .B2(new_n495), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(G169), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n466), .B1(new_n487), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n476), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n281), .A2(new_n482), .A3(new_n485), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n485), .B1(new_n281), .B2(new_n482), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n489), .B(new_n491), .C1(new_n497), .C2(new_n496), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n504), .A2(KEYINPUT21), .A3(G169), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n472), .A2(new_n475), .A3(G179), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n484), .B2(new_n486), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n505), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n500), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(G190), .B(new_n501), .C1(new_n502), .C2(new_n503), .ZN(new_n511));
  INV_X1    g0311(.A(new_n505), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n487), .C2(new_n403), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n465), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n504), .A2(G169), .A3(new_n505), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(new_n466), .B1(new_n505), .B2(new_n508), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n517), .A2(KEYINPUT85), .A3(new_n506), .A4(new_n513), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n209), .B(G87), .C1(new_n316), .C2(new_n317), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT22), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n284), .A2(new_n522), .A3(new_n209), .A4(G87), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G20), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n209), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n217), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(G20), .B1(new_n282), .B2(new_n283), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n522), .B1(new_n535), .B2(G87), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n520), .A2(KEYINPUT22), .ZN(new_n537));
  OAI211_X1 g0337(.A(KEYINPUT86), .B(new_n530), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT86), .B1(new_n524), .B2(new_n530), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n534), .B(new_n263), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n267), .A2(new_n217), .ZN(new_n542));
  XNOR2_X1  g0342(.A(new_n542), .B(KEYINPUT25), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n268), .A2(new_n488), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(new_n217), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n286), .C1(new_n316), .C2(new_n317), .ZN(new_n547));
  OAI211_X1 g0347(.A(G257), .B(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n548));
  AND2_X1   g0348(.A1(KEYINPUT87), .A2(G294), .ZN(new_n549));
  NOR2_X1   g0349(.A1(KEYINPUT87), .A2(G294), .ZN(new_n550));
  OAI21_X1  g0350(.A(G33), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n281), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n275), .A2(new_n208), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n467), .B2(new_n474), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G264), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n556), .A3(new_n475), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n403), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n553), .A2(new_n556), .A3(new_n459), .A4(new_n475), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n541), .A2(new_n546), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT88), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n557), .A2(new_n562), .A3(G169), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n553), .A2(new_n556), .A3(G179), .A4(new_n475), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n557), .B2(G169), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n546), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n531), .A2(new_n532), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n569), .A2(KEYINPUT24), .A3(new_n538), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n346), .B1(new_n540), .B2(new_n533), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n561), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n266), .A2(G97), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n544), .B2(new_n428), .ZN(new_n576));
  OAI21_X1  g0376(.A(G107), .B1(new_n362), .B2(new_n363), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  AND2_X1   g0378(.A1(G97), .A2(G107), .ZN(new_n579));
  NOR2_X1   g0379(.A1(G97), .A2(G107), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n583), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n576), .B1(new_n585), .B2(new_n263), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT4), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n587), .A2(G1698), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n588), .B(G244), .C1(new_n317), .C2(new_n316), .ZN(new_n589));
  INV_X1    g0389(.A(G244), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n282), .B2(new_n283), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n589), .B(new_n494), .C1(new_n591), .C2(KEYINPUT4), .ZN(new_n592));
  OAI21_X1  g0392(.A(G250), .B1(new_n316), .B2(new_n317), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n286), .B1(new_n593), .B2(KEYINPUT4), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n281), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n470), .A2(new_n471), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n475), .B1(new_n596), .B2(new_n477), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n598), .A3(G190), .ZN(new_n599));
  OAI21_X1  g0399(.A(G244), .B1(new_n316), .B2(new_n317), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n587), .B1(G33), .B2(G283), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n587), .B1(new_n284), .B2(G250), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n589), .C1(new_n286), .C2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n597), .B1(new_n603), .B2(new_n281), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n586), .B(new_n599), .C1(new_n403), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n595), .A2(new_n598), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n310), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n583), .A2(G20), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n259), .A2(G77), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n217), .B1(new_n353), .B2(new_n354), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n263), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n576), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n595), .A2(new_n598), .A3(new_n329), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(G87), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n580), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT19), .ZN(new_n619));
  NOR3_X1   g0419(.A1(new_n619), .A2(new_n252), .A3(new_n428), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n618), .B1(new_n620), .B2(G20), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n535), .A2(G68), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n428), .B1(new_n253), .B2(new_n254), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n621), .B(new_n622), .C1(KEYINPUT19), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n263), .ZN(new_n625));
  INV_X1    g0425(.A(new_n544), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n344), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n414), .A2(new_n415), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n335), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n625), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(G250), .B1(new_n291), .B2(G1), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT83), .B1(new_n554), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT83), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n265), .A2(G45), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n471), .A2(new_n633), .A3(G250), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n473), .A2(new_n467), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n590), .A2(G1698), .ZN(new_n638));
  OAI221_X1 g0438(.A(new_n638), .B1(G238), .B2(G1698), .C1(new_n316), .C2(new_n317), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n525), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n281), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n310), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT73), .B1(new_n275), .B2(new_n208), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n278), .A2(new_n277), .A3(new_n279), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n525), .B2(new_n639), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n632), .A2(new_n635), .A3(new_n636), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n329), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n630), .A2(new_n643), .A3(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n624), .A2(new_n263), .B1(new_n628), .B2(new_n335), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n637), .A2(new_n641), .A3(G190), .ZN(new_n653));
  OAI21_X1  g0453(.A(G200), .B1(new_n647), .B2(new_n648), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n626), .A2(G87), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n605), .A2(new_n616), .A3(new_n651), .A4(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n573), .A2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n464), .A2(new_n519), .A3(new_n658), .ZN(G372));
  AND2_X1   g0459(.A1(new_n651), .A2(new_n656), .ZN(new_n660));
  INV_X1    g0460(.A(new_n616), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(KEYINPUT26), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT26), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n651), .A2(new_n656), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(new_n664), .B2(new_n616), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n605), .A2(new_n616), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n561), .A3(new_n660), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n567), .A2(new_n572), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n510), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n666), .B(new_n651), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n464), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n312), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n391), .A2(new_n396), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n443), .A2(new_n456), .B1(new_n462), .B2(new_n348), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n402), .A2(new_n407), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n305), .A2(new_n308), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(G369));
  NAND2_X1  g0480(.A1(new_n452), .A2(new_n209), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n572), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT90), .ZN(new_n689));
  INV_X1    g0489(.A(new_n573), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n669), .A2(new_n686), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT89), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n686), .A2(new_n505), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n519), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n510), .A2(new_n505), .A3(new_n686), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n695), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n698), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT89), .A3(G330), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n694), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n510), .A2(new_n687), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n689), .A2(new_n690), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n669), .A2(new_n687), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n704), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n205), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  NOR4_X1   g0512(.A1(new_n712), .A2(new_n265), .A3(G116), .A4(new_n618), .ZN(new_n713));
  INV_X1    g0513(.A(new_n212), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n712), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT28), .Z(new_n716));
  NAND2_X1  g0516(.A1(new_n671), .A2(new_n687), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n651), .B1(new_n670), .B2(new_n668), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n662), .A2(new_n665), .A3(KEYINPUT93), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT93), .ZN(new_n722));
  OAI211_X1 g0522(.A(new_n722), .B(new_n663), .C1(new_n664), .C2(new_n616), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g0524(.A(KEYINPUT29), .B(new_n687), .C1(new_n720), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n507), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n502), .B2(new_n503), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n553), .A2(new_n556), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n728), .A2(new_n729), .A3(new_n642), .ZN(new_n730));
  AOI21_X1  g0530(.A(KEYINPUT30), .B1(new_n730), .B2(new_n604), .ZN(new_n731));
  AOI21_X1  g0531(.A(G179), .B1(new_n637), .B2(new_n641), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n504), .A2(new_n606), .A3(new_n732), .A4(new_n557), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n484), .A2(new_n486), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n553), .A2(new_n556), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(new_n735), .A3(new_n727), .A4(new_n649), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n604), .A2(KEYINPUT30), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT91), .B1(new_n731), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n736), .A2(new_n737), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n736), .B2(new_n606), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT91), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n740), .A2(new_n742), .A3(new_n743), .A4(new_n733), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n686), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT31), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n519), .A2(new_n658), .A3(new_n687), .ZN(new_n748));
  OAI211_X1 g0548(.A(KEYINPUT31), .B(new_n686), .C1(new_n731), .C2(new_n738), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  AND2_X1   g0551(.A1(new_n726), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n716), .B1(new_n752), .B2(G1), .ZN(G364));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n208), .B1(G20), .B2(new_n310), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n711), .A2(new_n284), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n294), .A2(new_n295), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n760), .B1(new_n213), .B2(new_n761), .C1(new_n243), .C2(new_n291), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n284), .A2(G355), .ZN(new_n763));
  MUX2_X1   g0563(.A(G116), .B(new_n763), .S(new_n205), .Z(new_n764));
  AOI21_X1  g0564(.A(new_n759), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n757), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n209), .A2(new_n459), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n329), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n209), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G58), .A2(new_n770), .B1(new_n773), .B2(G77), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n209), .A2(new_n329), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n774), .B1(new_n269), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT95), .Z(new_n778));
  INV_X1    g0578(.A(new_n771), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n329), .A2(new_n403), .A3(KEYINPUT96), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT96), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G179), .B2(G200), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n779), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G159), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n784), .A2(KEYINPUT32), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n459), .B1(new_n780), .B2(new_n782), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n209), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G97), .A2(new_n788), .B1(new_n784), .B2(KEYINPUT32), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n403), .A2(G179), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n771), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n767), .A2(new_n790), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n284), .B1(new_n791), .B2(new_n217), .C1(new_n617), .C2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n775), .A2(new_n459), .A3(G200), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(KEYINPUT97), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n793), .B1(new_n798), .B2(G68), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n778), .A2(new_n785), .A3(new_n789), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n769), .A2(new_n801), .B1(new_n772), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G303), .ZN(new_n804));
  INV_X1    g0604(.A(G326), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n318), .B1(new_n792), .B2(new_n804), .C1(new_n805), .C2(new_n776), .ZN(new_n806));
  INV_X1    g0606(.A(new_n791), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n803), .B(new_n806), .C1(G283), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n783), .A2(G329), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n549), .A2(new_n550), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n788), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n798), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n808), .A2(new_n809), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n766), .B1(new_n800), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n451), .A2(G20), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n265), .B1(new_n816), .B2(G45), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n712), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n765), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n756), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n702), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n702), .A2(G330), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT94), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n701), .A2(new_n703), .A3(new_n820), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT98), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n347), .A2(new_n686), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n348), .B1(new_n424), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n348), .A2(new_n687), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(KEYINPUT100), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n419), .B(new_n339), .C1(new_n328), .C2(new_n403), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n835), .A2(KEYINPUT77), .B1(G190), .B2(new_n328), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n836), .A2(new_n420), .B1(new_n347), .B2(new_n686), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(new_n831), .C1(new_n837), .C2(new_n348), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n717), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(new_n671), .A3(new_n687), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n819), .B1(new_n843), .B2(new_n751), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n751), .B2(new_n843), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n757), .A2(new_n754), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT99), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n819), .B1(G77), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(G294), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n769), .A2(new_n849), .B1(new_n772), .B2(new_n490), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n318), .B1(new_n791), .B2(new_n617), .C1(new_n776), .C2(new_n804), .ZN(new_n851));
  INV_X1    g0651(.A(new_n792), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n850), .B(new_n851), .C1(G107), .C2(new_n852), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n798), .A2(G283), .B1(G97), .B2(new_n788), .ZN(new_n854));
  INV_X1    g0654(.A(new_n783), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n853), .B(new_n854), .C1(new_n802), .C2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n770), .B1(new_n773), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n858), .B2(new_n776), .C1(new_n797), .C2(new_n258), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n284), .B1(new_n791), .B2(new_n351), .C1(new_n269), .C2(new_n792), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G132), .B2(new_n783), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n215), .C2(new_n787), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n859), .A2(new_n860), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n856), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n848), .B1(new_n866), .B2(new_n757), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n867), .B1(new_n839), .B2(new_n755), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n845), .A2(new_n868), .ZN(G384));
  XOR2_X1   g0669(.A(new_n583), .B(KEYINPUT101), .Z(new_n870));
  INV_X1    g0670(.A(KEYINPUT35), .ZN(new_n871));
  OAI211_X1 g0671(.A(G116), .B(new_n210), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT36), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n714), .B(G77), .C1(new_n215), .C2(new_n351), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n269), .A2(G68), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n265), .B(G13), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n816), .A2(new_n265), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n391), .A2(new_n396), .A3(new_n684), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  INV_X1    g0681(.A(new_n684), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n373), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n676), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n674), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n389), .A2(new_n400), .A3(new_n883), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n886), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n881), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT103), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT16), .B1(new_n364), .B2(new_n365), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n891), .B2(new_n346), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n361), .A2(KEYINPUT103), .A3(new_n263), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n366), .ZN(new_n894));
  INV_X1    g0694(.A(new_n371), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n684), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n391), .A2(KEYINPUT82), .A3(new_n396), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n402), .A2(new_n407), .A3(new_n409), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n389), .A2(new_n400), .A3(new_n887), .A4(new_n883), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n385), .A2(new_n388), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n895), .B2(new_n894), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n399), .B1(new_n394), .B2(new_n403), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n903), .A2(new_n373), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n902), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n900), .B1(new_n905), .B2(new_n887), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n899), .A2(new_n906), .A3(KEYINPUT38), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n889), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n894), .A2(new_n895), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n882), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n410), .B2(new_n397), .ZN(new_n913));
  AND4_X1   g0713(.A1(new_n887), .A2(new_n389), .A3(new_n400), .A4(new_n883), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n395), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n912), .A2(new_n915), .A3(new_n400), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n914), .B1(new_n916), .B2(KEYINPUT37), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n881), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n907), .A3(KEYINPUT39), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n457), .A2(new_n686), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n880), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(new_n907), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n456), .A2(new_n686), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n457), .A2(new_n462), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n462), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n456), .B(new_n686), .C1(new_n443), .C2(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n842), .A2(new_n831), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT102), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n651), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n657), .B1(new_n572), .B2(new_n560), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n570), .A2(new_n571), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n934), .A2(new_n568), .B1(new_n566), .B2(new_n565), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(new_n506), .A3(new_n517), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n932), .B1(new_n933), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n686), .B1(new_n937), .B2(new_n666), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n832), .B1(new_n938), .B2(new_n839), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n926), .A2(new_n928), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NOR3_X1   g0741(.A1(new_n939), .A2(KEYINPUT102), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n931), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n923), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n464), .A2(new_n725), .A3(new_n719), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n679), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n889), .A2(new_n907), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n739), .A2(new_n744), .A3(KEYINPUT31), .A4(new_n686), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n747), .A2(new_n748), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n940), .A2(new_n950), .A3(new_n839), .ZN(new_n951));
  OAI21_X1  g0751(.A(KEYINPUT40), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT40), .B1(new_n918), .B2(new_n907), .ZN(new_n953));
  AND3_X1   g0753(.A1(new_n940), .A2(new_n950), .A3(new_n839), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n464), .A2(new_n950), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n958), .A2(new_n959), .A3(new_n700), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n879), .B1(new_n947), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT104), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n961), .A2(new_n962), .B1(new_n947), .B2(new_n960), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n878), .B1(new_n963), .B2(new_n964), .ZN(G367));
  INV_X1    g0765(.A(new_n760), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n966), .A2(new_n237), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n759), .B1(new_n711), .B2(new_n344), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n820), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n652), .A2(new_n655), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n686), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n660), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n971), .A2(new_n651), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n798), .A2(new_n810), .B1(G107), .B2(new_n788), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n318), .B1(new_n791), .B2(new_n428), .ZN(new_n977));
  INV_X1    g0777(.A(G283), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n769), .A2(new_n804), .B1(new_n772), .B2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(G317), .C2(new_n783), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n792), .A2(new_n490), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n981), .A2(KEYINPUT46), .ZN(new_n982));
  INV_X1    g0782(.A(new_n776), .ZN(new_n983));
  AOI22_X1  g0783(.A1(KEYINPUT46), .A2(new_n981), .B1(new_n983), .B2(G311), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n976), .A2(new_n980), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n284), .B1(new_n769), .B2(new_n258), .ZN(new_n986));
  AOI22_X1  g0786(.A1(G58), .A2(new_n852), .B1(new_n773), .B2(G50), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n336), .B2(new_n791), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n986), .B(new_n988), .C1(G143), .C2(new_n983), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n858), .B2(new_n855), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n788), .A2(G68), .ZN(new_n991));
  INV_X1    g0791(.A(G159), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n991), .B1(new_n992), .B2(new_n797), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n985), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  OAI221_X1 g0795(.A(new_n969), .B1(new_n822), .B2(new_n975), .C1(new_n995), .C2(new_n766), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n667), .B1(new_n586), .B2(new_n687), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n661), .A2(new_n686), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n997), .B1(new_n709), .B2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n707), .A2(KEYINPUT45), .A3(new_n708), .A4(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1000), .B1(new_n707), .B2(new_n708), .ZN(new_n1005));
  XOR2_X1   g0805(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1004), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n704), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n701), .A2(new_n703), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n693), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1012), .A2(new_n1004), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n707), .B1(new_n693), .B2(new_n706), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT108), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1015), .A2(new_n701), .A3(KEYINPUT108), .A4(new_n703), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n752), .B1(new_n1014), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n712), .B(KEYINPUT41), .Z(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n818), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g0824(.A1(new_n707), .A2(new_n1001), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1025), .A2(KEYINPUT42), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n616), .B1(new_n998), .B2(new_n935), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1025), .A2(KEYINPUT42), .B1(new_n687), .B2(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1026), .A2(new_n1028), .B1(KEYINPUT43), .B2(new_n975), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n974), .A2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT106), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1034), .A2(new_n704), .A3(new_n1000), .A4(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n975), .A2(KEYINPUT43), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n1037), .A2(new_n1032), .A3(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1033), .A2(new_n1039), .B1(new_n1012), .B2(new_n1001), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n996), .B1(new_n1024), .B2(new_n1041), .ZN(G387));
  NAND3_X1  g0842(.A1(new_n1018), .A2(new_n752), .A3(new_n1019), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n712), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(KEYINPUT109), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT109), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1046), .A3(new_n712), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n752), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1020), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n694), .A2(new_n756), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n233), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(new_n318), .A3(new_n761), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n618), .A2(G116), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n291), .B1(new_n351), .B2(new_n336), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n250), .A2(KEYINPUT50), .A3(new_n269), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT50), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n340), .B2(G50), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1055), .B1(new_n1060), .B2(new_n284), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n711), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n758), .B1(new_n205), .B2(new_n217), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n819), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n792), .A2(new_n336), .B1(new_n772), .B2(new_n351), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n284), .B1(new_n791), .B2(new_n428), .C1(new_n776), .C2(new_n992), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n770), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n783), .A2(G150), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n788), .A2(new_n344), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n798), .A2(new_n250), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(G317), .A2(new_n770), .B1(new_n773), .B2(G303), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n801), .B2(new_n776), .C1(new_n797), .C2(new_n802), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n788), .A2(G283), .B1(new_n810), .B2(new_n852), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT49), .Z(new_n1079));
  OAI221_X1 g0879(.A(new_n318), .B1(new_n490), .B2(new_n791), .C1(new_n855), .C2(new_n805), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1071), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1064), .B1(new_n1081), .B2(new_n757), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1051), .A2(new_n818), .B1(new_n1052), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1050), .A2(new_n1083), .ZN(G393));
  NOR2_X1   g0884(.A1(new_n966), .A2(new_n247), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n758), .B1(new_n205), .B2(new_n428), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n819), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n798), .A2(G50), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n284), .B1(new_n791), .B2(new_n617), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n792), .A2(new_n351), .B1(new_n772), .B2(new_n340), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G143), .C2(new_n783), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n776), .A2(new_n258), .B1(new_n769), .B2(new_n992), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT51), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n788), .A2(G77), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1088), .A2(new_n1091), .A3(new_n1093), .A4(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n318), .B1(new_n791), .B2(new_n217), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n792), .A2(new_n978), .B1(new_n772), .B2(new_n849), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(G322), .C2(new_n783), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n490), .B2(new_n787), .C1(new_n804), .C2(new_n797), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n983), .A2(G317), .B1(new_n770), .B2(G311), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT110), .B(KEYINPUT52), .Z(new_n1101));
  XNOR2_X1  g0901(.A(new_n1100), .B(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1095), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1087), .B1(new_n1103), .B2(new_n757), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1000), .B2(new_n822), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1051), .A2(new_n752), .A3(new_n1013), .A4(new_n1010), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n712), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n1014), .A2(new_n1043), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1105), .B1(new_n817), .B2(new_n1014), .C1(new_n1107), .C2(new_n1108), .ZN(G390));
  AND2_X1   g0909(.A1(new_n950), .A2(new_n839), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1110), .A2(KEYINPUT111), .A3(G330), .A4(new_n940), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n940), .A2(new_n950), .A3(G330), .A4(new_n839), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT111), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n941), .B1(new_n751), .B2(new_n840), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n939), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n687), .B1(new_n720), .B2(new_n724), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n831), .B1(new_n1119), .B2(new_n840), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n751), .A2(new_n840), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n940), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT112), .ZN(new_n1123));
  AND3_X1   g0923(.A1(new_n950), .A2(new_n1123), .A3(G330), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n950), .B2(G330), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1124), .A2(new_n1125), .A3(new_n840), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1122), .B1(new_n1126), .B2(new_n940), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1118), .A2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n918), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT39), .B1(new_n889), .B2(new_n907), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1129), .A2(new_n1130), .B1(new_n929), .B2(new_n921), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1120), .A2(new_n940), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n921), .B1(new_n889), .B2(new_n907), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n950), .A2(G330), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n464), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n945), .A2(new_n679), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1121), .A2(new_n940), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1131), .A2(new_n1143), .A3(new_n1134), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1128), .A2(new_n1137), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1145), .A2(new_n712), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1128), .A2(new_n1142), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n922), .B1(new_n939), .B2(new_n941), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n920), .A2(new_n1148), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1136), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1144), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1147), .A2(KEYINPUT113), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT113), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1146), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1137), .A2(new_n818), .A3(new_n1144), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n819), .B1(new_n250), .B2(new_n847), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n852), .A2(G150), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1158), .A2(KEYINPUT53), .B1(new_n1159), .B2(new_n776), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(KEYINPUT53), .B2(new_n1158), .ZN(new_n1161));
  INV_X1    g0961(.A(G132), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n769), .A2(new_n1162), .B1(new_n791), .B2(new_n269), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(KEYINPUT54), .B(G143), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n318), .B(new_n1163), .C1(new_n773), .C2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(G125), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1161), .B(new_n1166), .C1(new_n1167), .C2(new_n855), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n797), .A2(new_n858), .B1(new_n992), .B2(new_n787), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n798), .A2(G107), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n769), .A2(new_n490), .B1(new_n772), .B2(new_n428), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n284), .B(new_n1171), .C1(G87), .C2(new_n852), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n983), .A2(G283), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1172), .A3(new_n1094), .A4(new_n1173), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n783), .A2(G294), .B1(new_n807), .B2(G68), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT114), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1168), .A2(new_n1169), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1157), .B1(new_n1177), .B2(new_n757), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n920), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n755), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1156), .A2(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1155), .A2(new_n1181), .ZN(G378));
  NOR2_X1   g0982(.A1(new_n309), .A2(new_n684), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n313), .B(new_n1183), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1184), .B(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n956), .B2(G330), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n700), .B(new_n1186), .C1(new_n952), .C2(new_n955), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n1188), .A2(new_n1189), .B1(new_n943), .B2(new_n923), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n954), .A2(new_n908), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(KEYINPUT40), .B1(new_n954), .B2(new_n953), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1186), .B1(new_n1192), .B2(new_n700), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n956), .A2(G330), .A3(new_n1187), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n944), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n818), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n820), .B1(new_n269), .B2(new_n846), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n318), .A2(new_n290), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G77), .B2(new_n852), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n215), .B2(new_n791), .C1(new_n978), .C2(new_n855), .ZN(new_n1201));
  XOR2_X1   g1001(.A(new_n1201), .B(KEYINPUT115), .Z(new_n1202));
  NAND2_X1  g1002(.A1(new_n344), .A2(new_n773), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n983), .A2(G116), .B1(new_n770), .B2(G107), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n991), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1202), .B(new_n1205), .C1(new_n428), .C2(new_n797), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1199), .B(new_n269), .C1(G33), .C2(G41), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n252), .B(new_n290), .C1(new_n791), .C2(new_n992), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n787), .A2(new_n258), .B1(new_n1167), .B2(new_n776), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT117), .Z(new_n1214));
  AOI22_X1  g1014(.A1(new_n798), .A2(G132), .B1(G137), .B2(new_n773), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n1159), .A2(new_n769), .B1(new_n792), .B2(new_n1164), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT116), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1217), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1212), .B(new_n1219), .C1(G124), .C2(new_n783), .ZN(new_n1220));
  OR2_X1    g1020(.A1(new_n1218), .A2(KEYINPUT59), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1208), .B(new_n1211), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1198), .B1(new_n766), .B2(new_n1222), .C1(new_n1187), .C2(new_n755), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT118), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1145), .B2(new_n1142), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1138), .A2(KEYINPUT112), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n950), .A2(new_n1123), .A3(G330), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1227), .A2(new_n839), .A3(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n941), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1117), .A2(new_n1116), .B1(new_n1230), .B2(new_n1122), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1225), .B(new_n1142), .C1(new_n1151), .C2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1226), .A2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1190), .A2(new_n1195), .A3(KEYINPUT119), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT119), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n944), .A2(new_n1193), .A3(new_n1236), .A4(new_n1194), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(KEYINPUT57), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n712), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1142), .B1(new_n1151), .B2(new_n1231), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(KEYINPUT118), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1232), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT57), .B1(new_n1242), .B2(new_n1196), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1224), .B1(new_n1239), .B2(new_n1243), .ZN(G375));
  NAND3_X1  g1044(.A1(new_n1118), .A2(new_n1127), .A3(new_n1141), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1147), .A2(new_n1023), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n941), .A2(new_n754), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n819), .B1(G68), .B2(new_n847), .ZN(new_n1248));
  OAI221_X1 g1048(.A(new_n318), .B1(new_n791), .B2(new_n336), .C1(new_n776), .C2(new_n849), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G97), .A2(new_n852), .B1(new_n770), .B2(G283), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n217), .B2(new_n772), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1249), .B(new_n1251), .C1(G303), .C2(new_n783), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n1069), .C1(new_n490), .C2(new_n797), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n776), .A2(new_n1162), .B1(new_n769), .B2(new_n858), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(new_n798), .B2(new_n1165), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1255), .B(KEYINPUT120), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n284), .B1(new_n791), .B2(new_n215), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n792), .A2(new_n992), .B1(new_n772), .B2(new_n258), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(G128), .C2(new_n783), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n269), .B2(new_n787), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1253), .B1(new_n1256), .B2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1248), .B1(new_n1261), .B2(new_n757), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT121), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1247), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1231), .B2(new_n817), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1246), .A2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(G375), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1155), .A2(new_n1181), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1270));
  INV_X1    g1070(.A(G396), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1050), .A2(new_n1271), .A3(new_n1083), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(G384), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT122), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1274), .ZN(G407));
  NAND2_X1  g1075(.A1(new_n685), .A2(G213), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1268), .A2(new_n1269), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(G213), .A3(new_n1278), .ZN(G409));
  NAND2_X1  g1079(.A1(G393), .A2(G396), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(G387), .A2(new_n1280), .A3(new_n1272), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1022), .B1(new_n1106), .B2(new_n752), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1036), .B(new_n1040), .C1(new_n1282), .C2(new_n818), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT125), .B1(new_n1283), .B2(new_n996), .ZN(new_n1284));
  AND3_X1   g1084(.A1(new_n1050), .A2(new_n1271), .A3(new_n1083), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1271), .B1(new_n1050), .B2(new_n1083), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1281), .B(G390), .C1(new_n1284), .C2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1280), .A2(new_n1272), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(G390), .B1(new_n1293), .B2(new_n1281), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1224), .C1(new_n1239), .C2(new_n1243), .ZN(new_n1296));
  AND3_X1   g1096(.A1(new_n1242), .A2(new_n1023), .A3(new_n1196), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1235), .A2(new_n818), .A3(new_n1237), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1223), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1269), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1296), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1276), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1277), .A2(G2897), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G384), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1245), .A2(KEYINPUT60), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT60), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1118), .A2(new_n1127), .A3(new_n1307), .A4(new_n1141), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n712), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1310), .B1(new_n1128), .B2(new_n1142), .ZN(new_n1311));
  AOI211_X1 g1111(.A(new_n1305), .B(new_n1265), .C1(new_n1309), .C2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1307), .B1(new_n1231), .B2(new_n1141), .ZN(new_n1313));
  AND4_X1   g1113(.A1(new_n1307), .A2(new_n1118), .A3(new_n1141), .A4(new_n1127), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1311), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1315), .B2(new_n1266), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1312), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT124), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1304), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n712), .B1(new_n1231), .B2(new_n1141), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1320), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1305), .B1(new_n1321), .B2(new_n1265), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1315), .A2(G384), .A3(new_n1266), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT124), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1319), .A2(new_n1325), .ZN(new_n1326));
  AND4_X1   g1126(.A1(new_n1318), .A2(new_n1322), .A3(new_n1323), .A4(new_n1304), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  AOI21_X1  g1129(.A(KEYINPUT61), .B1(new_n1302), .B2(new_n1329), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1301), .A2(new_n1276), .A3(new_n1317), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1332), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1331), .A2(KEYINPUT62), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1295), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1317), .A2(KEYINPUT63), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1301), .A2(new_n1276), .A3(new_n1337), .ZN(new_n1338));
  OR2_X1    g1138(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT61), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1277), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1327), .B1(new_n1319), .B2(new_n1325), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1341), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1340), .A2(new_n1344), .ZN(new_n1345));
  XOR2_X1   g1145(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1346));
  NAND2_X1  g1146(.A1(new_n1331), .A2(new_n1346), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1336), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1295), .B1(new_n1342), .B2(new_n1337), .ZN(new_n1349));
  AND4_X1   g1149(.A1(new_n1336), .A2(new_n1330), .A3(new_n1349), .A4(new_n1347), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1335), .B1(new_n1348), .B2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1339), .B(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1296), .B1(new_n1324), .B2(KEYINPUT127), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1354), .B1(new_n1269), .B2(G375), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1353), .B(new_n1355), .ZN(G402));
endmodule


