

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XNOR2_X1 U326 ( .A(n472), .B(n471), .ZN(n576) );
  XNOR2_X1 U327 ( .A(n312), .B(n311), .ZN(n361) );
  XNOR2_X1 U328 ( .A(n467), .B(n466), .ZN(n554) );
  XNOR2_X1 U329 ( .A(n432), .B(n431), .ZN(n583) );
  XNOR2_X1 U330 ( .A(n430), .B(n294), .ZN(n431) );
  XNOR2_X1 U331 ( .A(n476), .B(n475), .ZN(n477) );
  AND2_X1 U332 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U333 ( .A(n367), .B(n366), .Z(n295) );
  NOR2_X1 U334 ( .A1(n543), .A2(n507), .ZN(n388) );
  INV_X1 U335 ( .A(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U336 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U337 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U338 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n466) );
  XNOR2_X1 U339 ( .A(n406), .B(n405), .ZN(n408) );
  INV_X1 U340 ( .A(KEYINPUT64), .ZN(n471) );
  XNOR2_X1 U341 ( .A(n414), .B(n413), .ZN(n415) );
  OR2_X1 U342 ( .A1(n528), .A2(n496), .ZN(n451) );
  XNOR2_X1 U343 ( .A(n416), .B(n415), .ZN(n586) );
  XNOR2_X1 U344 ( .A(n566), .B(KEYINPUT113), .ZN(n572) );
  XNOR2_X1 U345 ( .A(n451), .B(KEYINPUT38), .ZN(n513) );
  XNOR2_X1 U346 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U347 ( .A(n452), .B(G29GAT), .ZN(n453) );
  XNOR2_X1 U348 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n454), .B(n453), .ZN(G1328GAT) );
  XOR2_X1 U350 ( .A(G57GAT), .B(G148GAT), .Z(n297) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(G127GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U353 ( .A(G85GAT), .B(G162GAT), .Z(n299) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(G155GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n320) );
  XOR2_X1 U357 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n303) );
  XNOR2_X1 U358 ( .A(KEYINPUT91), .B(KEYINPUT5), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n305) );
  XNOR2_X1 U361 ( .A(KEYINPUT93), .B(KEYINPUT92), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U363 ( .A(n307), .B(n306), .Z(n318) );
  XNOR2_X1 U364 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n308) );
  XNOR2_X1 U365 ( .A(n308), .B(KEYINPUT83), .ZN(n312) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(G120GAT), .ZN(n310) );
  XOR2_X1 U367 ( .A(G134GAT), .B(KEYINPUT77), .Z(n330) );
  XNOR2_X1 U368 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n313) );
  XNOR2_X1 U369 ( .A(n313), .B(KEYINPUT2), .ZN(n343) );
  XOR2_X1 U370 ( .A(n330), .B(n343), .Z(n315) );
  NAND2_X1 U371 ( .A1(G225GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U372 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n361), .B(n316), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U375 ( .A(n320), .B(n319), .Z(n555) );
  INV_X1 U376 ( .A(n555), .ZN(n469) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(G190GAT), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n321), .B(G218GAT), .ZN(n383) );
  XOR2_X1 U379 ( .A(n383), .B(G106GAT), .Z(n323) );
  NAND2_X1 U380 ( .A1(G232GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n337) );
  XOR2_X1 U382 ( .A(KEYINPUT67), .B(KEYINPUT76), .Z(n325) );
  XNOR2_X1 U383 ( .A(KEYINPUT65), .B(KEYINPUT78), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U385 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n327) );
  XNOR2_X1 U386 ( .A(G92GAT), .B(KEYINPUT74), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U388 ( .A(n329), .B(n328), .Z(n335) );
  XOR2_X1 U389 ( .A(G50GAT), .B(G162GAT), .Z(n346) );
  XOR2_X1 U390 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n332) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n430) );
  XNOR2_X1 U392 ( .A(n330), .B(n430), .ZN(n331) );
  XNOR2_X1 U393 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n346), .B(n333), .ZN(n334) );
  XNOR2_X1 U395 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U396 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U397 ( .A(KEYINPUT69), .B(KEYINPUT8), .Z(n339) );
  XNOR2_X1 U398 ( .A(G43GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U400 ( .A(KEYINPUT7), .B(n340), .ZN(n449) );
  XOR2_X1 U401 ( .A(n341), .B(n449), .Z(n490) );
  XNOR2_X1 U402 ( .A(KEYINPUT36), .B(n490), .ZN(n589) );
  XNOR2_X1 U403 ( .A(G22GAT), .B(G155GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n342), .B(G78GAT), .ZN(n410) );
  XNOR2_X1 U405 ( .A(n343), .B(n410), .ZN(n357) );
  XOR2_X1 U406 ( .A(G197GAT), .B(KEYINPUT21), .Z(n375) );
  XOR2_X1 U407 ( .A(G106GAT), .B(G148GAT), .Z(n422) );
  XOR2_X1 U408 ( .A(n375), .B(n422), .Z(n345) );
  NAND2_X1 U409 ( .A1(G228GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n347) );
  XOR2_X1 U411 ( .A(n347), .B(n346), .Z(n355) );
  XOR2_X1 U412 ( .A(KEYINPUT22), .B(G204GAT), .Z(n349) );
  XNOR2_X1 U413 ( .A(G218GAT), .B(KEYINPUT90), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U415 ( .A(KEYINPUT89), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U416 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U420 ( .A(n357), .B(n356), .ZN(n474) );
  XOR2_X1 U421 ( .A(G15GAT), .B(G127GAT), .Z(n401) );
  XOR2_X1 U422 ( .A(n401), .B(KEYINPUT20), .Z(n359) );
  NAND2_X1 U423 ( .A1(G227GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U425 ( .A(n360), .B(G99GAT), .Z(n363) );
  XNOR2_X1 U426 ( .A(G43GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U428 ( .A(G176GAT), .B(G71GAT), .Z(n365) );
  XNOR2_X1 U429 ( .A(G190GAT), .B(G134GAT), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U431 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n369) );
  XNOR2_X1 U432 ( .A(KEYINPUT17), .B(KEYINPUT86), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U434 ( .A(G169GAT), .B(n370), .Z(n387) );
  XOR2_X1 U435 ( .A(G183GAT), .B(KEYINPUT87), .Z(n372) );
  XNOR2_X1 U436 ( .A(KEYINPUT66), .B(KEYINPUT88), .ZN(n371) );
  XNOR2_X1 U437 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U438 ( .A(n387), .B(n373), .ZN(n374) );
  XOR2_X1 U439 ( .A(n295), .B(n374), .Z(n535) );
  INV_X1 U440 ( .A(n535), .ZN(n543) );
  XOR2_X1 U441 ( .A(KEYINPUT95), .B(n375), .Z(n377) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U443 ( .A(n377), .B(n376), .ZN(n380) );
  XOR2_X1 U444 ( .A(G211GAT), .B(KEYINPUT79), .Z(n379) );
  XNOR2_X1 U445 ( .A(G8GAT), .B(G183GAT), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n379), .B(n378), .ZN(n402) );
  XOR2_X1 U447 ( .A(n380), .B(n402), .Z(n385) );
  XOR2_X1 U448 ( .A(G64GAT), .B(G92GAT), .Z(n382) );
  XNOR2_X1 U449 ( .A(G176GAT), .B(G204GAT), .ZN(n381) );
  XNOR2_X1 U450 ( .A(n382), .B(n381), .ZN(n427) );
  XNOR2_X1 U451 ( .A(n427), .B(n383), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U453 ( .A(n387), .B(n386), .Z(n531) );
  INV_X1 U454 ( .A(n531), .ZN(n507) );
  XNOR2_X1 U455 ( .A(n388), .B(KEYINPUT98), .ZN(n389) );
  NOR2_X1 U456 ( .A1(n474), .A2(n389), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n390), .B(KEYINPUT25), .ZN(n393) );
  XOR2_X1 U458 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n391) );
  XOR2_X1 U459 ( .A(n531), .B(n391), .Z(n396) );
  NAND2_X1 U460 ( .A1(n474), .A2(n543), .ZN(n392) );
  XOR2_X1 U461 ( .A(KEYINPUT26), .B(n392), .Z(n575) );
  NAND2_X1 U462 ( .A1(n396), .A2(n575), .ZN(n556) );
  NAND2_X1 U463 ( .A1(n393), .A2(n556), .ZN(n394) );
  NAND2_X1 U464 ( .A1(n394), .A2(n469), .ZN(n395) );
  XNOR2_X1 U465 ( .A(KEYINPUT99), .B(n395), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n474), .B(KEYINPUT28), .ZN(n538) );
  INV_X1 U467 ( .A(n538), .ZN(n514) );
  NAND2_X1 U468 ( .A1(n396), .A2(n514), .ZN(n397) );
  NOR2_X1 U469 ( .A1(n469), .A2(n397), .ZN(n541) );
  NAND2_X1 U470 ( .A1(n543), .A2(n541), .ZN(n398) );
  XNOR2_X1 U471 ( .A(KEYINPUT97), .B(n398), .ZN(n399) );
  NOR2_X1 U472 ( .A1(n400), .A2(n399), .ZN(n493) );
  XNOR2_X1 U473 ( .A(n402), .B(n401), .ZN(n406) );
  AND2_X1 U474 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  INV_X1 U475 ( .A(KEYINPUT81), .ZN(n403) );
  XOR2_X1 U476 ( .A(KEYINPUT70), .B(G1GAT), .Z(n444) );
  XNOR2_X1 U477 ( .A(n444), .B(G64GAT), .ZN(n407) );
  XNOR2_X1 U478 ( .A(n408), .B(n407), .ZN(n416) );
  XNOR2_X1 U479 ( .A(G71GAT), .B(G57GAT), .ZN(n409) );
  XNOR2_X1 U480 ( .A(n409), .B(KEYINPUT13), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n410), .B(n426), .ZN(n414) );
  XOR2_X1 U482 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n412) );
  XNOR2_X1 U483 ( .A(KEYINPUT14), .B(KEYINPUT15), .ZN(n411) );
  XNOR2_X1 U484 ( .A(n412), .B(n411), .ZN(n413) );
  INV_X1 U485 ( .A(n586), .ZN(n566) );
  NOR2_X1 U486 ( .A1(n493), .A2(n566), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n417), .B(KEYINPUT103), .ZN(n418) );
  NOR2_X1 U488 ( .A1(n589), .A2(n418), .ZN(n419) );
  XNOR2_X1 U489 ( .A(KEYINPUT37), .B(n419), .ZN(n528) );
  XOR2_X1 U490 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n421) );
  XNOR2_X1 U491 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n420) );
  XNOR2_X1 U492 ( .A(n421), .B(n420), .ZN(n425) );
  XNOR2_X1 U493 ( .A(G120GAT), .B(G78GAT), .ZN(n423) );
  XNOR2_X1 U494 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U495 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U497 ( .A(n429), .B(n428), .ZN(n432) );
  XOR2_X1 U498 ( .A(KEYINPUT30), .B(KEYINPUT72), .Z(n434) );
  XNOR2_X1 U499 ( .A(KEYINPUT68), .B(KEYINPUT71), .ZN(n433) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n448) );
  XOR2_X1 U501 ( .A(G22GAT), .B(G141GAT), .Z(n436) );
  XNOR2_X1 U502 ( .A(G50GAT), .B(G36GAT), .ZN(n435) );
  XNOR2_X1 U503 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U504 ( .A(G15GAT), .B(G113GAT), .Z(n438) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(G197GAT), .ZN(n437) );
  XNOR2_X1 U506 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U507 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U508 ( .A(KEYINPUT29), .B(G8GAT), .Z(n442) );
  NAND2_X1 U509 ( .A1(G229GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U510 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U513 ( .A(n448), .B(n447), .ZN(n450) );
  XOR2_X1 U514 ( .A(n450), .B(n449), .Z(n577) );
  INV_X1 U515 ( .A(n577), .ZN(n559) );
  NAND2_X1 U516 ( .A1(n583), .A2(n559), .ZN(n496) );
  NOR2_X1 U517 ( .A1(n469), .A2(n513), .ZN(n454) );
  XNOR2_X1 U518 ( .A(KEYINPUT39), .B(KEYINPUT104), .ZN(n452) );
  INV_X1 U519 ( .A(n490), .ZN(n568) );
  XNOR2_X1 U520 ( .A(n583), .B(KEYINPUT41), .ZN(n561) );
  NAND2_X1 U521 ( .A1(n561), .A2(n559), .ZN(n455) );
  XNOR2_X1 U522 ( .A(n455), .B(KEYINPUT46), .ZN(n456) );
  XNOR2_X1 U523 ( .A(n456), .B(KEYINPUT114), .ZN(n457) );
  NAND2_X1 U524 ( .A1(n457), .A2(n572), .ZN(n458) );
  NOR2_X1 U525 ( .A1(n568), .A2(n458), .ZN(n459) );
  XNOR2_X1 U526 ( .A(n459), .B(KEYINPUT47), .ZN(n465) );
  NOR2_X1 U527 ( .A1(n589), .A2(n586), .ZN(n460) );
  XNOR2_X1 U528 ( .A(KEYINPUT45), .B(n460), .ZN(n461) );
  NAND2_X1 U529 ( .A1(n461), .A2(n583), .ZN(n462) );
  XNOR2_X1 U530 ( .A(KEYINPUT115), .B(n462), .ZN(n463) );
  NAND2_X1 U531 ( .A1(n463), .A2(n577), .ZN(n464) );
  NAND2_X1 U532 ( .A1(n465), .A2(n464), .ZN(n467) );
  AND2_X1 U533 ( .A1(n554), .A2(n531), .ZN(n468) );
  XNOR2_X1 U534 ( .A(KEYINPUT54), .B(n468), .ZN(n470) );
  NAND2_X1 U535 ( .A1(n470), .A2(n469), .ZN(n472) );
  INV_X1 U536 ( .A(n576), .ZN(n473) );
  NOR2_X1 U537 ( .A1(n474), .A2(n473), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n476) );
  INV_X1 U539 ( .A(KEYINPUT55), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U541 ( .A1(n543), .A2(n479), .ZN(n571) );
  NAND2_X1 U542 ( .A1(n571), .A2(n561), .ZN(n483) );
  XOR2_X1 U543 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n481) );
  XOR2_X1 U544 ( .A(G176GAT), .B(KEYINPUT56), .Z(n480) );
  XNOR2_X1 U545 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  NAND2_X1 U547 ( .A1(n571), .A2(n568), .ZN(n487) );
  XOR2_X1 U548 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n485) );
  XNOR2_X1 U549 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n484) );
  NAND2_X1 U550 ( .A1(n559), .A2(n571), .ZN(n489) );
  XNOR2_X1 U551 ( .A(KEYINPUT122), .B(G169GAT), .ZN(n488) );
  XNOR2_X1 U552 ( .A(n489), .B(n488), .ZN(G1348GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT100), .B(KEYINPUT34), .Z(n498) );
  XOR2_X1 U554 ( .A(KEYINPUT82), .B(KEYINPUT16), .Z(n492) );
  NAND2_X1 U555 ( .A1(n566), .A2(n490), .ZN(n491) );
  XNOR2_X1 U556 ( .A(n492), .B(n491), .ZN(n495) );
  INV_X1 U557 ( .A(n493), .ZN(n494) );
  NAND2_X1 U558 ( .A1(n495), .A2(n494), .ZN(n516) );
  NOR2_X1 U559 ( .A1(n496), .A2(n516), .ZN(n504) );
  NAND2_X1 U560 ( .A1(n504), .A2(n555), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U562 ( .A(G1GAT), .B(n499), .Z(G1324GAT) );
  NAND2_X1 U563 ( .A1(n504), .A2(n531), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n500), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT35), .B(KEYINPUT101), .Z(n502) );
  NAND2_X1 U566 ( .A1(n504), .A2(n535), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U568 ( .A(G15GAT), .B(n503), .Z(G1326GAT) );
  NAND2_X1 U569 ( .A1(n538), .A2(n504), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n505), .B(KEYINPUT102), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G22GAT), .B(n506), .ZN(G1327GAT) );
  NOR2_X1 U572 ( .A1(n513), .A2(n507), .ZN(n508) );
  XOR2_X1 U573 ( .A(G36GAT), .B(n508), .Z(G1329GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n510) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n512) );
  NOR2_X1 U577 ( .A1(n543), .A2(n513), .ZN(n511) );
  XOR2_X1 U578 ( .A(n512), .B(n511), .Z(G1330GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XOR2_X1 U580 ( .A(G50GAT), .B(n515), .Z(G1331GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT107), .B(KEYINPUT42), .Z(n518) );
  NAND2_X1 U582 ( .A1(n577), .A2(n561), .ZN(n527) );
  NOR2_X1 U583 ( .A1(n527), .A2(n516), .ZN(n522) );
  NAND2_X1 U584 ( .A1(n522), .A2(n555), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(n519), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n531), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U589 ( .A1(n535), .A2(n522), .ZN(n521) );
  XNOR2_X1 U590 ( .A(n521), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U592 ( .A1(n522), .A2(n538), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(n526) );
  XOR2_X1 U594 ( .A(G78GAT), .B(KEYINPUT109), .Z(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1335GAT) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(KEYINPUT110), .ZN(n530) );
  NOR2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n537), .A2(n555), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(G1336GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n533) );
  NAND2_X1 U601 ( .A1(n537), .A2(n531), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U603 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NAND2_X1 U604 ( .A1(n535), .A2(n537), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n536), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U606 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n539), .B(KEYINPUT44), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n540), .ZN(G1339GAT) );
  NAND2_X1 U609 ( .A1(n541), .A2(n554), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n543), .A2(n542), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n559), .A2(n551), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n544), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U614 ( .A1(n551), .A2(n561), .ZN(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U616 ( .A(G120GAT), .B(n547), .Z(G1341GAT) );
  INV_X1 U617 ( .A(n551), .ZN(n548) );
  NOR2_X1 U618 ( .A1(n572), .A2(n548), .ZN(n549) );
  XOR2_X1 U619 ( .A(KEYINPUT50), .B(n549), .Z(n550) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n553) );
  NAND2_X1 U622 ( .A1(n551), .A2(n568), .ZN(n552) );
  XNOR2_X1 U623 ( .A(n553), .B(n552), .ZN(G1343GAT) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n557) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT118), .ZN(n569) );
  NAND2_X1 U627 ( .A1(n569), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n560), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U630 ( .A1(n569), .A2(n561), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n565) );
  XOR2_X1 U632 ( .A(G148GAT), .B(KEYINPUT53), .Z(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(G1345GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G162GAT), .ZN(G1347GAT) );
  INV_X1 U638 ( .A(n571), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U640 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n588) );
  NOR2_X1 U642 ( .A1(n577), .A2(n588), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT126), .B(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n588), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

