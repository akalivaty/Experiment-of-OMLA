//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1315, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1324, new_n1325, new_n1326, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT0), .ZN(new_n207));
  AND2_X1   g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G20), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT65), .Z(new_n211));
  OAI22_X1  g0011(.A1(new_n206), .A2(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(new_n207), .B2(new_n206), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT67), .B(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n221), .A2(G77), .B1(G68), .B2(G238), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT66), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n219), .B2(KEYINPUT68), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n204), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n213), .B1(KEYINPUT1), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n234), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT70), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT71), .ZN(new_n242));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n244), .B(new_n248), .ZN(G351));
  OR2_X1    g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  AOI21_X1  g0051(.A(G1698), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n251), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G223), .A3(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n253), .B(new_n255), .C1(new_n256), .C2(new_n254), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT73), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n208), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  INV_X1    g0066(.A(G41), .ZN(new_n267));
  INV_X1    g0067(.A(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(new_n269), .B1(new_n208), .B2(new_n262), .ZN(new_n270));
  OR2_X1    g0070(.A1(KEYINPUT72), .A2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT72), .A2(G45), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n267), .A3(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n266), .A2(G274), .ZN(new_n274));
  AOI22_X1  g0074(.A1(new_n270), .A2(G226), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n265), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G200), .ZN(new_n277));
  INV_X1    g0077(.A(G190), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n277), .B1(new_n278), .B2(new_n276), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n259), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n266), .A2(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(G50), .A3(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n283), .ZN(new_n290));
  XOR2_X1   g0090(.A(KEYINPUT8), .B(G58), .Z(new_n291));
  INV_X1    g0091(.A(KEYINPUT74), .ZN(new_n292));
  INV_X1    g0092(.A(G33), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n292), .B1(new_n293), .B2(G20), .ZN(new_n294));
  INV_X1    g0094(.A(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(KEYINPUT74), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G58), .ZN(new_n299));
  INV_X1    g0099(.A(G68), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n287), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n301), .A2(G20), .B1(G150), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n290), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n289), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n306));
  NAND2_X1  g0106(.A1(KEYINPUT78), .A2(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n289), .B2(new_n304), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(KEYINPUT78), .A2(KEYINPUT10), .ZN(new_n311));
  OR3_X1    g0111(.A1(new_n279), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n311), .B1(new_n279), .B2(new_n310), .ZN(new_n313));
  INV_X1    g0113(.A(G169), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n305), .B1(new_n276), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G179), .B2(new_n276), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT76), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n280), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n266), .A2(KEYINPUT76), .A3(G13), .A4(G20), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n283), .B1(new_n319), .B2(new_n320), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n256), .B1(new_n266), .B2(G20), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n322), .A2(new_n256), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT8), .B(G58), .ZN(new_n326));
  INV_X1    g0126(.A(new_n302), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n326), .A2(new_n327), .B1(new_n295), .B2(new_n256), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT15), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G87), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT75), .ZN(new_n332));
  AOI21_X1  g0132(.A(KEYINPUT75), .B1(new_n329), .B2(new_n331), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n328), .B1(new_n334), .B2(new_n297), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n325), .B1(new_n335), .B2(new_n290), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n270), .A2(new_n221), .B1(new_n273), .B2(new_n274), .ZN(new_n338));
  INV_X1    g0138(.A(G1698), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G238), .ZN(new_n340));
  NOR2_X1   g0140(.A1(G232), .A2(G1698), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n340), .A2(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G107), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n250), .A2(new_n345), .A3(new_n251), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n344), .A2(new_n260), .A3(new_n263), .A4(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n349), .A2(G169), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n348), .A2(G179), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n337), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G200), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n338), .B2(new_n347), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT77), .B1(new_n336), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n348), .A2(G200), .ZN(new_n356));
  INV_X1    g0156(.A(new_n328), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n329), .A2(new_n331), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT75), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n329), .A2(new_n331), .A3(KEYINPUT75), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n297), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n283), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT77), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n356), .A2(new_n364), .A3(new_n365), .A4(new_n325), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n349), .A2(G190), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n355), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n317), .A2(new_n352), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n297), .A2(G77), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n302), .A2(G50), .B1(G20), .B2(new_n300), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n283), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT11), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n323), .A2(G68), .A3(new_n285), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT12), .B1(new_n321), .B2(G68), .ZN(new_n379));
  INV_X1    g0179(.A(G13), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(G1), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n381), .A2(new_n382), .A3(G20), .A4(new_n300), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n379), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n260), .A2(new_n263), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  INV_X1    g0187(.A(G226), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(new_n339), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n231), .A2(G1698), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n389), .B(new_n390), .C1(new_n342), .C2(new_n343), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n386), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n273), .A2(new_n274), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n269), .A2(new_n266), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n208), .A2(new_n262), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G238), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n393), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n392), .B2(new_n398), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n399), .A2(G190), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n391), .A2(new_n387), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n264), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n270), .A2(G238), .B1(new_n273), .B2(new_n274), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n385), .B1(new_n400), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n399), .A2(KEYINPUT79), .A3(new_n405), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT79), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n402), .A2(new_n408), .A3(new_n403), .A4(new_n404), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n407), .A2(G200), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n407), .A2(G169), .A3(new_n409), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT14), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT14), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n407), .A2(new_n414), .A3(G169), .A4(new_n409), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n399), .A2(G179), .A3(new_n405), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n385), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n370), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n250), .A2(new_n295), .A3(new_n251), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT7), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n295), .A4(new_n251), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n300), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n299), .A2(new_n300), .ZN(new_n426));
  NOR2_X1   g0226(.A1(G58), .A2(G68), .ZN(new_n427));
  OAI21_X1  g0227(.A(G20), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n302), .A2(G159), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n420), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n342), .A2(new_n343), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT7), .B1(new_n432), .B2(new_n295), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n342), .A2(new_n343), .A3(new_n422), .A4(G20), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n430), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n435), .A2(KEYINPUT16), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n431), .A2(new_n437), .A3(new_n283), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n326), .A2(new_n281), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n291), .A2(new_n285), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n290), .A2(new_n280), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT80), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT80), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n439), .C1(new_n440), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n438), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G87), .ZN(new_n448));
  OR2_X1    g0248(.A1(G223), .A2(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n388), .A2(G1698), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n254), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n386), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n393), .B1(new_n396), .B2(new_n231), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n452), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n449), .A2(new_n450), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n448), .B1(new_n456), .B2(new_n432), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n264), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n270), .A2(G232), .B1(new_n273), .B2(new_n274), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT81), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n314), .B1(new_n455), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n459), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G179), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n447), .A2(KEYINPUT18), .A3(new_n461), .A4(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n454), .B1(new_n452), .B2(new_n453), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n459), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n463), .B1(new_n470), .B2(new_n314), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n471), .A2(KEYINPUT82), .A3(new_n447), .A4(KEYINPUT18), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT18), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n461), .A2(new_n464), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n435), .A2(new_n436), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n290), .B1(new_n475), .B2(new_n420), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n476), .A2(new_n437), .B1(new_n443), .B2(new_n445), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n467), .A2(new_n472), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(G200), .B1(new_n468), .B2(new_n469), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n462), .A2(G190), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n438), .B(new_n446), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT17), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n353), .B1(new_n455), .B2(new_n460), .ZN(new_n485));
  INV_X1    g0285(.A(new_n481), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(KEYINPUT17), .B1(new_n487), .B2(new_n477), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n479), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n419), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n268), .A2(G1), .ZN(new_n493));
  AND2_X1   g0293(.A1(KEYINPUT5), .A2(G41), .ZN(new_n494));
  NOR2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n496), .A2(G270), .A3(new_n395), .ZN(new_n497));
  XNOR2_X1  g0297(.A(KEYINPUT5), .B(G41), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n498), .A2(new_n395), .A3(G274), .A4(new_n493), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n502));
  OAI211_X1 g0302(.A(G257), .B(new_n339), .C1(new_n342), .C2(new_n343), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n250), .A2(G303), .A3(new_n251), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT84), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n505), .A2(new_n264), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n505), .B2(new_n264), .ZN(new_n508));
  OAI211_X1 g0308(.A(G190), .B(new_n501), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n510), .B1(new_n266), .B2(G33), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n322), .A2(new_n510), .B1(new_n323), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n282), .A2(new_n259), .B1(G20), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(new_n295), .C1(G33), .C2(new_n217), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT20), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n513), .A2(KEYINPUT20), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n264), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT84), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n505), .A2(new_n264), .A3(new_n506), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n500), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n509), .B(new_n522), .C1(new_n526), .C2(new_n353), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n525), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n497), .A2(new_n499), .A3(G179), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n521), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n501), .B1(new_n507), .B2(new_n508), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n314), .B1(new_n512), .B2(new_n520), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT21), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n531), .B2(new_n532), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n527), .B(new_n530), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n531), .A2(new_n532), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT21), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(KEYINPUT85), .A3(new_n530), .A4(new_n527), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n538), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n280), .A2(G97), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n266), .A2(G33), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n284), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n549), .B2(new_n217), .ZN(new_n550));
  OAI21_X1  g0350(.A(G107), .B1(new_n433), .B2(new_n434), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n327), .A2(new_n256), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT6), .ZN(new_n553));
  AND2_X1   g0353(.A1(G97), .A2(G107), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G97), .A2(G107), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n345), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n552), .B1(new_n558), .B2(G20), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n550), .B1(new_n560), .B2(new_n283), .ZN(new_n561));
  OAI211_X1 g0361(.A(G250), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n562));
  OAI211_X1 g0362(.A(G244), .B(new_n339), .C1(new_n342), .C2(new_n343), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n514), .B(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(KEYINPUT4), .B1(new_n252), .B2(G244), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n264), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n258), .A2(new_n259), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n568), .B1(new_n493), .B2(new_n498), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n395), .A2(G274), .A3(new_n493), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(G257), .B1(new_n570), .B2(new_n498), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n567), .A2(new_n278), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(G200), .B1(new_n567), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n561), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n567), .A2(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n314), .ZN(new_n576));
  INV_X1    g0376(.A(new_n552), .ZN(new_n577));
  INV_X1    g0377(.A(new_n557), .ZN(new_n578));
  XNOR2_X1  g0378(.A(G97), .B(G107), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n578), .B1(new_n553), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n577), .B1(new_n580), .B2(new_n295), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n345), .B1(new_n423), .B2(new_n424), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n283), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n550), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G179), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n567), .A2(new_n571), .A3(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n576), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n395), .A2(G274), .A3(new_n493), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n293), .A2(new_n510), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G238), .A2(G1698), .ZN(new_n591));
  INV_X1    g0391(.A(G244), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(G1698), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n590), .B1(new_n593), .B2(new_n254), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n589), .B1(new_n594), .B2(new_n386), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  OAI21_X1  g0396(.A(G250), .B1(new_n268), .B2(G1), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n596), .B1(new_n568), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n216), .B1(new_n266), .B2(G45), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n395), .A2(new_n599), .A3(KEYINPUT83), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n314), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n592), .A2(G1698), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G238), .B2(G1698), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n604), .A2(new_n432), .B1(new_n293), .B2(new_n510), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n570), .B1(new_n605), .B2(new_n264), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n598), .A2(new_n600), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n586), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT19), .B1(new_n297), .B2(G97), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n295), .B1(new_n387), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n555), .A2(new_n215), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n295), .B(G68), .C1(new_n342), .C2(new_n343), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n283), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n334), .A2(new_n284), .A3(new_n548), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n360), .A2(new_n361), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n322), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n602), .A2(new_n608), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(G200), .B1(new_n595), .B2(new_n601), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n217), .B1(new_n294), .B2(new_n296), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n614), .B(new_n613), .C1(new_n623), .C2(KEYINPUT19), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n624), .A2(new_n283), .B1(new_n618), .B2(new_n322), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n284), .A2(G87), .A3(new_n548), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n605), .A2(new_n264), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n627), .A2(G190), .A3(new_n607), .A4(new_n589), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n622), .A2(new_n625), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n574), .A2(new_n588), .A3(new_n621), .A4(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT23), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n295), .B2(G107), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n345), .A2(KEYINPUT23), .A3(G20), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n590), .A2(new_n295), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT22), .ZN(new_n637));
  AOI21_X1  g0437(.A(G20), .B1(new_n250), .B2(new_n251), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(G87), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n295), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n640), .A2(KEYINPUT22), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n636), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT86), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT24), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n634), .A2(new_n635), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(KEYINPUT22), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n254), .A2(new_n637), .A3(new_n295), .A4(G87), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT24), .B1(new_n649), .B2(KEYINPUT86), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n643), .B(new_n646), .C1(new_n647), .C2(new_n648), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n645), .B(new_n283), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n281), .A2(new_n345), .ZN(new_n653));
  XNOR2_X1  g0453(.A(new_n653), .B(KEYINPUT25), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n549), .A2(new_n345), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n496), .A2(G264), .A3(new_n395), .ZN(new_n657));
  NOR2_X1   g0457(.A1(G250), .A2(G1698), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n218), .B2(G1698), .ZN(new_n659));
  XNOR2_X1  g0459(.A(KEYINPUT87), .B(G294), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n659), .A2(new_n254), .B1(new_n660), .B2(G33), .ZN(new_n661));
  OAI211_X1 g0461(.A(new_n499), .B(new_n657), .C1(new_n661), .C2(new_n386), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n353), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(G190), .B2(new_n662), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n652), .A2(new_n656), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n656), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n649), .A2(KEYINPUT86), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n290), .B1(new_n667), .B2(new_n644), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n642), .A2(new_n643), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n649), .A2(KEYINPUT86), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(KEYINPUT24), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n666), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n662), .A2(new_n673), .A3(G169), .ZN(new_n674));
  XOR2_X1   g0474(.A(KEYINPUT87), .B(G294), .Z(new_n675));
  NAND2_X1  g0475(.A1(new_n218), .A2(G1698), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n676), .B1(G250), .B2(G1698), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n675), .A2(new_n293), .B1(new_n677), .B2(new_n432), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n264), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(G179), .A3(new_n499), .A4(new_n657), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n674), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n673), .B1(new_n662), .B2(G169), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n665), .B1(new_n672), .B2(new_n683), .ZN(new_n684));
  NOR4_X1   g0484(.A1(new_n492), .A2(new_n545), .A3(new_n630), .A4(new_n684), .ZN(G372));
  NAND2_X1  g0485(.A1(new_n482), .A2(new_n483), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n487), .A2(new_n477), .A3(KEYINPUT17), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n411), .A2(new_n352), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n688), .B1(new_n418), .B2(new_n689), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n471), .A2(KEYINPUT18), .A3(new_n447), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT18), .B1(new_n471), .B2(new_n447), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n313), .B(new_n312), .C1(new_n690), .C2(new_n693), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n694), .A2(new_n316), .ZN(new_n695));
  INV_X1    g0495(.A(new_n587), .ZN(new_n696));
  AOI21_X1  g0496(.A(G169), .B1(new_n567), .B2(new_n571), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n696), .A2(new_n561), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(KEYINPUT26), .A3(new_n621), .A4(new_n629), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT26), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n629), .A2(new_n621), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n588), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n704));
  INV_X1    g0504(.A(new_n682), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n674), .A2(new_n680), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(new_n652), .B2(new_n656), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n629), .A2(new_n621), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n709), .A2(new_n665), .A3(new_n588), .A4(new_n574), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n703), .B(new_n621), .C1(new_n708), .C2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n695), .B1(new_n492), .B2(new_n712), .ZN(G369));
  INV_X1    g0513(.A(new_n684), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n381), .A2(new_n295), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT27), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(KEYINPUT27), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G213), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G343), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n672), .A2(KEYINPUT90), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT90), .B1(new_n672), .B2(new_n721), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n714), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n707), .A2(new_n720), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n704), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n521), .A2(new_n720), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n544), .B2(new_n729), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(KEYINPUT89), .A3(G330), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT89), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n734), .B1(new_n731), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n727), .B1(new_n733), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n720), .B1(new_n542), .B2(new_n530), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n714), .A2(new_n738), .A3(new_n722), .A4(new_n723), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n707), .A2(new_n721), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n737), .A2(new_n741), .ZN(G399));
  INV_X1    g0542(.A(new_n205), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G41), .ZN(new_n744));
  NOR4_X1   g0544(.A1(new_n744), .A2(new_n266), .A3(G116), .A4(new_n612), .ZN(new_n745));
  INV_X1    g0545(.A(new_n210), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n744), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  NAND2_X1  g0548(.A1(new_n711), .A2(new_n721), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n699), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n702), .A2(KEYINPUT93), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT93), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n754), .B(new_n700), .C1(new_n701), .C2(new_n588), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n621), .B1(new_n708), .B2(new_n710), .ZN(new_n757));
  OAI211_X1 g0557(.A(KEYINPUT29), .B(new_n721), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n567), .A2(KEYINPUT30), .A3(new_n571), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n595), .A2(new_n601), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n657), .B1(new_n661), .B2(new_n386), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n762), .A2(new_n586), .A3(new_n500), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n760), .A2(new_n528), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(G179), .B1(new_n606), .B2(new_n607), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n531), .A2(new_n575), .A3(new_n765), .A4(new_n662), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n678), .A2(new_n264), .B1(new_n569), .B2(G264), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n768), .A2(new_n529), .A3(new_n606), .A4(new_n607), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n507), .A2(new_n508), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n575), .ZN(new_n772));
  AOI21_X1  g0572(.A(KEYINPUT30), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(KEYINPUT91), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n772), .A2(new_n528), .A3(new_n761), .A4(new_n763), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT30), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT91), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n777), .A2(new_n778), .A3(new_n766), .A4(new_n764), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n774), .A2(new_n779), .A3(new_n720), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT31), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n684), .A2(new_n630), .A3(new_n720), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n544), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g0584(.A(KEYINPUT31), .B(new_n720), .C1(new_n767), .C2(new_n773), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G330), .ZN(new_n787));
  AND2_X1   g0587(.A1(new_n759), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n748), .B1(new_n788), .B2(G1), .ZN(G364));
  NOR2_X1   g0589(.A1(new_n380), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n266), .B1(new_n790), .B2(G45), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n744), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n259), .B1(G20), .B2(new_n314), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n295), .A2(new_n586), .A3(new_n353), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n278), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G326), .ZN(new_n801));
  INV_X1    g0601(.A(G283), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n295), .A2(G179), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n803), .A2(new_n278), .A3(G200), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n803), .A2(G190), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(G303), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n295), .A2(G190), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n586), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  INV_X1    g0612(.A(G322), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n810), .A2(G20), .A3(G190), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n432), .B1(new_n811), .B2(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n809), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n586), .A2(new_n353), .A3(KEYINPUT96), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT96), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(G179), .B2(G200), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n815), .B1(G329), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g0621(.A1(new_n808), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n278), .B1(new_n817), .B2(new_n819), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n295), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n798), .A2(KEYINPUT97), .A3(G190), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT97), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n797), .B2(new_n278), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g0628(.A(KEYINPUT33), .B(G317), .Z(new_n829));
  OAI221_X1 g0629(.A(new_n822), .B1(new_n675), .B2(new_n824), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n814), .ZN(new_n831));
  INV_X1    g0631(.A(new_n811), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n831), .A2(G58), .B1(new_n832), .B2(G77), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n800), .B2(new_n287), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT95), .Z(new_n835));
  NAND2_X1  g0635(.A1(new_n820), .A2(G159), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT32), .ZN(new_n837));
  INV_X1    g0637(.A(new_n824), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G97), .A2(new_n838), .B1(new_n836), .B2(KEYINPUT32), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n804), .A2(new_n345), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n254), .B1(new_n806), .B2(new_n215), .ZN(new_n841));
  INV_X1    g0641(.A(new_n828), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n840), .B(new_n841), .C1(new_n842), .C2(G68), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n835), .A2(new_n837), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n796), .B1(new_n830), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(G13), .A2(G33), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n847), .A2(G20), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n795), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n743), .A2(new_n254), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n271), .A2(new_n272), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n211), .B2(new_n851), .C1(new_n244), .C2(new_n268), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n205), .A2(G355), .A3(new_n254), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n853), .C1(G116), .C2(new_n205), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n794), .B(new_n845), .C1(new_n849), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n848), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n855), .B1(new_n732), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n731), .A2(new_n735), .ZN(new_n858));
  XOR2_X1   g0658(.A(new_n858), .B(KEYINPUT94), .Z(new_n859));
  NAND3_X1  g0659(.A1(new_n733), .A2(new_n736), .A3(new_n794), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n857), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT98), .ZN(G396));
  NAND2_X1  g0662(.A1(new_n336), .A2(new_n720), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n352), .B1(new_n368), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n352), .A2(new_n721), .ZN(new_n865));
  OAI21_X1  g0665(.A(KEYINPUT100), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT100), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n352), .A2(new_n721), .ZN(new_n868));
  INV_X1    g0668(.A(new_n863), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n356), .A2(new_n364), .A3(new_n325), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n870), .A2(KEYINPUT77), .B1(G190), .B2(new_n349), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n871), .B2(new_n366), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n867), .B(new_n868), .C1(new_n872), .C2(new_n352), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n749), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n874), .A2(new_n711), .A3(new_n721), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n793), .B1(new_n878), .B2(new_n787), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n787), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n795), .A2(new_n846), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT99), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n793), .B1(G77), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(G294), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n432), .B1(new_n811), .B2(new_n510), .C1(new_n884), .C2(new_n814), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n804), .A2(new_n215), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n886), .B1(new_n799), .B2(G303), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n345), .B2(new_n806), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n885), .B(new_n888), .C1(G311), .C2(new_n820), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n889), .B1(new_n217), .B2(new_n824), .C1(new_n802), .C2(new_n828), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n831), .A2(G143), .B1(new_n832), .B2(G159), .ZN(new_n891));
  INV_X1    g0691(.A(G137), .ZN(new_n892));
  INV_X1    g0692(.A(G150), .ZN(new_n893));
  OAI221_X1 g0693(.A(new_n891), .B1(new_n892), .B2(new_n800), .C1(new_n828), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT34), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n254), .B1(new_n806), .B2(new_n287), .C1(new_n300), .C2(new_n804), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(G132), .B2(new_n820), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n896), .B(new_n898), .C1(new_n299), .C2(new_n824), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n894), .A2(new_n895), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n890), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n883), .B1(new_n901), .B2(new_n795), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n874), .B2(new_n847), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n880), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(G384));
  NOR2_X1   g0705(.A1(new_n209), .A2(new_n510), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n558), .B(KEYINPUT101), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT35), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n909), .B2(new_n908), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT36), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n746), .B(G77), .C1(new_n299), .C2(new_n300), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n287), .A2(G68), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n266), .B(G13), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n790), .A2(new_n266), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT39), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n471), .A2(new_n447), .ZN(new_n919));
  INV_X1    g0719(.A(new_n718), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n447), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT37), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n919), .A2(new_n482), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT103), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT16), .B1(new_n435), .B2(new_n436), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n290), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n431), .A2(KEYINPUT103), .A3(new_n283), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n437), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n442), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n920), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n471), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n933), .A3(new_n482), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n924), .B1(new_n934), .B2(KEYINPUT37), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n932), .B1(new_n479), .B2(new_n489), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT38), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n921), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n693), .B2(new_n688), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n919), .A2(new_n482), .A3(new_n921), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT37), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n923), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n918), .B1(new_n938), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n418), .A2(new_n720), .ZN(new_n946));
  INV_X1    g0746(.A(new_n437), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n431), .A2(new_n283), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n948), .B2(new_n925), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n442), .B1(new_n949), .B2(new_n928), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n950), .A2(new_n718), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n490), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n482), .B1(new_n950), .B2(new_n474), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT37), .B1(new_n953), .B2(new_n951), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n923), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n955), .A3(KEYINPUT38), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n937), .B1(new_n935), .B2(new_n936), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT39), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n945), .A2(new_n946), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n693), .A2(new_n718), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n956), .A2(new_n957), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n385), .A2(new_n720), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n418), .A2(new_n411), .A3(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n411), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n385), .B(new_n720), .C1(new_n964), .C2(new_n417), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(new_n868), .B2(new_n877), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT102), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n961), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n877), .A2(new_n868), .ZN(new_n970));
  INV_X1    g0770(.A(new_n966), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(KEYINPUT102), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n959), .B(new_n960), .C1(new_n969), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n491), .A2(new_n758), .A3(new_n751), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n695), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n974), .B(new_n976), .Z(new_n977));
  NAND4_X1  g0777(.A1(new_n774), .A2(new_n779), .A3(KEYINPUT31), .A4(new_n720), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n782), .A2(new_n784), .A3(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n963), .A2(new_n965), .B1(new_n873), .B2(new_n866), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n961), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT40), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n940), .A2(new_n943), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n937), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n956), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g0786(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT40), .ZN(new_n987));
  AOI22_X1  g0787(.A1(new_n982), .A2(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n988), .A2(new_n491), .A3(new_n979), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n988), .B1(new_n491), .B2(new_n979), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n989), .A2(new_n990), .A3(new_n735), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n917), .B1(new_n977), .B2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT104), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n992), .A2(new_n993), .B1(new_n977), .B2(new_n991), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n916), .B1(new_n994), .B2(new_n995), .ZN(G367));
  INV_X1    g0796(.A(new_n850), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n238), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n849), .B1(new_n205), .B2(new_n618), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n793), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n800), .A2(new_n1001), .B1(new_n256), .B2(new_n804), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(G58), .B2(new_n807), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n254), .B1(new_n811), .B2(new_n287), .C1(new_n893), .C2(new_n814), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G137), .B2(new_n820), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n842), .A2(G159), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n838), .A2(G68), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n807), .A2(G116), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT46), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n345), .B2(new_n824), .C1(new_n675), .C2(new_n828), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n804), .A2(new_n217), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n799), .B2(G311), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n820), .A2(G317), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n832), .A2(G283), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n254), .B1(new_n831), .B2(G303), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1008), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1000), .B1(new_n1019), .B2(new_n795), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n625), .A2(new_n626), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n720), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n709), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n1022), .A2(new_n621), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n848), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1020), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT45), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n574), .B(new_n588), .C1(new_n561), .C2(new_n721), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n698), .A2(new_n720), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1027), .B1(new_n741), .B2(new_n1031), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n739), .A2(KEYINPUT45), .A3(new_n740), .A4(new_n1030), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1030), .B1(new_n739), .B2(new_n740), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(new_n737), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n733), .A2(new_n736), .A3(KEYINPUT108), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n739), .B1(new_n726), .B2(new_n738), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n733), .A2(new_n736), .A3(KEYINPUT108), .A4(new_n1042), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n788), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n744), .B(KEYINPUT41), .Z(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n792), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1023), .A2(new_n1051), .A3(new_n1024), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT106), .Z(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n739), .A2(new_n1031), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n652), .A2(new_n656), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n705), .A2(new_n680), .A3(new_n674), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n588), .B1(new_n1028), .B2(new_n1058), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n1055), .A2(KEYINPUT42), .B1(new_n721), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(KEYINPUT42), .B2(new_n1055), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(KEYINPUT43), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1054), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1061), .A2(new_n1054), .A3(new_n1063), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1065), .A2(new_n737), .A3(new_n1030), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n737), .A2(new_n1030), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1066), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n1064), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1026), .B1(new_n1050), .B2(new_n1071), .ZN(G387));
  NAND3_X1  g0872(.A1(new_n1044), .A2(new_n788), .A3(new_n1045), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n744), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(KEYINPUT109), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT109), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1073), .A2(new_n1076), .A3(new_n744), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1046), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1075), .B(new_n1077), .C1(new_n788), .C2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n727), .A2(new_n848), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n234), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1081), .A2(new_n432), .A3(new_n851), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n612), .A2(G116), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n268), .B1(new_n300), .B2(new_n256), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n291), .A2(KEYINPUT50), .A3(new_n287), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT50), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n326), .B2(G50), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1083), .B1(new_n1088), .B2(new_n254), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n743), .B1(new_n1082), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n849), .B1(new_n205), .B2(new_n345), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n793), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n842), .A2(new_n291), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n806), .A2(new_n256), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1012), .B(new_n1094), .C1(G159), .C2(new_n799), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n254), .B1(new_n811), .B2(new_n300), .C1(new_n287), .C2(new_n814), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G150), .B2(new_n820), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n838), .A2(new_n334), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1093), .A2(new_n1095), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n831), .A2(G317), .B1(new_n832), .B2(G303), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1100), .B1(new_n813), .B2(new_n800), .C1(new_n828), .C2(new_n812), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT48), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n838), .A2(G283), .B1(new_n660), .B2(new_n807), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT49), .Z(new_n1107));
  INV_X1    g0907(.A(new_n820), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n432), .B1(new_n510), .B2(new_n804), .C1(new_n1108), .C2(new_n801), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1099), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1092), .B1(new_n1110), .B2(new_n795), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1078), .A2(new_n792), .B1(new_n1080), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1079), .A2(new_n1112), .ZN(G393));
  NOR2_X1   g0913(.A1(new_n997), .A2(new_n248), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n849), .B1(new_n205), .B2(new_n217), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n793), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(G159), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n800), .A2(new_n893), .B1(new_n1117), .B2(new_n814), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT51), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1118), .A2(new_n1119), .B1(G77), .B2(new_n838), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n1119), .B2(new_n1118), .C1(new_n287), .C2(new_n828), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n432), .B(new_n886), .C1(new_n291), .C2(new_n832), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n300), .B2(new_n806), .C1(new_n1001), .C2(new_n1108), .ZN(new_n1123));
  AOI211_X1 g0923(.A(new_n254), .B(new_n840), .C1(G294), .C2(new_n832), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n802), .B2(new_n806), .C1(new_n813), .C2(new_n1108), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n799), .A2(G317), .B1(G311), .B2(new_n831), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n842), .A2(G303), .B1(G116), .B2(new_n838), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n1121), .A2(new_n1123), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1116), .B1(new_n1131), .B2(new_n795), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1030), .B2(new_n856), .ZN(new_n1133));
  AND2_X1   g0933(.A1(new_n1040), .A2(new_n1073), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n744), .B1(new_n1040), .B2(new_n1073), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1133), .B1(new_n791), .B2(new_n1040), .C1(new_n1134), .C2(new_n1135), .ZN(G390));
  INV_X1    g0936(.A(new_n744), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n979), .A2(new_n980), .A3(G330), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT111), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT111), .A4(G330), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n946), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n945), .A2(new_n958), .B1(new_n972), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n874), .B(new_n721), .C1(new_n756), .C2(new_n757), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n966), .B1(new_n1145), .B2(new_n868), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n490), .A2(new_n951), .B1(new_n954), .B2(new_n923), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n944), .B1(new_n1147), .B2(KEYINPUT38), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1146), .A2(new_n1148), .A3(new_n946), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1142), .B1(new_n1144), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g0950(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT39), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT39), .B1(new_n956), .B2(new_n985), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1151), .A2(new_n1152), .B1(new_n967), .B2(new_n946), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1145), .A2(new_n868), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1143), .B(new_n986), .C1(new_n1154), .C2(new_n966), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n971), .A2(G330), .A3(new_n786), .A4(new_n874), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1150), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n979), .A2(G330), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n975), .B(new_n695), .C1(new_n492), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(KEYINPUT112), .ZN(new_n1162));
  INV_X1    g0962(.A(KEYINPUT112), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n979), .A2(new_n1163), .A3(G330), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n874), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n966), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1156), .A2(new_n1154), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n786), .A2(G330), .A3(new_n874), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n966), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1140), .A2(new_n1171), .A3(new_n1141), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n970), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1161), .B1(new_n1169), .B2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1137), .B1(new_n1159), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n875), .B1(new_n1160), .B2(KEYINPUT112), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n971), .B1(new_n1176), .B2(new_n1164), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1173), .B1(new_n1177), .B2(new_n1167), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1161), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1180), .A2(KEYINPUT113), .A3(new_n1158), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT113), .B1(new_n1180), .B2(new_n1158), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1159), .A2(new_n792), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n846), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n793), .B1(new_n291), .B2(new_n882), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n432), .B1(new_n814), .B2(new_n510), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n800), .A2(new_n802), .B1(new_n215), .B2(new_n806), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(G97), .C2(new_n832), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n256), .B2(new_n824), .C1(new_n345), .C2(new_n828), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n804), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n820), .A2(G294), .B1(new_n1191), .B2(G68), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT114), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT54), .B(G143), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n254), .B1(new_n811), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n799), .A2(G128), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n287), .B2(new_n804), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G132), .C2(new_n831), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n892), .B2(new_n828), .C1(new_n1117), .C2(new_n824), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n820), .A2(G125), .ZN(new_n1200));
  OR3_X1    g1000(.A1(new_n806), .A2(KEYINPUT53), .A3(new_n893), .ZN(new_n1201));
  OAI21_X1  g1001(.A(KEYINPUT53), .B1(new_n806), .B2(new_n893), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1190), .A2(new_n1193), .B1(new_n1199), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1186), .B1(new_n1204), .B2(new_n795), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1185), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1183), .A2(new_n1184), .A3(new_n1206), .ZN(G378));
  NAND2_X1  g1007(.A1(new_n432), .A2(new_n267), .ZN(new_n1208));
  AOI211_X1 g1008(.A(new_n1208), .B(new_n1094), .C1(G58), .C2(new_n1191), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n802), .B2(new_n1108), .ZN(new_n1210));
  XOR2_X1   g1010(.A(new_n1210), .B(KEYINPUT115), .Z(new_n1211));
  NAND2_X1  g1011(.A1(new_n334), .A2(new_n832), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n799), .A2(G116), .B1(G107), .B2(new_n831), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1007), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1211), .B(new_n1214), .C1(new_n217), .C2(new_n828), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT58), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1208), .B(new_n287), .C1(G33), .C2(G41), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n838), .A2(G150), .B1(G125), .B2(new_n799), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT117), .ZN(new_n1222));
  INV_X1    g1022(.A(G128), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n806), .A2(new_n1194), .B1(new_n814), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT116), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n842), .A2(G132), .B1(G137), .B2(new_n832), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1222), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n293), .B(new_n267), .C1(new_n804), .C2(new_n1117), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1227), .A2(KEYINPUT59), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1229), .B(new_n1230), .C1(G124), .C2(new_n820), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1220), .B1(new_n1228), .B2(new_n1231), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n796), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n794), .B(new_n1233), .C1(new_n287), .C2(new_n881), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n305), .A2(new_n718), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n317), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1235), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n312), .A2(new_n313), .A3(new_n316), .A4(new_n1237), .ZN(new_n1238));
  XNOR2_X1  g1038(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1239), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n846), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1234), .A2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n987), .A2(new_n986), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n979), .A2(new_n980), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n956), .B2(new_n957), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(G330), .C1(new_n1248), .C2(KEYINPUT40), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n1242), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT40), .B1(new_n981), .B2(new_n961), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1242), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1252), .A2(G330), .A3(new_n1246), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n959), .A2(new_n960), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n969), .A2(new_n973), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1250), .A2(new_n1254), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1250), .A2(new_n1257), .A3(new_n1256), .A4(new_n1254), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1245), .B1(new_n1261), .B2(new_n792), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT118), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1178), .A2(new_n1157), .A3(new_n1150), .A4(new_n1179), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n1179), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1166), .A2(new_n1168), .B1(new_n1172), .B2(new_n970), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1264), .B(new_n1179), .C1(new_n1158), .C2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1261), .B1(new_n1266), .B2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT57), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1137), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1253), .B1(new_n988), .B2(G330), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT40), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1148), .A2(new_n1274), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1251), .A2(new_n1275), .A3(new_n735), .A4(new_n1242), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1273), .A2(new_n1276), .A3(new_n974), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT119), .B1(new_n1277), .B2(new_n1258), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT119), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1260), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1179), .B1(new_n1158), .B2(new_n1267), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(KEYINPUT118), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1268), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1281), .A2(new_n1284), .A3(KEYINPUT57), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1263), .B1(new_n1272), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(G375));
  NAND2_X1  g1087(.A1(new_n1267), .A2(new_n1161), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1180), .A2(new_n1288), .A3(new_n1049), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n966), .A2(new_n846), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n793), .B1(G68), .B2(new_n882), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n842), .A2(G116), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n804), .A2(new_n256), .B1(new_n806), .B2(new_n217), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1293), .B1(G294), .B2(new_n799), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n432), .B1(new_n811), .B2(new_n345), .C1(new_n802), .C2(new_n814), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(G303), .B2(new_n820), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1292), .A2(new_n1098), .A3(new_n1294), .A4(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n432), .B1(new_n832), .B2(G150), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n1298), .B1(new_n299), .B2(new_n804), .C1(new_n1117), .C2(new_n806), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(G128), .B2(new_n820), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n799), .A2(G132), .B1(G137), .B2(new_n831), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n828), .B2(new_n1194), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT120), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n838), .A2(G50), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1300), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1297), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1291), .B1(new_n1308), .B2(new_n795), .ZN(new_n1309));
  XNOR2_X1  g1109(.A(new_n1309), .B(KEYINPUT121), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(new_n1310), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1311), .B1(new_n1267), .B2(new_n791), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1289), .A2(new_n1313), .ZN(G381));
  INV_X1    g1114(.A(G378), .ZN(new_n1315));
  NOR3_X1   g1115(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(G396), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1079), .A2(new_n1318), .A3(new_n1112), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n904), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT122), .ZN(new_n1321));
  OR2_X1    g1121(.A1(new_n1320), .A2(KEYINPUT122), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1317), .A2(new_n1286), .A3(new_n1321), .A4(new_n1322), .ZN(G407));
  NAND2_X1  g1123(.A1(new_n719), .A2(G213), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1286), .A2(new_n1315), .A3(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(G407), .A2(G213), .A3(new_n1326), .ZN(G409));
  AOI22_X1  g1127(.A1(new_n1283), .A2(new_n1268), .B1(new_n1260), .B2(new_n1259), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n744), .B1(new_n1328), .B2(KEYINPUT57), .ZN(new_n1329));
  AND3_X1   g1129(.A1(new_n1281), .A2(new_n1284), .A3(KEYINPUT57), .ZN(new_n1330));
  OAI211_X1 g1130(.A(G378), .B(new_n1262), .C1(new_n1329), .C2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1049), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1245), .B1(new_n1281), .B2(new_n792), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1315), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1331), .A2(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(new_n1324), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1325), .A2(G2897), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1169), .A2(KEYINPUT60), .A3(new_n1173), .A4(new_n1161), .ZN(new_n1340));
  AND2_X1   g1140(.A1(new_n1340), .A2(new_n744), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT60), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1288), .B1(new_n1174), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1341), .A2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(G384), .B1(new_n1344), .B2(new_n1313), .ZN(new_n1345));
  AOI211_X1 g1145(.A(new_n904), .B(new_n1312), .C1(new_n1341), .C2(new_n1343), .ZN(new_n1346));
  OAI21_X1  g1146(.A(KEYINPUT124), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1340), .A2(new_n744), .ZN(new_n1348));
  OAI21_X1  g1148(.A(KEYINPUT60), .B1(new_n1267), .B2(new_n1161), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1348), .B1(new_n1288), .B2(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n904), .B1(new_n1350), .B2(new_n1312), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1344), .A2(G384), .A3(new_n1313), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT124), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1351), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  AOI21_X1  g1154(.A(new_n1339), .B1(new_n1347), .B2(new_n1354), .ZN(new_n1355));
  NOR2_X1   g1155(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1338), .B1(new_n1356), .B2(new_n1353), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1355), .A2(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(KEYINPUT61), .B1(new_n1337), .B2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1325), .B1(new_n1331), .B2(new_n1335), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT62), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1360), .A2(new_n1361), .A3(new_n1356), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1336), .A2(new_n1324), .A3(new_n1356), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1363), .A2(KEYINPUT62), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1359), .A2(new_n1362), .A3(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n788), .ZN(new_n1366));
  AND2_X1   g1166(.A1(new_n1039), .A2(new_n737), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1039), .A2(new_n737), .ZN(new_n1368));
  NOR2_X1   g1168(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1366), .B1(new_n1369), .B2(new_n1078), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n791), .B1(new_n1370), .B2(new_n1048), .ZN(new_n1371));
  INV_X1    g1171(.A(new_n1071), .ZN(new_n1372));
  AOI22_X1  g1172(.A1(new_n1371), .A2(new_n1372), .B1(new_n1025), .B2(new_n1020), .ZN(new_n1373));
  AOI21_X1  g1173(.A(new_n1318), .B1(new_n1079), .B2(new_n1112), .ZN(new_n1374));
  OAI22_X1  g1174(.A1(new_n1373), .A2(KEYINPUT125), .B1(new_n1319), .B2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(G393), .A2(G396), .ZN(new_n1376));
  NAND3_X1  g1176(.A1(new_n1079), .A2(new_n1318), .A3(new_n1112), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1376), .A2(G387), .A3(new_n1377), .ZN(new_n1378));
  AND3_X1   g1178(.A1(new_n1375), .A2(G390), .A3(new_n1378), .ZN(new_n1379));
  AOI21_X1  g1179(.A(G390), .B1(new_n1375), .B2(new_n1378), .ZN(new_n1380));
  NOR2_X1   g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1365), .A2(new_n1381), .ZN(new_n1382));
  XOR2_X1   g1182(.A(KEYINPUT123), .B(KEYINPUT63), .Z(new_n1383));
  NAND2_X1  g1183(.A1(new_n1363), .A2(new_n1383), .ZN(new_n1384));
  AND2_X1   g1184(.A1(new_n1356), .A2(KEYINPUT63), .ZN(new_n1385));
  AOI21_X1  g1185(.A(new_n1381), .B1(new_n1360), .B2(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT61), .ZN(new_n1387));
  AOI21_X1  g1187(.A(G378), .B1(new_n1332), .B2(new_n1333), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1388), .B1(new_n1286), .B2(G378), .ZN(new_n1389));
  OAI21_X1  g1189(.A(new_n1358), .B1(new_n1389), .B2(new_n1325), .ZN(new_n1390));
  NAND4_X1  g1190(.A1(new_n1384), .A2(new_n1386), .A3(new_n1387), .A4(new_n1390), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT126), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1391), .A2(new_n1392), .ZN(new_n1393));
  NAND4_X1  g1193(.A1(new_n1359), .A2(new_n1384), .A3(KEYINPUT126), .A4(new_n1386), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1382), .A2(new_n1393), .A3(new_n1394), .ZN(G405));
  INV_X1    g1195(.A(new_n1356), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1396), .A2(KEYINPUT127), .ZN(new_n1397));
  XOR2_X1   g1197(.A(new_n1381), .B(new_n1397), .Z(new_n1398));
  OAI21_X1  g1198(.A(new_n1331), .B1(KEYINPUT127), .B2(new_n1396), .ZN(new_n1399));
  AOI21_X1  g1199(.A(new_n1399), .B1(new_n1315), .B2(G375), .ZN(new_n1400));
  XNOR2_X1  g1200(.A(new_n1398), .B(new_n1400), .ZN(G402));
endmodule


