//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n507, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G125), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n470), .A2(new_n474), .ZN(G160));
  OAI211_X1 g050(.A(G124), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT67), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT68), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G112), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n479), .B1(new_n480), .B2(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(new_n468), .B2(G136), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n477), .A2(new_n478), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n478), .B1(new_n477), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(G162));
  INV_X1    g061(.A(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n487), .C1(new_n465), .C2(new_n466), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n487), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G543), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(new_n500), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(G166));
  INV_X1    g081(.A(KEYINPUT69), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n501), .A2(KEYINPUT69), .A3(new_n502), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(new_n511), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n510), .A2(new_n511), .A3(new_n514), .A4(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n516), .A2(G51), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(KEYINPUT6), .B(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n497), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G89), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n519), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n517), .A2(new_n524), .ZN(G168));
  NAND2_X1  g100(.A1(new_n516), .A2(G52), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n500), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n530), .A2(new_n531), .B1(new_n501), .B2(new_n502), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G90), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n526), .A2(new_n528), .A3(new_n533), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  NAND2_X1  g110(.A1(new_n516), .A2(G43), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(G81), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  AND2_X1   g114(.A1(KEYINPUT5), .A2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n529), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n539), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n500), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OAI211_X1 g120(.A(KEYINPUT71), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n538), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT72), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND4_X1  g130(.A1(new_n510), .A2(new_n511), .A3(G53), .A4(G543), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G543), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n558), .B1(new_n521), .B2(new_n507), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n559), .A2(new_n560), .A3(G53), .A4(new_n511), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  AND2_X1   g137(.A1(G78), .A2(G543), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n497), .B2(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT74), .B1(new_n564), .B2(new_n500), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n530), .B2(new_n531), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(G651), .C1(new_n568), .C2(new_n563), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n522), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n532), .A2(KEYINPUT73), .A3(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n562), .A2(new_n570), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND3_X1  g153(.A1(new_n559), .A2(G49), .A3(new_n511), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n532), .A2(G87), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(G288));
  AOI22_X1  g157(.A1(new_n497), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n583), .A2(new_n500), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n521), .A2(G48), .A3(G543), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n532), .A2(G86), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G305));
  AOI22_X1  g164(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n590), .A2(new_n500), .B1(new_n522), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n516), .B2(G47), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(KEYINPUT75), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(KEYINPUT75), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(G54), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n513), .B2(new_n515), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n541), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  AOI21_X1  g178(.A(KEYINPUT10), .B1(new_n532), .B2(G92), .ZN(new_n604));
  AND4_X1   g179(.A1(KEYINPUT10), .A2(new_n497), .A3(new_n521), .A4(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n597), .B1(G868), .B2(new_n607), .ZN(G284));
  OAI21_X1  g183(.A(new_n597), .B1(G868), .B2(new_n607), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G168), .B2(new_n610), .ZN(G280));
  XOR2_X1   g187(.A(G280), .B(KEYINPUT76), .Z(G297));
  XNOR2_X1  g188(.A(KEYINPUT77), .B(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(G860), .B2(new_n614), .ZN(G148));
  NAND2_X1  g190(.A1(new_n548), .A2(new_n610), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n607), .A2(new_n614), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n610), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT78), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g195(.A1(new_n467), .A2(new_n487), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G123), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  INV_X1    g200(.A(G111), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G2105), .ZN(new_n627));
  AOI21_X1  g202(.A(new_n627), .B1(new_n468), .B2(G135), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT79), .B(KEYINPUT12), .ZN(new_n633));
  NOR3_X1   g208(.A1(new_n463), .A2(new_n464), .A3(G2105), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n629), .A2(G2096), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n632), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT81), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(KEYINPUT14), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n655), .A2(new_n656), .A3(G14), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT82), .Z(G401));
  INV_X1    g233(.A(KEYINPUT18), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n662), .A2(KEYINPUT17), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n660), .A2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n637), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n662), .B2(KEYINPUT18), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n631), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1971), .B(G1976), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  AND2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n673), .A2(new_n674), .ZN(new_n678));
  NOR3_X1   g253(.A1(new_n672), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n672), .B2(new_n678), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(G229));
  XNOR2_X1  g262(.A(KEYINPUT31), .B(G11), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT30), .B(G28), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n688), .B(new_n691), .C1(new_n629), .C2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G16), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G21), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G168), .B2(new_n693), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n692), .B1(new_n695), .B2(G1966), .ZN(new_n696));
  NOR2_X1   g271(.A1(G171), .A2(new_n693), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G5), .B2(new_n693), .ZN(new_n698));
  INV_X1    g273(.A(G1961), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n696), .B1(G1966), .B2(new_n695), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT94), .Z(new_n701));
  NOR2_X1   g276(.A1(G29), .A2(G32), .ZN(new_n702));
  AOI22_X1  g277(.A1(new_n468), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT26), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  AOI22_X1  g282(.A1(new_n621), .A2(G129), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(KEYINPUT92), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n703), .A2(new_n708), .A3(KEYINPUT92), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(KEYINPUT93), .A3(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n713));
  INV_X1    g288(.A(new_n711), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(new_n709), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n702), .B1(new_n717), .B2(G29), .ZN(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT27), .B(G1996), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n693), .A2(G4), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n607), .B2(new_n693), .ZN(new_n722));
  INV_X1    g297(.A(G1348), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n693), .A2(G20), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT23), .Z(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G299), .B2(G16), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1956), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n720), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n690), .A2(G33), .ZN(new_n730));
  AND3_X1   g305(.A1(new_n468), .A2(KEYINPUT89), .A3(G139), .ZN(new_n731));
  AOI21_X1  g306(.A(KEYINPUT89), .B1(new_n468), .B2(G139), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n487), .A2(G103), .A3(G2104), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT25), .Z(new_n735));
  INV_X1    g310(.A(new_n467), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n736), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n735), .B1(new_n737), .B2(new_n487), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(new_n690), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G2072), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n690), .B1(new_n742), .B2(G34), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT90), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n742), .A2(G34), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT91), .Z(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G160), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2084), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n690), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n690), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2078), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n690), .A2(G26), .ZN(new_n754));
  XOR2_X1   g329(.A(new_n754), .B(KEYINPUT28), .Z(new_n755));
  NAND2_X1  g330(.A1(new_n468), .A2(G140), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n621), .A2(G128), .ZN(new_n757));
  OR2_X1    g332(.A1(G104), .A2(G2105), .ZN(new_n758));
  OAI211_X1 g333(.A(new_n758), .B(G2104), .C1(G116), .C2(new_n487), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n755), .B1(new_n760), .B2(G29), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR4_X1   g338(.A1(new_n741), .A2(new_n750), .A3(new_n753), .A4(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G29), .A2(G35), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G162), .B2(G29), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT29), .B(G2090), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n766), .A2(new_n767), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n699), .B2(new_n698), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n549), .B2(G16), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(G1341), .Z(new_n773));
  NAND4_X1  g348(.A1(new_n764), .A2(new_n768), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NOR3_X1   g349(.A1(new_n701), .A2(new_n729), .A3(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT34), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n693), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n693), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT86), .Z(new_n780));
  INV_X1    g355(.A(G1971), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G23), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT85), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G288), .B2(new_n693), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT33), .B(G1976), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n782), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n693), .A2(G6), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n588), .B2(new_n693), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT84), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(KEYINPUT32), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n793), .A2(G1981), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(G1981), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n777), .B(new_n789), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n693), .A2(G24), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n594), .A2(new_n595), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n693), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(G1986), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(G1986), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n690), .A2(G25), .ZN(new_n803));
  OAI211_X1 g378(.A(G131), .B(new_n487), .C1(new_n465), .C2(new_n466), .ZN(new_n804));
  OAI211_X1 g379(.A(G119), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(new_n487), .B2(G107), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT83), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n808), .A2(G95), .A3(G2105), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(G95), .B2(G2105), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n807), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n803), .B1(new_n812), .B2(new_n690), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT35), .B(G1991), .Z(new_n814));
  XOR2_X1   g389(.A(new_n813), .B(new_n814), .Z(new_n815));
  NOR3_X1   g390(.A1(new_n801), .A2(new_n802), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n797), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(KEYINPUT87), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n797), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT88), .B(KEYINPUT36), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n821), .A2(new_n823), .A3(new_n825), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n776), .B1(new_n827), .B2(new_n828), .ZN(G311));
  INV_X1    g404(.A(new_n828), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n825), .B1(new_n821), .B2(new_n823), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n775), .B1(new_n830), .B2(new_n831), .ZN(G150));
  INV_X1    g407(.A(G55), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n513), .B2(new_n515), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n541), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n837), .A2(G651), .B1(new_n532), .B2(G93), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n607), .A2(G559), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT38), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n543), .A2(new_n544), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n546), .A3(G651), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n537), .ZN(new_n848));
  INV_X1    g423(.A(G43), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(new_n513), .B2(new_n515), .ZN(new_n850));
  OAI22_X1  g425(.A1(new_n848), .A2(new_n850), .B1(new_n834), .B2(new_n839), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n514), .B1(new_n559), .B2(new_n511), .ZN(new_n852));
  INV_X1    g427(.A(new_n515), .ZN(new_n853));
  OAI21_X1  g428(.A(G55), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n536), .A2(new_n547), .A3(new_n854), .A4(new_n838), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n845), .B(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT95), .Z(new_n860));
  OAI21_X1  g435(.A(new_n841), .B1(new_n857), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n843), .B1(new_n860), .B2(new_n861), .ZN(G145));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n739), .A2(new_n714), .A3(new_n709), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n716), .B2(new_n739), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n812), .A2(KEYINPUT98), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT98), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n806), .B2(new_n811), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n468), .A2(G142), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n621), .A2(G130), .ZN(new_n871));
  OR2_X1    g446(.A1(G106), .A2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n872), .B(G2104), .C1(G118), .C2(new_n487), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n866), .A2(new_n874), .A3(new_n868), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n493), .A2(KEYINPUT97), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n493), .A2(KEYINPUT97), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n489), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n760), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n760), .A2(new_n880), .A3(new_n489), .A4(new_n881), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n635), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n884), .A2(new_n635), .A3(new_n885), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n879), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n884), .A2(new_n635), .A3(new_n885), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n890), .A2(new_n886), .A3(new_n878), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n865), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT93), .B1(new_n710), .B2(new_n711), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n714), .A2(new_n713), .A3(new_n709), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n739), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n864), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n887), .A2(new_n879), .A3(new_n888), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n878), .B1(new_n890), .B2(new_n886), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n470), .A2(new_n474), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n484), .B2(new_n485), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n477), .A2(new_n482), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT68), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n905), .A2(G160), .A3(new_n483), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT96), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n903), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n629), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n484), .A2(new_n485), .A3(new_n902), .ZN(new_n911));
  AOI21_X1  g486(.A(G160), .B1(new_n905), .B2(new_n483), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT96), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n903), .A2(new_n906), .A3(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(new_n630), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n910), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n908), .A2(new_n909), .A3(new_n629), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n630), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT99), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n901), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT100), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n901), .A2(new_n920), .A3(KEYINPUT100), .A4(new_n917), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n910), .A2(new_n915), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n892), .A3(new_n900), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n863), .B1(new_n925), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI211_X1 g507(.A(KEYINPUT101), .B(new_n929), .C1(new_n923), .C2(new_n924), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g511(.A1(new_n799), .A2(G305), .ZN(new_n937));
  INV_X1    g512(.A(G288), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(G166), .ZN(new_n939));
  NAND2_X1  g514(.A1(G290), .A2(new_n588), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n937), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n939), .B1(new_n937), .B2(new_n940), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT42), .Z(new_n944));
  INV_X1    g519(.A(KEYINPUT104), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n856), .B(new_n617), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n607), .A2(G299), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n565), .A2(new_n569), .B1(new_n573), .B2(new_n574), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n949), .B(new_n562), .C1(new_n599), .C2(new_n606), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT41), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT102), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n948), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n599), .A2(new_n606), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n562), .A2(new_n570), .A3(new_n575), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT102), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n954), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n951), .B2(new_n954), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT103), .A4(KEYINPUT41), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n953), .B1(new_n947), .B2(new_n964), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n946), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n944), .A2(new_n945), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n967), .B1(new_n946), .B2(new_n965), .ZN(new_n968));
  OAI21_X1  g543(.A(G868), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G868), .B2(new_n840), .ZN(G295));
  OAI21_X1  g545(.A(new_n969), .B1(G868), .B2(new_n840), .ZN(G331));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT106), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n856), .A2(G171), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n851), .A2(new_n855), .A3(G301), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(G168), .A3(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n851), .A2(new_n855), .A3(G301), .ZN(new_n977));
  AOI21_X1  g552(.A(G301), .B1(new_n851), .B2(new_n855), .ZN(new_n978));
  OAI21_X1  g553(.A(G286), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n964), .A2(new_n973), .A3(new_n976), .A4(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n976), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(new_n951), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n979), .A2(new_n976), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n973), .B1(new_n984), .B2(new_n964), .ZN(new_n985));
  OR3_X1    g560(.A1(new_n983), .A2(new_n985), .A3(new_n943), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n988));
  AND3_X1   g563(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT106), .B1(new_n989), .B2(new_n981), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n990), .A2(new_n982), .A3(new_n980), .ZN(new_n991));
  AOI211_X1 g566(.A(new_n988), .B(G37), .C1(new_n991), .C2(new_n943), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n943), .B1(new_n983), .B2(new_n985), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT107), .B1(new_n993), .B2(new_n928), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n986), .B(new_n987), .C1(new_n992), .C2(new_n994), .ZN(new_n995));
  OR2_X1    g570(.A1(new_n956), .A2(new_n959), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n984), .A2(KEYINPUT41), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n943), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n952), .B1(new_n981), .B2(new_n954), .ZN(new_n999));
  AOI21_X1  g574(.A(G37), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n986), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT43), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n972), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n1000), .A2(new_n986), .A3(new_n987), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n986), .B1(new_n992), .B2(new_n994), .ZN(new_n1005));
  INV_X1    g580(.A(new_n987), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1003), .B1(new_n972), .B2(new_n1007), .ZN(G397));
  NOR2_X1   g583(.A1(G290), .A2(G1986), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G160), .A2(new_n1011), .A3(G40), .ZN(new_n1012));
  INV_X1    g587(.A(G40), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT109), .B1(new_n902), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n882), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n1017), .B2(KEYINPUT108), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(KEYINPUT108), .B2(new_n1017), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1010), .A2(new_n1015), .A3(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1019), .A2(new_n1015), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n760), .B(G2067), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n714), .A2(new_n709), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(G1996), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(G1996), .B2(new_n716), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n812), .B(new_n814), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1022), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1021), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n812), .A2(new_n814), .ZN(new_n1032));
  OAI22_X1  g607(.A1(new_n1027), .A2(new_n1032), .B1(G2067), .B2(new_n760), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1022), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  OR3_X1    g610(.A1(new_n1019), .A2(G1996), .A3(new_n1015), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT126), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1022), .B1(new_n1025), .B2(new_n1023), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1042), .A2(KEYINPUT47), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1035), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  INV_X1    g624(.A(G1981), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n586), .A2(new_n1050), .A3(new_n587), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT113), .B(G86), .Z(new_n1052));
  OAI211_X1 g627(.A(new_n584), .B(new_n585), .C1(new_n522), .C2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G1981), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1051), .A2(new_n1054), .A3(KEYINPUT49), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT49), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1048), .A2(new_n1049), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1057), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n882), .A2(new_n1016), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1014), .A3(new_n1012), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(new_n1062), .A3(G8), .A4(new_n1055), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT114), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1059), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n938), .A2(G1976), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(G8), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT112), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1062), .A2(new_n1069), .A3(G8), .A4(new_n1066), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(KEYINPUT52), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(G1976), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT52), .B1(G288), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1067), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1065), .A2(new_n1071), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n495), .A2(new_n1016), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT45), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(new_n1014), .A3(new_n1012), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1017), .A2(new_n1079), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n781), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1061), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2090), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1078), .A2(KEYINPUT50), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G166), .A2(new_n1047), .ZN(new_n1091));
  NOR2_X1   g666(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1092));
  AND2_X1   g667(.A1(KEYINPUT111), .A2(KEYINPUT55), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(G8), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n495), .A2(new_n1085), .A3(new_n1016), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1084), .A2(new_n1087), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1047), .B1(new_n1083), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1096), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(KEYINPUT125), .B1(new_n1077), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1083), .A2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1095), .B1(new_n1103), .B2(G8), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1095), .A2(G8), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1075), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1071), .A4(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT117), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1088), .A2(new_n1014), .A3(new_n1012), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1084), .A2(new_n1086), .A3(KEYINPUT117), .A4(new_n1088), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1114), .A2(new_n1115), .A3(new_n699), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT53), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1061), .A2(KEYINPUT45), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1084), .A2(new_n1118), .A3(new_n1080), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1119), .B2(G2078), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1012), .B(new_n1014), .C1(new_n1079), .C2(new_n1078), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1061), .A2(KEYINPUT45), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1117), .A2(G2078), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1116), .B(new_n1120), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1125), .A2(G171), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1102), .A2(new_n1110), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1966), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1129));
  INV_X1    g704(.A(G2084), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1084), .A2(new_n1086), .A3(new_n1130), .A4(new_n1088), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(G168), .A2(new_n1047), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT123), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1047), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1135), .B(KEYINPUT51), .C1(new_n1136), .C2(new_n1134), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1136), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1134), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1138), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1137), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT62), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT124), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1137), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1127), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1136), .A2(new_n1152), .A3(G168), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1096), .B1(new_n1153), .B2(new_n1104), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(new_n1071), .A3(new_n1109), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1136), .B(G168), .C1(new_n1090), .C2(new_n1095), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT63), .B1(new_n1077), .B2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g732(.A(G1976), .B(G288), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1051), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1048), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1155), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1151), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(G301), .B(KEYINPUT54), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1082), .A2(new_n1013), .A3(new_n902), .A4(new_n1124), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1163), .B1(new_n1165), .B2(new_n1019), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1125), .A2(new_n1163), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1102), .A2(new_n1110), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n562), .A2(KEYINPUT115), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n562), .A2(KEYINPUT115), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n949), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT57), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT116), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n958), .A2(KEYINPUT57), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1173), .A2(KEYINPUT116), .A3(new_n1174), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(KEYINPUT56), .B(G2072), .ZN(new_n1181));
  NAND4_X1  g756(.A1(new_n1084), .A2(new_n1118), .A3(new_n1080), .A4(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1084), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1183));
  INV_X1    g758(.A(G1956), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1180), .A2(new_n1182), .A3(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1114), .A2(new_n1115), .A3(new_n723), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1046), .A2(new_n762), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n957), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT118), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1185), .A2(new_n1182), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1192), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1186), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1197), .A2(new_n607), .ZN(new_n1198));
  OAI21_X1  g773(.A(KEYINPUT60), .B1(new_n1198), .B2(new_n1189), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT121), .ZN(new_n1200));
  XOR2_X1   g775(.A(KEYINPUT119), .B(G1996), .Z(new_n1201));
  NAND4_X1  g776(.A1(new_n1084), .A2(new_n1118), .A3(new_n1080), .A4(new_n1201), .ZN(new_n1202));
  XOR2_X1   g777(.A(KEYINPUT58), .B(G1341), .Z(new_n1203));
  NAND2_X1  g778(.A1(new_n1062), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n548), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT59), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1200), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT120), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  OAI21_X1  g785(.A(KEYINPUT59), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1207), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1213), .A2(new_n549), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1206), .B1(new_n1214), .B2(KEYINPUT120), .ZN(new_n1215));
  NAND3_X1  g790(.A1(new_n1215), .A2(new_n1200), .A3(new_n1209), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1193), .A2(KEYINPUT61), .A3(new_n1186), .ZN(new_n1217));
  NAND4_X1  g792(.A1(new_n1199), .A2(new_n1212), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  AND2_X1   g793(.A1(new_n1193), .A2(new_n1186), .ZN(new_n1219));
  OR2_X1    g794(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n1220));
  OAI22_X1  g795(.A1(new_n1219), .A2(KEYINPUT61), .B1(new_n1197), .B2(new_n1220), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1196), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1170), .B1(KEYINPUT122), .B2(new_n1222), .ZN(new_n1223));
  OR2_X1    g798(.A1(new_n1222), .A2(KEYINPUT122), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1162), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(G290), .A2(G1986), .ZN(new_n1226));
  AND3_X1   g801(.A1(new_n1010), .A2(KEYINPUT110), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g802(.A(new_n1022), .B1(KEYINPUT110), .B2(new_n1226), .ZN(new_n1228));
  OAI21_X1  g803(.A(new_n1029), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g804(.A(new_n1045), .B1(new_n1225), .B2(new_n1229), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g805(.A(new_n1004), .ZN(new_n1232));
  INV_X1    g806(.A(new_n986), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n928), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n1234), .A2(new_n988), .ZN(new_n1235));
  NAND3_X1  g809(.A1(new_n993), .A2(KEYINPUT107), .A3(new_n928), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  OAI21_X1  g811(.A(new_n1232), .B1(new_n1237), .B2(new_n987), .ZN(new_n1238));
  OR3_X1    g812(.A1(new_n657), .A2(new_n461), .A3(G227), .ZN(new_n1239));
  OR2_X1    g813(.A1(G229), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g814(.A(new_n1240), .B1(new_n932), .B2(new_n934), .ZN(new_n1241));
  AOI21_X1  g815(.A(KEYINPUT127), .B1(new_n1238), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1243));
  NOR2_X1   g817(.A1(G229), .A2(new_n1239), .ZN(new_n1244));
  OAI21_X1  g818(.A(new_n1244), .B1(new_n931), .B2(new_n933), .ZN(new_n1245));
  NOR3_X1   g819(.A1(new_n1007), .A2(new_n1243), .A3(new_n1245), .ZN(new_n1246));
  NOR2_X1   g820(.A1(new_n1242), .A2(new_n1246), .ZN(G308));
  NAND3_X1  g821(.A1(new_n1238), .A2(new_n1241), .A3(KEYINPUT127), .ZN(new_n1248));
  OAI21_X1  g822(.A(new_n1243), .B1(new_n1007), .B2(new_n1245), .ZN(new_n1249));
  NAND2_X1  g823(.A1(new_n1248), .A2(new_n1249), .ZN(G225));
endmodule


