//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  INV_X1    g000(.A(G169gat), .ZN(new_n202));
  INV_X1    g001(.A(G176gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT23), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G169gat), .B2(G176gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  AND4_X1   g006(.A1(KEYINPUT25), .A2(new_n204), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT24), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(G183gat), .A3(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n214));
  OR3_X1    g013(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n208), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  INV_X1    g017(.A(G183gat), .ZN(new_n219));
  INV_X1    g018(.A(G190gat), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n210), .A2(new_n212), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n218), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n203), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(KEYINPUT66), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  NOR2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n202), .A3(new_n203), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(KEYINPUT67), .A3(new_n225), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n228), .A2(new_n232), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n219), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(new_n220), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n242), .A2(KEYINPUT65), .ZN(new_n243));
  AOI22_X1  g042(.A1(new_n241), .A2(new_n243), .B1(G183gat), .B2(G190gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT27), .B(G183gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n245), .A2(new_n246), .A3(new_n220), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n237), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n224), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT75), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n224), .A2(KEYINPUT75), .A3(new_n248), .ZN(new_n252));
  NAND2_X1  g051(.A1(G226gat), .A2(G233gat), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(KEYINPUT29), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n258));
  XOR2_X1   g057(.A(G197gat), .B(G204gat), .Z(new_n259));
  AOI21_X1  g058(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(G197gat), .ZN(new_n262));
  INV_X1    g061(.A(G204gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G197gat), .A2(G204gat), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n260), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n257), .B1(new_n261), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n257), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n266), .B2(KEYINPUT73), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT74), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n259), .A2(new_n258), .A3(new_n260), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n267), .A2(new_n257), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n241), .A2(new_n243), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n247), .A2(new_n279), .A3(new_n209), .ZN(new_n280));
  AOI22_X1  g079(.A1(new_n280), .A2(new_n237), .B1(new_n217), .B2(new_n223), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(new_n254), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n256), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT76), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n251), .A2(new_n252), .A3(new_n254), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT29), .B1(new_n224), .B2(new_n248), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT77), .B1(new_n287), .B2(new_n254), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n289), .B(new_n253), .C1(new_n281), .C2(KEYINPUT29), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n271), .A2(new_n277), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n286), .A2(new_n288), .A3(new_n290), .A4(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n256), .A2(KEYINPUT76), .A3(new_n278), .A4(new_n282), .ZN(new_n293));
  XNOR2_X1  g092(.A(G8gat), .B(G36gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(G64gat), .B(G92gat), .ZN(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  NAND4_X1  g095(.A1(new_n285), .A2(new_n292), .A3(new_n293), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT30), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n292), .A2(new_n293), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n299), .A2(new_n300), .A3(new_n285), .A4(new_n296), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT78), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n283), .A2(new_n284), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n292), .A2(new_n293), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n285), .A2(KEYINPUT78), .A3(new_n292), .A4(new_n293), .ZN(new_n307));
  INV_X1    g106(.A(new_n296), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n302), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT84), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT84), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n302), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n316), .B2(new_n317), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT79), .B1(new_n320), .B2(G148gat), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(new_n323), .A3(G141gat), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n321), .B(new_n324), .C1(G141gat), .C2(new_n323), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n320), .A2(G148gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n323), .A2(G141gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n315), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G155gat), .B(G162gat), .Z(new_n329));
  AOI22_X1  g128(.A1(new_n319), .A2(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n268), .B2(new_n270), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n333), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n331), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n278), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G228gat), .ZN(new_n339));
  INV_X1    g138(.A(G233gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n335), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n271), .A2(new_n277), .B1(new_n331), .B2(new_n336), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n343), .A2(new_n334), .B1(new_n339), .B2(new_n340), .ZN(new_n344));
  INV_X1    g143(.A(G22gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT83), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n342), .A2(new_n344), .A3(new_n348), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n342), .A2(new_n344), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(G22gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G78gat), .B(G106gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT31), .B(G50gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  XOR2_X1   g154(.A(new_n355), .B(KEYINPUT82), .Z(new_n356));
  AOI21_X1  g155(.A(new_n355), .B1(new_n350), .B2(G22gat), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n352), .A2(new_n356), .B1(new_n346), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G113gat), .ZN(new_n363));
  INV_X1    g162(.A(G113gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G120gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367));
  XNOR2_X1  g166(.A(G127gat), .B(G134gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n366), .B(new_n367), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G134gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G127gat), .ZN(new_n372));
  INV_X1    g171(.A(G127gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G134gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(new_n367), .ZN(new_n376));
  XNOR2_X1  g175(.A(G113gat), .B(G120gat), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(KEYINPUT1), .ZN(new_n378));
  AND2_X1   g177(.A1(new_n370), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n224), .A2(new_n379), .A3(new_n248), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT69), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT69), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n224), .A2(new_n248), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n370), .A2(new_n378), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n249), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n361), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT33), .B1(new_n386), .B2(new_n387), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(KEYINPUT70), .ZN(new_n391));
  XOR2_X1   g190(.A(G71gat), .B(G99gat), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n388), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  AOI221_X4 g194(.A(new_n361), .B1(KEYINPUT33), .B2(new_n393), .C1(new_n386), .C2(new_n387), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n386), .A2(new_n387), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n397), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n386), .A2(new_n387), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT33), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n388), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n396), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n399), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n360), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n397), .B1(new_n395), .B2(new_n396), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n405), .A3(new_n399), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n359), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n358), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G1gat), .B(G29gat), .Z(new_n412));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G57gat), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n325), .A2(new_n319), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n328), .A2(new_n329), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT3), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n336), .A3(new_n384), .ZN(new_n422));
  NAND2_X1  g221(.A1(G225gat), .A2(G233gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n420), .B2(new_n384), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n379), .A2(KEYINPUT4), .A3(new_n330), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n422), .A2(new_n423), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n423), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n420), .A2(new_n384), .ZN(new_n429));
  AOI22_X1  g228(.A1(new_n418), .A2(new_n419), .B1(new_n370), .B2(new_n378), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT5), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n426), .A2(new_n425), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(KEYINPUT5), .A3(new_n423), .A4(new_n422), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n417), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n433), .A2(new_n417), .A3(new_n435), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT6), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n446), .A2(KEYINPUT35), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n314), .A2(new_n411), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT35), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n302), .A3(new_n309), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n451), .B2(new_n411), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n352), .A2(new_n356), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n357), .A2(new_n346), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT38), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n306), .A2(KEYINPUT37), .A3(new_n307), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n285), .A2(new_n458), .A3(new_n292), .A4(new_n293), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n459), .A2(new_n308), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n286), .A2(new_n288), .A3(new_n290), .A4(new_n278), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n256), .A2(new_n291), .A3(new_n282), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n462), .A2(KEYINPUT37), .A3(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n459), .A2(new_n464), .A3(new_n456), .A4(new_n308), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n442), .A2(new_n465), .A3(new_n444), .A4(new_n297), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n455), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n313), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n312), .B1(new_n302), .B2(new_n309), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n434), .A2(new_n422), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n428), .ZN(new_n472));
  OR3_X1    g271(.A1(new_n429), .A2(new_n430), .A3(new_n428), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(KEYINPUT39), .A3(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n416), .C1(KEYINPUT39), .C2(new_n472), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT40), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n475), .A2(new_n476), .ZN(new_n478));
  NOR3_X1   g277(.A1(new_n477), .A2(new_n478), .A3(new_n443), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n467), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n481));
  OR2_X1    g280(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n408), .A2(new_n359), .A3(new_n409), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n359), .B1(new_n408), .B2(new_n409), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n450), .A2(new_n358), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n407), .A2(KEYINPUT72), .A3(KEYINPUT36), .A4(new_n410), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI22_X1  g287(.A1(new_n448), .A2(new_n452), .B1(new_n480), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  INV_X1    g289(.A(G43gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(G50gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(KEYINPUT88), .B(G43gat), .ZN(new_n495));
  INV_X1    g294(.A(G50gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT15), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(G43gat), .B2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT86), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT14), .ZN(new_n503));
  NAND2_X1  g302(.A1(G29gat), .A2(G36gat), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  INV_X1    g306(.A(G36gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT86), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n502), .A3(KEYINPUT14), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(new_n506), .A3(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n498), .A2(new_n500), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT90), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT90), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n514), .B1(new_n511), .B2(new_n500), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n513), .B(KEYINPUT17), .C1(new_n515), .C2(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT92), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n512), .A2(new_n515), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT92), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(KEYINPUT17), .A4(new_n513), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT16), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n523), .B2(G1gat), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(G1gat), .B2(new_n522), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(G8gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n518), .A2(new_n513), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT91), .B(KEYINPUT17), .Z(new_n528));
  AOI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(G229gat), .A2(G233gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n526), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n530), .A2(KEYINPUT18), .A3(new_n531), .A4(new_n532), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n527), .B(new_n526), .ZN(new_n537));
  XOR2_X1   g336(.A(new_n531), .B(KEYINPUT13), .Z(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G113gat), .B(G141gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G197gat), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT11), .B(G169gat), .Z(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT12), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n540), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n540), .B2(KEYINPUT85), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n490), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n540), .A2(KEYINPUT85), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n545), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n540), .A2(KEYINPUT85), .A3(new_n546), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(KEYINPUT93), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n489), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G232gat), .A2(G233gat), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT96), .Z(new_n557));
  INV_X1    g356(.A(KEYINPUT41), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G190gat), .B(G218gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT99), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n559), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(new_n527), .B2(new_n528), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n521), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT98), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n521), .A2(new_n577), .A3(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n557), .A2(new_n558), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n580), .B1(new_n527), .B2(new_n573), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n560), .A2(KEYINPUT99), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G134gat), .B(G162gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n581), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n588), .B1(new_n576), .B2(new_n578), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n589), .B2(new_n583), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n562), .B1(new_n587), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n590), .A3(new_n562), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XOR2_X1   g393(.A(G57gat), .B(G64gat), .Z(new_n595));
  NAND2_X1  g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G71gat), .B(G78gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n601), .B(KEYINPUT94), .Z(new_n602));
  AOI21_X1  g401(.A(new_n526), .B1(new_n602), .B2(KEYINPUT21), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT95), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n316), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n604), .B(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(new_n373), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n607), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n594), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n573), .A2(new_n601), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n573), .A2(new_n601), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n602), .A2(KEYINPUT10), .A3(new_n573), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n627), .B(KEYINPUT100), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  OAI211_X1 g432(.A(new_n630), .B(new_n633), .C1(new_n629), .C2(new_n622), .ZN(new_n634));
  INV_X1    g433(.A(new_n633), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n628), .B(KEYINPUT101), .Z(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n624), .B2(new_n625), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n629), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n635), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n619), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n555), .A2(KEYINPUT102), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT102), .B1(new_n555), .B2(new_n641), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n445), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT103), .B(G1gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1324gat));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n470), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(G8gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT16), .B(G8gat), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT42), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n653), .B1(KEYINPUT42), .B2(new_n652), .ZN(G1325gat));
  NAND2_X1  g453(.A1(new_n407), .A2(new_n410), .ZN(new_n655));
  AOI21_X1  g454(.A(G15gat), .B1(new_n648), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n485), .A2(new_n487), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(G15gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT104), .Z(new_n660));
  AOI21_X1  g459(.A(new_n656), .B1(new_n648), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n455), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  INV_X1    g463(.A(new_n640), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n617), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n594), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT105), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n555), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(new_n507), .A3(new_n446), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT45), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n480), .B2(new_n488), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n457), .A2(new_n460), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT38), .ZN(new_n676));
  AND4_X1   g475(.A1(new_n442), .A2(new_n465), .A3(new_n444), .A4(new_n297), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n358), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n311), .A2(new_n313), .A3(new_n479), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n657), .A2(new_n680), .A3(KEYINPUT106), .A4(new_n486), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n455), .B1(new_n483), .B2(new_n484), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT35), .B1(new_n682), .B2(new_n450), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n314), .A2(new_n411), .A3(new_n447), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT107), .ZN(new_n685));
  AND3_X1   g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n683), .B2(new_n684), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n674), .B(new_n681), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT108), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT107), .B1(new_n448), .B2(new_n452), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n674), .A4(new_n681), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n594), .A2(KEYINPUT44), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n689), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n593), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n591), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n489), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n666), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n547), .A2(new_n548), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(KEYINPUT109), .A3(new_n705), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n445), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n672), .B1(new_n711), .B2(new_n507), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT110), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT110), .B(new_n672), .C1(new_n711), .C2(new_n507), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(G1328gat));
  OAI21_X1  g515(.A(G36gat), .B1(new_n710), .B2(new_n314), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n669), .A2(G36gat), .A3(new_n314), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1329gat));
  OAI21_X1  g519(.A(new_n495), .B1(new_n706), .B2(new_n657), .ZN(new_n721));
  INV_X1    g520(.A(new_n655), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n669), .A2(new_n722), .A3(new_n495), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(KEYINPUT47), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n708), .A2(new_n658), .A3(new_n709), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n723), .B1(new_n726), .B2(new_n495), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g527(.A1(new_n455), .A2(G50gat), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT111), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n730), .B1(new_n670), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n669), .A2(KEYINPUT111), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT48), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n708), .A2(new_n358), .A3(new_n709), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n736), .B1(new_n737), .B2(G50gat), .ZN(new_n738));
  OAI21_X1  g537(.A(G50gat), .B1(new_n706), .B2(new_n455), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(new_n734), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(KEYINPUT112), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT48), .B1(new_n732), .B2(new_n733), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT109), .B1(new_n701), .B2(new_n705), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n707), .B(new_n704), .C1(new_n696), .C2(new_n700), .ZN(new_n745));
  NOR3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(new_n455), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(new_n496), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n739), .A2(new_n734), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT48), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n742), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n741), .A2(new_n750), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n689), .A2(new_n694), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n619), .A2(new_n703), .A3(new_n665), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT113), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n445), .ZN(new_n756));
  XOR2_X1   g555(.A(new_n756), .B(G57gat), .Z(G1332gat));
  NAND3_X1  g556(.A1(new_n752), .A2(new_n754), .A3(new_n470), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT49), .B(G64gat), .Z(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n758), .B2(new_n760), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n755), .B2(new_n657), .ZN(new_n762));
  OR2_X1    g561(.A1(new_n722), .A2(G71gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n755), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g564(.A1(new_n755), .A2(new_n455), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g566(.A1(new_n618), .A2(new_n703), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n701), .A2(new_n640), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n445), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n618), .A2(new_n594), .A3(new_n703), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n688), .A2(KEYINPUT51), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT51), .B1(new_n688), .B2(new_n771), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n446), .A2(new_n568), .A3(new_n640), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  OR4_X1    g575(.A1(G92gat), .A2(new_n774), .A3(new_n314), .A4(new_n665), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n769), .A2(new_n314), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n569), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g579(.A1(new_n769), .A2(new_n657), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT114), .B(G99gat), .Z(new_n782));
  NAND3_X1  g581(.A1(new_n655), .A2(new_n640), .A3(new_n782), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n781), .A2(new_n782), .B1(new_n774), .B2(new_n783), .ZN(G1338gat));
  OAI21_X1  g583(.A(G106gat), .B1(new_n769), .B2(new_n455), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n665), .A2(new_n455), .A3(G106gat), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  INV_X1    g589(.A(new_n636), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n626), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n635), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n626), .B2(new_n791), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n624), .A2(KEYINPUT115), .A3(new_n625), .A4(new_n636), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n790), .B1(new_n626), .B2(new_n629), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n634), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n801), .B(new_n793), .C1(new_n797), .C2(new_n798), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n540), .A2(new_n545), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n530), .A2(new_n532), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n805), .A2(new_n531), .B1(new_n537), .B2(new_n538), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n804), .B1(new_n544), .B2(new_n806), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n698), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n803), .A2(new_n703), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n640), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n698), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n617), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  OR3_X1    g611(.A1(new_n619), .A2(new_n703), .A3(new_n640), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n470), .A2(new_n445), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n411), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n554), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n816), .A2(new_n364), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n814), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n819), .A2(new_n445), .A3(new_n470), .A4(new_n682), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n703), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n818), .B1(new_n821), .B2(new_n364), .ZN(G1340gat));
  NOR3_X1   g621(.A1(new_n816), .A2(new_n362), .A3(new_n665), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n640), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n362), .ZN(G1341gat));
  NAND3_X1  g624(.A1(new_n820), .A2(new_n373), .A3(new_n618), .ZN(new_n826));
  OAI21_X1  g625(.A(G127gat), .B1(new_n816), .B2(new_n617), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1342gat));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n371), .A3(new_n698), .ZN(new_n829));
  OR2_X1    g628(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n816), .B2(new_n594), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(KEYINPUT56), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(G1343gat));
  NOR2_X1   g632(.A1(new_n819), .A2(new_n445), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n658), .A2(new_n455), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n554), .A2(new_n320), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n470), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n657), .A2(new_n815), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n814), .A2(new_n358), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n549), .A2(new_n553), .A3(new_n803), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n698), .B1(new_n846), .B2(new_n810), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n617), .B1(new_n847), .B2(new_n808), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n848), .A2(new_n813), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT57), .B1(new_n849), .B2(new_n455), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n703), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n840), .B1(new_n853), .B2(G141gat), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT58), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n320), .B1(new_n852), .B2(new_n554), .ZN(new_n856));
  XOR2_X1   g655(.A(KEYINPUT118), .B(KEYINPUT58), .Z(new_n857));
  NAND2_X1  g656(.A1(new_n834), .A2(new_n835), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n835), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n860), .A2(new_n314), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n857), .B1(new_n862), .B2(new_n836), .ZN(new_n863));
  OAI22_X1  g662(.A1(new_n854), .A2(new_n855), .B1(new_n856), .B2(new_n863), .ZN(G1344gat));
  INV_X1    g663(.A(new_n862), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n323), .A3(new_n640), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n323), .C1(new_n852), .C2(new_n640), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n455), .A2(KEYINPUT57), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n846), .A2(new_n810), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n594), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n698), .A2(new_n803), .A3(new_n807), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT120), .B1(new_n847), .B2(new_n808), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n617), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n641), .A2(new_n817), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n844), .B1(new_n814), .B2(new_n358), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n665), .B1(new_n841), .B2(KEYINPUT119), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(KEYINPUT119), .B2(new_n841), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n868), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n866), .B1(new_n867), .B2(new_n887), .ZN(G1345gat));
  OAI21_X1  g687(.A(G155gat), .B1(new_n851), .B2(new_n617), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n618), .A2(new_n316), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n862), .B2(new_n890), .ZN(G1346gat));
  AOI21_X1  g690(.A(G162gat), .B1(new_n865), .B2(new_n698), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n594), .A2(new_n317), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n852), .B2(new_n893), .ZN(G1347gat));
  NOR2_X1   g693(.A1(new_n314), .A2(new_n446), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n682), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n814), .A2(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n898), .A2(new_n202), .A3(new_n817), .ZN(new_n899));
  INV_X1    g698(.A(new_n898), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n703), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n899), .B1(new_n202), .B2(new_n901), .ZN(G1348gat));
  NOR2_X1   g701(.A1(new_n898), .A2(new_n665), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(new_n203), .ZN(G1349gat));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n905), .B2(KEYINPUT122), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n900), .A2(new_n245), .A3(new_n618), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n908));
  OAI21_X1  g707(.A(G183gat), .B1(new_n898), .B2(new_n617), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(KEYINPUT121), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n905), .A2(KEYINPUT123), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n906), .B2(new_n911), .ZN(G1350gat));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n594), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n220), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT61), .Z(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n220), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1351gat));
  NOR2_X1   g719(.A1(new_n658), .A2(new_n896), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n880), .A2(new_n882), .A3(new_n921), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n262), .A3(new_n817), .ZN(new_n923));
  INV_X1    g722(.A(new_n921), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n842), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925), .B2(new_n703), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n923), .A2(new_n926), .ZN(G1352gat));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n263), .A3(new_n640), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT62), .Z(new_n929));
  OAI21_X1  g728(.A(G204gat), .B1(new_n922), .B2(new_n665), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1353gat));
  NOR4_X1   g730(.A1(new_n879), .A2(new_n881), .A3(new_n617), .A4(new_n924), .ZN(new_n932));
  OAI21_X1  g731(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n933));
  OAI211_X1 g732(.A(KEYINPUT126), .B(KEYINPUT63), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n935));
  INV_X1    g734(.A(new_n933), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n936), .C1(new_n922), .C2(new_n617), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n617), .A2(G211gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n925), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT125), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT127), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n934), .A2(new_n937), .A3(new_n940), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1354gat));
  OAI21_X1  g744(.A(G218gat), .B1(new_n922), .B2(new_n594), .ZN(new_n946));
  INV_X1    g745(.A(G218gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n925), .A2(new_n947), .A3(new_n698), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n946), .A2(new_n948), .ZN(G1355gat));
endmodule


