//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT64), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT71), .ZN(new_n204));
  INV_X1    g003(.A(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G134gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT70), .B(G134gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(new_n205), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n204), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G113gat), .B(G120gat), .Z(new_n213));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n206), .A2(KEYINPUT70), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n206), .A2(KEYINPUT70), .ZN(new_n217));
  OAI21_X1  g016(.A(G127gat), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n215), .A2(new_n218), .A3(KEYINPUT71), .A4(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G127gat), .B(G134gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n213), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT72), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT72), .ZN(new_n224));
  INV_X1    g023(.A(new_n222), .ZN(new_n225));
  AOI211_X1 g024(.A(new_n224), .B(new_n225), .C1(new_n212), .C2(new_n219), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT68), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT24), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  INV_X1    g035(.A(G169gat), .ZN(new_n237));
  INV_X1    g036(.A(G176gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n238), .A3(KEYINPUT23), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n233), .A2(new_n234), .A3(new_n236), .A4(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n241));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(KEYINPUT23), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n244), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g045(.A(KEYINPUT67), .B(new_n230), .C1(new_n240), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n239), .A2(new_n236), .A3(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n232), .A2(KEYINPUT24), .ZN(new_n249));
  NOR2_X1   g048(.A1(G183gat), .A2(G190gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n245), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n239), .A2(new_n236), .A3(new_n234), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(new_n253), .A3(new_n233), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT67), .B1(new_n257), .B2(new_n230), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n228), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n230), .B1(new_n240), .B2(new_n246), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n262), .A2(KEYINPUT68), .A3(new_n254), .A4(new_n247), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT27), .B(G183gat), .ZN(new_n265));
  INV_X1    g064(.A(G190gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT28), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n267), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n267), .A2(new_n269), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n242), .A2(KEYINPUT26), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n234), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n242), .A2(KEYINPUT26), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n232), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n227), .B1(new_n264), .B2(new_n278), .ZN(new_n279));
  AOI211_X1 g078(.A(new_n277), .B(new_n223), .C1(new_n259), .C2(new_n263), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n203), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT32), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(KEYINPUT73), .B(G71gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(G99gat), .ZN(new_n286));
  XOR2_X1   g085(.A(G15gat), .B(G43gat), .Z(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n223), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n229), .B1(new_n252), .B2(new_n253), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n256), .A2(new_n253), .A3(new_n233), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n291), .A2(KEYINPUT67), .B1(new_n292), .B2(KEYINPUT25), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT68), .B1(new_n293), .B2(new_n262), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n255), .A2(new_n228), .A3(new_n258), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n278), .B(new_n290), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n203), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n277), .B1(new_n259), .B2(new_n263), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(new_n227), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT34), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n300), .B1(new_n297), .B2(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g101(.A1(new_n298), .A2(new_n227), .ZN(new_n303));
  INV_X1    g102(.A(new_n301), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n303), .A2(new_n297), .A3(new_n296), .A4(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n288), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n281), .B(KEYINPUT32), .C1(new_n283), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n289), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n289), .A2(new_n306), .A3(KEYINPUT76), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n306), .B1(new_n289), .B2(new_n308), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT84), .ZN(new_n317));
  XNOR2_X1  g116(.A(G197gat), .B(G204gat), .ZN(new_n318));
  INV_X1    g117(.A(G211gat), .ZN(new_n319));
  INV_X1    g118(.A(G218gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(KEYINPUT22), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G211gat), .B(G218gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G155gat), .ZN(new_n325));
  INV_X1    g124(.A(G162gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n330));
  INV_X1    g129(.A(G148gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G141gat), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G148gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT79), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(KEYINPUT79), .A3(G148gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n327), .A2(KEYINPUT80), .A3(new_n328), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n343));
  INV_X1    g142(.A(new_n328), .ZN(new_n344));
  NOR2_X1   g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n328), .A2(KEYINPUT2), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n341), .A2(new_n342), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n324), .B1(new_n350), .B2(KEYINPUT29), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT3), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n352), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n349), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G22gat), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n351), .A2(new_n354), .A3(G228gat), .A4(G233gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT83), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT31), .B(G50gat), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n363), .B(new_n364), .Z(new_n365));
  AOI21_X1  g164(.A(new_n317), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AND2_X1   g166(.A1(new_n357), .A2(new_n359), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n368), .A2(new_n358), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n362), .A2(new_n317), .A3(new_n365), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n367), .A2(new_n360), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n368), .B(new_n358), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n362), .A2(new_n317), .A3(new_n365), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n366), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n316), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT35), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n220), .A2(new_n222), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n346), .A2(new_n342), .A3(new_n347), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n336), .B1(new_n380), .B2(new_n341), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n352), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n220), .A2(new_n222), .A3(new_n381), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(G225gat), .A2(G233gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT81), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n225), .B1(new_n212), .B2(new_n219), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n383), .A2(new_n386), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n384), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n390), .A2(new_n381), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n388), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n392), .A2(new_n395), .A3(KEYINPUT5), .ZN(new_n396));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(KEYINPUT0), .ZN(new_n398));
  XNOR2_X1  g197(.A(G57gat), .B(G85gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  AOI22_X1  g199(.A1(new_n220), .A2(new_n222), .B1(new_n381), .B2(new_n352), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n388), .B1(new_n401), .B2(new_n379), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n384), .A2(new_n385), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT5), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n405), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n402), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n396), .A2(new_n400), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n400), .B1(new_n396), .B2(new_n407), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI211_X1 g211(.A(new_n409), .B(new_n400), .C1(new_n396), .C2(new_n407), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G8gat), .B(G36gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G64gat), .B(G92gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT77), .ZN(new_n419));
  INV_X1    g218(.A(new_n324), .ZN(new_n420));
  INV_X1    g219(.A(G226gat), .ZN(new_n421));
  INV_X1    g220(.A(G233gat), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI211_X1 g223(.A(new_n277), .B(new_n424), .C1(new_n259), .C2(new_n263), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(KEYINPUT29), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n293), .A2(new_n262), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n278), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n419), .B(new_n420), .C1(new_n425), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n278), .ZN(new_n431));
  OAI221_X1 g230(.A(new_n324), .B1(new_n431), .B2(new_n424), .C1(new_n298), .C2(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n264), .A2(new_n278), .ZN(new_n434));
  INV_X1    g233(.A(new_n431), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n434), .A2(new_n424), .B1(new_n435), .B2(new_n427), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n419), .B1(new_n436), .B2(new_n420), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n418), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n429), .B1(new_n298), .B2(new_n423), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT77), .B1(new_n439), .B2(new_n324), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n440), .A2(new_n432), .A3(new_n430), .A4(new_n417), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(KEYINPUT30), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n432), .A3(new_n430), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n417), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n414), .B1(new_n442), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n376), .A2(new_n377), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n289), .A2(new_n308), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n306), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n289), .A2(KEYINPUT74), .A3(new_n308), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n371), .A2(new_n374), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n313), .A2(new_n454), .A3(new_n447), .A4(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n456), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT86), .B1(new_n456), .B2(KEYINPUT35), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n448), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT36), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n313), .A2(new_n460), .A3(new_n315), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n306), .B1(new_n449), .B2(new_n450), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n453), .A2(new_n462), .B1(new_n311), .B2(new_n312), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n463), .B2(new_n460), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n418), .A2(KEYINPUT37), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n438), .A2(new_n466), .B1(KEYINPUT37), .B2(new_n443), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT38), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT37), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n444), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n418), .B1(new_n443), .B2(KEYINPUT37), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT85), .B(KEYINPUT38), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n411), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(new_n409), .A3(new_n408), .ZN(new_n475));
  INV_X1    g274(.A(new_n413), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n441), .ZN(new_n477));
  INV_X1    g276(.A(new_n472), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n434), .A2(new_n426), .B1(new_n435), .B2(new_n423), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n470), .B1(new_n479), .B2(new_n420), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n436), .A2(new_n324), .ZN(new_n481));
  AOI21_X1  g280(.A(KEYINPUT38), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n477), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n469), .A2(new_n473), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n383), .B(new_n406), .C1(new_n384), .C2(new_n385), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n388), .ZN(new_n486));
  OR3_X1    g285(.A1(new_n393), .A2(new_n394), .A3(new_n388), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT39), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT39), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(new_n489), .A3(new_n388), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n400), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n488), .A2(KEYINPUT40), .A3(new_n400), .A4(new_n490), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n493), .A2(new_n494), .A3(new_n474), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n495), .A2(new_n442), .A3(new_n446), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n496), .A2(new_n455), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n484), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n447), .A2(new_n455), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n459), .B1(new_n464), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G22gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(KEYINPUT88), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT16), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n504), .B1(new_n505), .B2(G1gat), .ZN(new_n506));
  INV_X1    g305(.A(G8gat), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT88), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n503), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(G1gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n507), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n507), .B1(new_n506), .B2(new_n511), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(KEYINPUT87), .B(G36gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  OR3_X1    g318(.A1(new_n518), .A2(G29gat), .A3(G36gat), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT15), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  XNOR2_X1  g323(.A(G43gat), .B(G50gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n527));
  OR3_X1    g326(.A1(new_n521), .A2(new_n522), .A3(new_n525), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n515), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT89), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  INV_X1    g332(.A(new_n515), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n526), .A2(new_n528), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n515), .B(new_n537), .C1(new_n529), .C2(new_n530), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n532), .A2(new_n533), .A3(new_n536), .A4(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n515), .B(new_n535), .Z(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(new_n533), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n539), .A2(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n536), .A2(new_n538), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n532), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G113gat), .B(G141gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G197gat), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT11), .B(G169gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n551), .B(KEYINPUT12), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n552), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n544), .A2(new_n554), .A3(new_n546), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(G57gat), .A2(G64gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(G57gat), .A2(G64gat), .ZN(new_n558));
  AND2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n557), .B(new_n558), .C1(new_n559), .C2(KEYINPUT9), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(KEYINPUT91), .B2(new_n559), .ZN(new_n561));
  NOR2_X1   g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n561), .B(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g364(.A1(G231gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n565), .B(new_n566), .Z(new_n567));
  XNOR2_X1  g366(.A(G127gat), .B(G155gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT20), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n569), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G183gat), .B(G211gat), .Z(new_n573));
  OR2_X1    g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n573), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n534), .B1(KEYINPUT21), .B2(new_n564), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n574), .A2(new_n579), .A3(new_n575), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT93), .B(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n589), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  AOI22_X1  g395(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n590), .A2(new_n592), .A3(new_n593), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT94), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n590), .A2(new_n593), .A3(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n591), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT95), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT95), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(new_n603), .A3(new_n591), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n599), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n564), .A2(KEYINPUT10), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n564), .A2(new_n598), .A3(new_n601), .ZN(new_n608));
  INV_X1    g407(.A(new_n564), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n587), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI211_X1 g414(.A(KEYINPUT10), .B(new_n608), .C1(new_n605), .C2(new_n609), .ZN(new_n616));
  OAI211_X1 g415(.A(KEYINPUT97), .B(new_n613), .C1(new_n616), .C2(new_n607), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n610), .A2(new_n613), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n586), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n586), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n613), .B1(new_n616), .B2(new_n607), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n605), .B1(new_n529), .B2(new_n530), .ZN(new_n626));
  NAND4_X1  g425(.A1(new_n535), .A2(new_n599), .A3(new_n602), .A4(new_n604), .ZN(new_n627));
  NAND3_X1  g426(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G134gat), .B(G162gat), .Z(new_n634));
  AOI21_X1  g433(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(KEYINPUT96), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n636), .B(KEYINPUT96), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n631), .A2(new_n632), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n583), .A2(new_n625), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n583), .A2(new_n625), .A3(KEYINPUT98), .A4(new_n642), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n502), .A2(new_n556), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(new_n414), .B(KEYINPUT99), .Z(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(new_n510), .ZN(G1324gat));
  NAND2_X1  g450(.A1(new_n442), .A2(new_n446), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(G8gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT16), .B(G8gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT42), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(KEYINPUT42), .B2(new_n656), .ZN(G1325gat));
  AOI21_X1  g457(.A(new_n460), .B1(new_n313), .B2(new_n454), .ZN(new_n659));
  AOI211_X1 g458(.A(KEYINPUT36), .B(new_n314), .C1(new_n311), .C2(new_n312), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT100), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n461), .B(new_n662), .C1(new_n463), .C2(new_n460), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n661), .A2(new_n663), .A3(KEYINPUT101), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT101), .B1(new_n661), .B2(new_n663), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(G15gat), .B1(new_n647), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n316), .A2(G15gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n647), .B2(new_n669), .ZN(G1326gat));
  NOR2_X1   g469(.A1(new_n647), .A2(new_n455), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT102), .ZN(new_n672));
  XNOR2_X1  g471(.A(KEYINPUT43), .B(G22gat), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(new_n583), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n625), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n642), .ZN(new_n677));
  INV_X1    g476(.A(new_n447), .ZN(new_n678));
  NOR4_X1   g477(.A1(new_n316), .A2(new_n678), .A3(new_n375), .A4(KEYINPUT35), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT86), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n456), .A2(KEYINPUT86), .A3(KEYINPUT35), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n679), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n501), .A2(new_n464), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n556), .B(new_n677), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(G29gat), .A3(new_n649), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT45), .Z(new_n688));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n642), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n691));
  AND3_X1   g490(.A1(new_n544), .A2(new_n554), .A3(new_n546), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n554), .B1(new_n544), .B2(new_n546), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n676), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n499), .B1(new_n484), .B2(new_n497), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n661), .A2(new_n663), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n642), .B1(new_n459), .B2(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n691), .B(new_n696), .C1(new_n699), .C2(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n649), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n688), .A2(new_n701), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n686), .A2(new_n652), .A3(new_n516), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n516), .B1(new_n700), .B2(new_n652), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  AND2_X1   g505(.A1(new_n661), .A2(new_n663), .ZN(new_n707));
  OAI21_X1  g506(.A(G43gat), .B1(new_n700), .B2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n686), .A2(G43gat), .A3(new_n316), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n700), .A2(new_n667), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n709), .B1(new_n713), .B2(G43gat), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n712), .B1(new_n714), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g514(.A1(new_n455), .A2(G50gat), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT48), .B1(new_n686), .B2(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n661), .A2(new_n663), .A3(new_n697), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n641), .B1(new_n684), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n689), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n721), .A2(new_n375), .A3(new_n691), .A4(new_n696), .ZN(new_n722));
  AOI211_X1 g521(.A(KEYINPUT105), .B(new_n718), .C1(new_n722), .C2(G50gat), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT105), .ZN(new_n724));
  OAI21_X1  g523(.A(G50gat), .B1(new_n700), .B2(new_n455), .ZN(new_n725));
  INV_X1    g524(.A(new_n718), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n728), .B(G50gat), .C1(new_n700), .C2(new_n455), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT48), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n686), .B2(new_n717), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n732), .B1(new_n722), .B2(G50gat), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n723), .A2(new_n727), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI221_X1 g535(.A(KEYINPUT106), .B1(new_n731), .B2(new_n733), .C1(new_n723), .C2(new_n727), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1331gat));
  NAND4_X1  g537(.A1(new_n583), .A2(new_n694), .A3(new_n642), .A4(new_n624), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n739), .B1(new_n459), .B2(new_n698), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n648), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT107), .B(G57gat), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1332gat));
  INV_X1    g542(.A(new_n652), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n746));
  AND2_X1   g545(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n745), .B2(new_n746), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT108), .ZN(G1333gat));
  NAND2_X1  g549(.A1(new_n740), .A2(new_n666), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n316), .A2(G71gat), .ZN(new_n752));
  AOI22_X1  g551(.A1(new_n751), .A2(G71gat), .B1(new_n740), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n740), .A2(new_n375), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n583), .A2(new_n556), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n721), .A2(new_n624), .A3(new_n691), .A4(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n649), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n699), .A2(new_n757), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT51), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n699), .A2(new_n762), .A3(new_n757), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n761), .A2(new_n763), .A3(new_n624), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n648), .A2(new_n595), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n759), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n758), .B2(new_n652), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n652), .A2(G92gat), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n761), .A2(new_n763), .A3(new_n624), .A4(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT109), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT109), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n767), .A2(new_n773), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n771), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n758), .B2(new_n667), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n316), .A2(G99gat), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n764), .B2(new_n780), .ZN(G1338gat));
  OR3_X1    g580(.A1(new_n764), .A2(G106gat), .A3(new_n455), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n758), .B2(new_n455), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n786), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1339gat));
  NOR2_X1   g587(.A1(new_n694), .A2(G113gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n463), .A2(new_n455), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n615), .A2(new_n792), .A3(new_n617), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n612), .A2(new_n614), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n622), .A3(KEYINPUT54), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n586), .A4(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n623), .B(new_n796), .C1(new_n692), .C2(new_n693), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n615), .A2(new_n792), .A3(new_n617), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT54), .B1(new_n612), .B2(new_n614), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n616), .A2(new_n613), .A3(new_n607), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n586), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n798), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT111), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n793), .A2(new_n586), .A3(new_n795), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n805), .A2(new_n806), .A3(new_n798), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n797), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n533), .B1(new_n545), .B2(new_n532), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n541), .A2(new_n543), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n551), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n555), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n620), .B2(new_n623), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n642), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n804), .A2(new_n807), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n796), .A2(new_n623), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n642), .A2(new_n812), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n583), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n643), .A2(new_n556), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n791), .B(new_n648), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n805), .A2(new_n806), .A3(new_n798), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n806), .B1(new_n805), .B2(new_n798), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n817), .B(new_n556), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n812), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n624), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n641), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n675), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(new_n821), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n649), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(KEYINPUT112), .A3(new_n791), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n824), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n652), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(KEYINPUT113), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n789), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n832), .A2(new_n833), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n376), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n744), .A3(new_n649), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n694), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(G1340gat));
  NOR2_X1   g645(.A1(new_n625), .A2(G120gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n847), .B1(new_n838), .B2(new_n839), .ZN(new_n848));
  OAI21_X1  g647(.A(G120gat), .B1(new_n844), .B2(new_n625), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n844), .B2(new_n675), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n583), .A2(new_n205), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n837), .B2(new_n852), .ZN(G1342gat));
  AOI21_X1  g652(.A(new_n206), .B1(new_n843), .B2(new_n641), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n641), .A2(new_n210), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT112), .B1(new_n834), .B2(new_n791), .ZN(new_n857));
  INV_X1    g656(.A(new_n797), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n813), .B1(new_n858), .B2(new_n815), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n819), .B1(new_n859), .B2(new_n641), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n821), .B1(new_n860), .B2(new_n675), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n861), .A2(new_n823), .A3(new_n790), .A4(new_n649), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n652), .B(new_n856), .C1(new_n857), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n854), .B1(new_n863), .B2(KEYINPUT56), .ZN(new_n864));
  AOI211_X1 g663(.A(new_n744), .B(new_n855), .C1(new_n824), .C2(new_n835), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT114), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n863), .A2(new_n868), .A3(KEYINPUT56), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n864), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g671(.A(KEYINPUT115), .B(new_n864), .C1(new_n867), .C2(new_n869), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1343gat));
  AND3_X1   g673(.A1(new_n707), .A2(new_n652), .A3(new_n648), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n455), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n803), .A2(KEYINPUT116), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n805), .A2(new_n880), .A3(new_n798), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n817), .A2(new_n879), .A3(new_n556), .A4(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n641), .B1(new_n882), .B2(new_n829), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n819), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n881), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n880), .B1(new_n805), .B2(new_n798), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n813), .B1(new_n888), .B2(new_n858), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n889), .A2(KEYINPUT117), .A3(new_n641), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n675), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n878), .B1(new_n891), .B2(new_n833), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n841), .B2(new_n375), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n556), .B(new_n875), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G141gat), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n375), .B1(new_n664), .B2(new_n665), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT118), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(KEYINPUT118), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n861), .A2(new_n744), .A3(new_n649), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n694), .A2(G141gat), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n897), .A2(new_n898), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n895), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT58), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n894), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT117), .B1(new_n889), .B2(new_n641), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n883), .A2(new_n884), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n819), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n821), .B1(new_n908), .B2(new_n675), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n861), .A2(new_n455), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n909), .A2(new_n878), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n911), .A2(KEYINPUT119), .A3(new_n556), .A4(new_n875), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n905), .A2(G141gat), .A3(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n901), .A2(new_n914), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n913), .A2(KEYINPUT120), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT120), .B1(new_n913), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n903), .B1(new_n916), .B2(new_n917), .ZN(G1344gat));
  AND2_X1   g717(.A1(new_n897), .A2(new_n899), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n919), .A2(new_n331), .A3(new_n624), .A4(new_n898), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n875), .A2(new_n624), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n675), .B1(new_n883), .B2(new_n831), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n645), .A2(new_n694), .A3(new_n646), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n455), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n925), .B2(KEYINPUT57), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n841), .A2(new_n877), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT121), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n923), .A2(new_n924), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n929), .B(new_n876), .C1(new_n930), .C2(new_n455), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n922), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n331), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n931), .A2(new_n927), .A3(new_n926), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n624), .A3(new_n875), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT122), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n921), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n911), .A2(new_n875), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(new_n625), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n940), .A2(KEYINPUT59), .A3(new_n331), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n920), .B1(new_n938), .B2(new_n941), .ZN(G1345gat));
  NAND4_X1  g741(.A1(new_n919), .A2(new_n325), .A3(new_n583), .A4(new_n898), .ZN(new_n943));
  OAI21_X1  g742(.A(G155gat), .B1(new_n939), .B2(new_n675), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  NAND4_X1  g744(.A1(new_n919), .A2(new_n326), .A3(new_n641), .A4(new_n898), .ZN(new_n946));
  OAI21_X1  g745(.A(G162gat), .B1(new_n939), .B2(new_n642), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(G1347gat));
  NOR2_X1   g747(.A1(new_n648), .A2(new_n652), .ZN(new_n949));
  AND3_X1   g748(.A1(new_n841), .A2(new_n791), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n556), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n841), .A2(new_n376), .A3(new_n949), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(new_n237), .A3(new_n694), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n953), .ZN(G1348gat));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n238), .A3(new_n624), .ZN(new_n955));
  OAI21_X1  g754(.A(G176gat), .B1(new_n952), .B2(new_n625), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1349gat));
  NAND3_X1  g756(.A1(new_n950), .A2(new_n265), .A3(new_n583), .ZN(new_n958));
  OAI21_X1  g757(.A(G183gat), .B1(new_n952), .B2(new_n675), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT60), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n960), .A2(KEYINPUT123), .A3(new_n961), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT124), .B1(new_n960), .B2(new_n961), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n960), .A2(KEYINPUT124), .A3(new_n961), .ZN(new_n967));
  OAI22_X1  g766(.A1(new_n964), .A2(new_n965), .B1(new_n966), .B2(new_n967), .ZN(G1350gat));
  OAI21_X1  g767(.A(G190gat), .B1(new_n952), .B2(new_n642), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT125), .Z(new_n970));
  OR2_X1    g769(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g770(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n950), .A2(new_n266), .A3(new_n641), .ZN(new_n974));
  OAI211_X1 g773(.A(new_n973), .B(new_n974), .C1(new_n970), .C2(new_n971), .ZN(G1351gat));
  NAND3_X1  g774(.A1(new_n667), .A2(new_n910), .A3(new_n949), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n556), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n935), .A2(new_n667), .A3(new_n949), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n556), .A2(G197gat), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  NOR3_X1   g781(.A1(new_n976), .A2(G204gat), .A3(new_n625), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  OAI21_X1  g783(.A(G204gat), .B1(new_n979), .B2(new_n625), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n977), .A2(new_n319), .A3(new_n583), .ZN(new_n987));
  NAND4_X1  g786(.A1(new_n935), .A2(new_n583), .A3(new_n667), .A4(new_n949), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(G211gat), .ZN(new_n989));
  NOR2_X1   g788(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n989), .A2(new_n990), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(G1354gat));
  OAI21_X1  g794(.A(G218gat), .B1(new_n979), .B2(new_n642), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n977), .A2(new_n320), .A3(new_n641), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1355gat));
endmodule


