//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1044,
    new_n1045;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT26), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT68), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT68), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT26), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AND2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n213), .B(KEYINPUT67), .C1(new_n214), .C2(KEYINPUT26), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n216), .B1(new_n217), .B2(new_n209), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n210), .A2(new_n215), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT27), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G183gat), .ZN(new_n223));
  INV_X1    g022(.A(G183gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT27), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT65), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT65), .B1(new_n224), .B2(KEYINPUT27), .ZN(new_n227));
  NOR2_X1   g026(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n226), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT28), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT27), .B(G183gat), .ZN(new_n232));
  INV_X1    g031(.A(G190gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n227), .B(new_n228), .C1(new_n232), .C2(KEYINPUT65), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n223), .A2(new_n225), .A3(new_n233), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(KEYINPUT28), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n221), .B1(new_n235), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT23), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n214), .B1(new_n213), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n233), .ZN(new_n245));
  NAND3_X1  g044(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n245), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  AOI211_X1 g048(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n242), .B(new_n244), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT25), .ZN(new_n252));
  INV_X1    g051(.A(new_n247), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n245), .A3(new_n246), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n243), .B1(G169gat), .B2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  AND4_X1   g055(.A1(KEYINPUT25), .A2(new_n242), .A3(new_n255), .A4(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n251), .A2(new_n252), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n203), .B1(new_n241), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n220), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n213), .B1(new_n214), .B2(KEYINPUT26), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n261), .A2(new_n216), .B1(new_n208), .B2(new_n209), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n262), .B2(new_n215), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n236), .A2(new_n237), .A3(new_n239), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n237), .B1(new_n236), .B2(new_n239), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n258), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT29), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n259), .B1(new_n268), .B2(new_n203), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270));
  OR2_X1    g069(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT22), .B1(new_n273), .B2(G218gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT72), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n280), .B1(new_n271), .B2(new_n272), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n275), .C1(new_n281), .C2(KEYINPUT22), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n274), .A2(new_n276), .ZN(new_n284));
  INV_X1    g083(.A(new_n278), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(new_n279), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n270), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n270), .A3(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n269), .A2(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n283), .A2(new_n270), .A3(new_n286), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n235), .A2(new_n240), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n258), .B1(new_n294), .B2(new_n263), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n202), .B1(new_n295), .B2(KEYINPUT29), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n296), .A3(new_n259), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G8gat), .B(G36gat), .ZN(new_n301));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n291), .A2(KEYINPUT74), .A3(new_n297), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n303), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n269), .A2(new_n290), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n296), .A2(new_n259), .B1(new_n288), .B2(new_n289), .ZN(new_n308));
  OAI211_X1 g107(.A(KEYINPUT30), .B(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT75), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n303), .B1(new_n291), .B2(new_n297), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(KEYINPUT30), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n305), .B1(new_n310), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n309), .A2(KEYINPUT75), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n312), .A2(new_n311), .A3(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n319), .A3(new_n305), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT77), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n321), .B1(new_n298), .B2(new_n306), .ZN(new_n322));
  AOI211_X1 g121(.A(KEYINPUT77), .B(new_n303), .C1(new_n291), .C2(new_n297), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n325));
  XNOR2_X1  g124(.A(G155gat), .B(G162gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G141gat), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT2), .ZN(new_n331));
  NAND2_X1  g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT2), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n326), .A2(new_n330), .A3(new_n337), .A4(new_n332), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  XOR2_X1   g140(.A(G127gat), .B(G134gat), .Z(new_n342));
  INV_X1    g141(.A(G120gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G113gat), .ZN(new_n344));
  INV_X1    g143(.A(G113gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G120gat), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n344), .A2(new_n346), .A3(KEYINPUT69), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT69), .B1(new_n344), .B2(new_n346), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n342), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n342), .A2(KEYINPUT1), .ZN(new_n352));
  OR3_X1    g151(.A1(new_n343), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT70), .B1(new_n343), .B2(G113gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n346), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  AOI22_X1  g156(.A1(new_n340), .A2(new_n341), .B1(new_n351), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n334), .A2(new_n338), .A3(KEYINPUT79), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(KEYINPUT3), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n351), .A2(new_n357), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n365), .A2(KEYINPUT4), .A3(new_n340), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n340), .A2(new_n351), .A3(new_n357), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n363), .A2(new_n364), .A3(new_n366), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n360), .A2(new_n361), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n371), .B2(new_n365), .ZN(new_n372));
  INV_X1    g171(.A(new_n364), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n376));
  XNOR2_X1  g175(.A(G1gat), .B(G29gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(G57gat), .B(G85gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n370), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n376), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n370), .B2(new_n374), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n381), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n386), .A2(new_n387), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n324), .A2(new_n325), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n315), .A2(new_n320), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n315), .A2(KEYINPUT81), .A3(new_n393), .A4(new_n320), .ZN(new_n397));
  INV_X1    g196(.A(G228gat), .ZN(new_n398));
  INV_X1    g197(.A(G233gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT29), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n283), .A2(new_n401), .A3(new_n286), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n340), .B1(new_n403), .B2(new_n341), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n293), .A2(new_n402), .B1(new_n404), .B2(KEYINPUT82), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n341), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n339), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT82), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n400), .B1(new_n405), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n293), .A2(new_n402), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n406), .A2(new_n360), .A3(new_n361), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n400), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(G22gat), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n404), .A2(KEYINPUT82), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n409), .A2(new_n411), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n400), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n413), .ZN(new_n421));
  XOR2_X1   g220(.A(G78gat), .B(G106gat), .Z(new_n422));
  XNOR2_X1  g221(.A(KEYINPUT31), .B(G50gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT83), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n415), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  OAI221_X1 g226(.A(G22gat), .B1(new_n425), .B2(new_n424), .C1(new_n410), .C2(new_n414), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n419), .A2(new_n420), .A3(new_n413), .A4(new_n424), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n295), .A2(new_n365), .ZN(new_n432));
  AND2_X1   g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n365), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n241), .B2(new_n258), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n437), .B(KEYINPUT34), .ZN(new_n438));
  XOR2_X1   g237(.A(G15gat), .B(G43gat), .Z(new_n439));
  XNOR2_X1  g238(.A(G71gat), .B(G99gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n434), .B1(new_n432), .B2(new_n436), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(KEYINPUT33), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT32), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n443), .A2(new_n445), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n438), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n443), .A2(new_n445), .ZN(new_n450));
  INV_X1    g249(.A(new_n438), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n446), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n431), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n396), .A2(new_n397), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n312), .A2(new_n321), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n325), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n460), .A2(new_n318), .A3(new_n305), .ZN(new_n461));
  INV_X1    g260(.A(new_n453), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT35), .ZN(new_n463));
  XOR2_X1   g262(.A(new_n381), .B(KEYINPUT84), .Z(new_n464));
  NAND3_X1  g263(.A1(new_n376), .A2(new_n384), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n388), .A3(new_n389), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n388), .A3(KEYINPUT87), .A4(new_n389), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n392), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(new_n431), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n319), .B1(new_n318), .B2(new_n305), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n390), .A2(new_n392), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n460), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT81), .B1(new_n477), .B2(new_n320), .ZN(new_n478));
  INV_X1    g277(.A(new_n397), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n431), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n453), .B(KEYINPUT36), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n318), .A3(new_n305), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n363), .A2(new_n366), .A3(new_n369), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n373), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT39), .B1(new_n372), .B2(new_n373), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n464), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT39), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n483), .A2(new_n488), .A3(new_n373), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT40), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n490), .A2(KEYINPUT85), .B1(new_n391), .B2(new_n464), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n381), .B(KEYINPUT84), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n483), .A2(new_n373), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n489), .B(new_n492), .C1(new_n493), .C2(new_n485), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT86), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT86), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n487), .A2(new_n497), .A3(KEYINPUT40), .A4(new_n489), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT85), .ZN(new_n500));
  INV_X1    g299(.A(new_n494), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n500), .B1(new_n501), .B2(KEYINPUT40), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n491), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  AND2_X1   g302(.A1(new_n427), .A2(new_n429), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n482), .A2(new_n503), .B1(new_n504), .B2(new_n428), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT37), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n306), .B1(new_n298), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n291), .A2(KEYINPUT37), .A3(new_n297), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT38), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n291), .A2(new_n297), .A3(KEYINPUT88), .A4(KEYINPUT37), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n507), .A2(new_n510), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n324), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n300), .A2(KEYINPUT37), .A3(new_n304), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n511), .B1(new_n515), .B2(new_n507), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n470), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n481), .B1(new_n505), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n456), .A2(new_n473), .B1(new_n480), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G50gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(G43gat), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n524), .B1(G43gat), .B2(new_n521), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(G29gat), .ZN(new_n528));
  INV_X1    g327(.A(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT90), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n534), .A2(new_n535), .B1(new_n528), .B2(new_n529), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n526), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(KEYINPUT91), .A2(G43gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(KEYINPUT91), .A2(G43gat), .ZN(new_n539));
  AOI21_X1  g338(.A(G50gat), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n524), .B1(new_n540), .B2(new_n522), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT92), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n534), .A2(KEYINPUT92), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n523), .A2(new_n525), .B1(G29gat), .B2(G36gat), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n541), .A2(new_n543), .A3(new_n544), .A4(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n537), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n549), .B1(new_n537), .B2(new_n546), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT8), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(G85gat), .B2(G92gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT95), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n555), .B1(new_n556), .B2(KEYINPUT7), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n555), .A3(KEYINPUT7), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT96), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n561), .B1(new_n556), .B2(KEYINPUT7), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n563), .A2(KEYINPUT96), .A3(G85gat), .A4(G92gat), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n560), .A2(KEYINPUT97), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n556), .A2(new_n555), .A3(KEYINPUT7), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(new_n557), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n562), .A2(new_n564), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n566), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n554), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(G99gat), .B(G106gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT98), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AOI211_X1 g374(.A(new_n554), .B(new_n573), .C1(new_n565), .C2(new_n570), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n551), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT99), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n537), .A2(new_n546), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n565), .A2(new_n570), .ZN(new_n585));
  INV_X1    g384(.A(new_n554), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n573), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n574), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n547), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n582), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n578), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT100), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n578), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n590), .A2(KEYINPUT99), .A3(new_n582), .ZN(new_n597));
  AOI21_X1  g396(.A(KEYINPUT99), .B1(new_n590), .B2(new_n582), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT100), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(new_n593), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n594), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n604), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n595), .A2(new_n601), .A3(new_n606), .A4(new_n602), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G134gat), .B(G162gat), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n615));
  XOR2_X1   g414(.A(G57gat), .B(G64gat), .Z(new_n616));
  INV_X1    g415(.A(KEYINPUT9), .ZN(new_n617));
  INV_X1    g416(.A(G71gat), .ZN(new_n618));
  INV_X1    g417(.A(G78gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G71gat), .B(G78gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n616), .A2(new_n622), .A3(new_n620), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n624), .B2(new_n626), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(G231gat), .B(G233gat), .C1(new_n629), .C2(KEYINPUT21), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT21), .ZN(new_n632));
  INV_X1    g431(.A(G231gat), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n631), .B(new_n632), .C1(new_n633), .C2(new_n399), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(new_n637), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n615), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  INV_X1    g441(.A(new_n615), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n642), .A2(new_n638), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G15gat), .B(G22gat), .ZN(new_n645));
  INV_X1    g444(.A(G1gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(KEYINPUT16), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G8gat), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n650), .B1(new_n629), .B2(KEYINPUT21), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n641), .A2(new_n644), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n652), .B1(new_n641), .B2(new_n644), .ZN(new_n655));
  XOR2_X1   g454(.A(G183gat), .B(G211gat), .Z(new_n656));
  OR3_X1    g455(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n654), .B2(new_n655), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n614), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n649), .B1(new_n548), .B2(new_n550), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n650), .A2(new_n547), .ZN(new_n662));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n661), .A2(KEYINPUT18), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(KEYINPUT13), .Z(new_n665));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n547), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n580), .A2(new_n649), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT93), .ZN(new_n673));
  XOR2_X1   g472(.A(G113gat), .B(G141gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT11), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT89), .ZN(new_n676));
  XOR2_X1   g475(.A(G169gat), .B(G197gat), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT89), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n675), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT12), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n679), .B2(new_n682), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n669), .B(new_n672), .C1(new_n673), .C2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n664), .A2(new_n673), .A3(new_n668), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n684), .A2(new_n685), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n670), .A2(new_n671), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n664), .A2(new_n668), .ZN(new_n691));
  OAI211_X1 g490(.A(new_n688), .B(new_n689), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n687), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n624), .A2(new_n626), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n588), .A2(new_n694), .A3(new_n589), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n631), .B1(new_n575), .B2(new_n576), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT10), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n577), .A2(KEYINPUT10), .A3(new_n629), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(G230gat), .A2(G233gat), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT101), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n703));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n703), .B(new_n704), .C1(new_n698), .C2(new_n699), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n701), .B1(new_n695), .B2(new_n696), .ZN(new_n707));
  XNOR2_X1  g506(.A(G120gat), .B(G148gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(G176gat), .B(G204gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n704), .B1(new_n698), .B2(new_n699), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n710), .B1(new_n713), .B2(new_n707), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR4_X1   g514(.A1(new_n520), .A2(new_n660), .A3(new_n693), .A4(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT102), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n475), .B(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g520(.A1(new_n716), .A2(new_n482), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT16), .B(G8gat), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(KEYINPUT42), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT42), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n722), .B2(G8gat), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n726), .B1(new_n725), .B2(new_n728), .ZN(G1325gat));
  INV_X1    g528(.A(G15gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n716), .A2(new_n730), .A3(new_n462), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n481), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(new_n730), .ZN(G1326gat));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n431), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT103), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT43), .B(G22gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1327gat));
  NOR2_X1   g537(.A1(new_n520), .A2(new_n614), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n659), .A2(new_n693), .A3(new_n715), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(G29gat), .A3(new_n718), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(KEYINPUT45), .Z(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n520), .B2(new_n614), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n472), .B1(new_n455), .B2(KEYINPUT35), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT36), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n748), .B1(new_n449), .B2(new_n452), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n491), .A2(new_n499), .A3(new_n502), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n430), .B1(new_n461), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n752), .B2(new_n517), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n396), .A2(new_n397), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n753), .B1(new_n754), .B2(new_n431), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT44), .B(new_n613), .C1(new_n746), .C2(new_n755), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n745), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n719), .A3(new_n740), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(KEYINPUT104), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(KEYINPUT104), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G29gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n743), .B1(new_n759), .B2(new_n761), .ZN(G1328gat));
  NOR3_X1   g561(.A1(new_n741), .A2(G36gat), .A3(new_n461), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT46), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n757), .A2(new_n482), .A3(new_n740), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n529), .B2(new_n765), .ZN(G1329gat));
  NAND4_X1  g565(.A1(new_n745), .A2(new_n481), .A3(new_n740), .A4(new_n756), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n538), .A2(new_n539), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n453), .A2(new_n768), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n769), .B(KEYINPUT47), .C1(new_n741), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(KEYINPUT106), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n767), .A2(new_n774), .A3(new_n768), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(new_n741), .B2(new_n771), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n739), .A2(KEYINPUT107), .A3(new_n740), .A4(new_n770), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n773), .A2(new_n775), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(G1330gat));
  NAND3_X1  g580(.A1(new_n757), .A2(new_n431), .A3(new_n740), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G50gat), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT108), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n739), .A2(new_n521), .A3(new_n431), .A4(new_n740), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n783), .B(new_n785), .C1(KEYINPUT108), .C2(KEYINPUT48), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1331gat));
  NAND2_X1  g589(.A1(new_n687), .A2(new_n692), .ZN(new_n791));
  INV_X1    g590(.A(new_n715), .ZN(new_n792));
  NOR4_X1   g591(.A1(new_n520), .A2(new_n660), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(new_n719), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g594(.A(new_n482), .B(KEYINPUT109), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n799));
  AND2_X1   g598(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n800));
  NOR3_X1   g599(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n799), .B2(new_n798), .ZN(G1333gat));
  NAND3_X1  g601(.A1(new_n793), .A2(new_n618), .A3(new_n462), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n793), .A2(new_n481), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n804), .B1(G71gat), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g606(.A1(new_n793), .A2(new_n431), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g608(.A1(new_n718), .A2(G85gat), .A3(new_n792), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n520), .B2(new_n614), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n659), .A2(new_n791), .ZN(new_n813));
  OAI211_X1 g612(.A(KEYINPUT110), .B(new_n613), .C1(new_n746), .C2(new_n755), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n810), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n659), .A2(new_n791), .A3(new_n792), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n757), .A2(new_n719), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G85gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(G1336gat));
  INV_X1    g623(.A(KEYINPUT112), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n456), .A2(new_n473), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n480), .A2(new_n519), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT110), .B1(new_n828), .B2(new_n613), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n813), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n825), .B(KEYINPUT51), .C1(new_n829), .C2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n815), .B2(new_n825), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n796), .A2(G92gat), .A3(new_n792), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n745), .A2(new_n482), .A3(new_n756), .A4(new_n821), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(G92gat), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(KEYINPUT52), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n834), .B1(new_n818), .B2(new_n819), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n757), .A2(new_n797), .A3(new_n821), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n845), .B2(G92gat), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n843), .A2(new_n847), .ZN(G1337gat));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n757), .A2(new_n481), .A3(new_n821), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G99gat), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n792), .A2(G99gat), .A3(new_n453), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n815), .A2(new_n816), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(new_n817), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n849), .B1(new_n852), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n853), .B1(new_n818), .B2(new_n819), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(KEYINPUT113), .A3(new_n851), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(G1338gat));
  NOR3_X1   g659(.A1(new_n792), .A2(new_n430), .A3(G106gat), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n832), .A2(new_n833), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n745), .A2(new_n431), .A3(new_n756), .A4(new_n821), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(G106gat), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT53), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n861), .B1(new_n818), .B2(new_n819), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n865), .A2(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n866), .A2(new_n869), .ZN(G1339gat));
  AND2_X1   g669(.A1(new_n657), .A2(new_n658), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n871), .A2(new_n613), .A3(new_n791), .A4(new_n715), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n700), .A2(new_n701), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n710), .B1(new_n873), .B2(KEYINPUT54), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n698), .A2(new_n699), .A3(new_n704), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT54), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n874), .B1(new_n706), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n791), .B1(new_n877), .B2(KEYINPUT55), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n873), .A2(new_n703), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n713), .A2(KEYINPUT101), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n879), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n874), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT55), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n712), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n669), .A2(new_n686), .A3(new_n672), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n663), .B1(new_n661), .B2(new_n662), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n666), .A2(new_n667), .A3(new_n665), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n679), .B(new_n682), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  OAI22_X1  g688(.A1(new_n878), .A2(new_n884), .B1(new_n792), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n612), .A3(new_n610), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n877), .A2(KEYINPUT55), .B1(new_n706), .B2(new_n711), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n881), .A2(new_n882), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT55), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n613), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n659), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  OR2_X1    g697(.A1(new_n872), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n719), .A3(new_n796), .ZN(new_n900));
  INV_X1    g699(.A(new_n454), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n791), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G113gat), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n904), .A2(KEYINPUT114), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(KEYINPUT114), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n905), .A2(new_n906), .B1(G113gat), .B2(new_n903), .ZN(G1340gat));
  NAND2_X1  g706(.A1(new_n902), .A2(new_n715), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g708(.A1(new_n902), .A2(new_n659), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g710(.A1(new_n902), .A2(new_n613), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G134gat), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n899), .A2(new_n461), .A3(new_n613), .A4(new_n719), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n901), .A2(G134gat), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n918), .B1(new_n917), .B2(new_n914), .ZN(new_n919));
  NOR4_X1   g718(.A1(new_n915), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n916), .ZN(new_n920));
  OAI221_X1 g719(.A(new_n913), .B1(new_n914), .B2(new_n917), .C1(new_n919), .C2(new_n920), .ZN(G1343gat));
  NAND2_X1  g720(.A1(new_n750), .A2(new_n431), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n900), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n328), .A3(new_n791), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT58), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n796), .A2(new_n750), .A3(new_n719), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n899), .A2(new_n431), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT57), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT57), .B(new_n431), .C1(new_n872), .C2(new_n898), .ZN(new_n930));
  AOI211_X1 g729(.A(new_n693), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  OAI221_X1 g730(.A(new_n924), .B1(KEYINPUT116), .B2(new_n925), .C1(new_n931), .C2(new_n328), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n925), .B1(new_n924), .B2(KEYINPUT116), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n328), .B1(new_n934), .B2(new_n791), .ZN(new_n935));
  INV_X1    g734(.A(new_n924), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n937), .ZN(G1344gat));
  NAND3_X1  g737(.A1(new_n923), .A2(new_n329), .A3(new_n715), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT59), .B(new_n329), .C1(new_n934), .C2(new_n715), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT59), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n891), .A2(new_n897), .A3(KEYINPUT117), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT117), .B1(new_n891), .B2(new_n897), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n871), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n872), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n430), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n930), .B1(new_n946), .B2(KEYINPUT57), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n926), .A2(new_n792), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n941), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n939), .B1(new_n940), .B2(new_n950), .ZN(G1345gat));
  NAND3_X1  g750(.A1(new_n923), .A2(new_n335), .A3(new_n659), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n934), .A2(new_n659), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n952), .B1(new_n953), .B2(new_n335), .ZN(G1346gat));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n336), .B1(new_n934), .B2(new_n613), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n915), .A2(G162gat), .A3(new_n922), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(new_n957), .ZN(new_n959));
  AOI211_X1 g758(.A(new_n614), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n959), .B(KEYINPUT118), .C1(new_n960), .C2(new_n336), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(G1347gat));
  NAND3_X1  g761(.A1(new_n718), .A2(new_n462), .A3(new_n482), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AND2_X1   g763(.A1(new_n964), .A2(KEYINPUT120), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n964), .A2(KEYINPUT120), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n965), .A2(new_n966), .A3(new_n431), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n899), .A2(G169gat), .A3(new_n791), .A4(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n899), .A2(new_n718), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n901), .A2(new_n796), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT119), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n970), .A2(new_n791), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(new_n969), .B1(new_n973), .B2(new_n211), .ZN(G1348gat));
  NAND2_X1  g773(.A1(new_n970), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n212), .B1(new_n975), .B2(new_n792), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n977));
  OR2_X1    g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n899), .A2(G176gat), .A3(new_n715), .A4(new_n967), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n980), .B(KEYINPUT122), .Z(new_n981));
  AND3_X1   g780(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(G1349gat));
  INV_X1    g781(.A(KEYINPUT123), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n659), .A2(new_n232), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n899), .A2(new_n659), .A3(new_n967), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(G183gat), .ZN(new_n987));
  INV_X1    g786(.A(new_n984), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n970), .A2(KEYINPUT123), .A3(new_n972), .A4(new_n988), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n985), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT60), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n985), .A2(new_n987), .A3(new_n992), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n991), .A2(new_n993), .ZN(G1350gat));
  NAND3_X1  g793(.A1(new_n899), .A2(new_n613), .A3(new_n967), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n995), .A2(new_n996), .A3(G190gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n996), .B1(new_n995), .B2(G190gat), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n613), .A2(new_n233), .ZN(new_n999));
  OAI22_X1  g798(.A1(new_n997), .A2(new_n998), .B1(new_n975), .B2(new_n999), .ZN(G1351gat));
  INV_X1    g799(.A(new_n930), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT117), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n889), .B1(new_n712), .B2(new_n714), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n693), .B1(new_n893), .B2(new_n894), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1003), .B1(new_n892), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n613), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n892), .A2(new_n895), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n1007), .B1(new_n612), .B2(new_n610), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1002), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n891), .A2(new_n897), .A3(KEYINPUT117), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n659), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n431), .B1(new_n1011), .B2(new_n872), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n1001), .B1(new_n1012), .B2(new_n928), .ZN(new_n1013));
  NOR3_X1   g812(.A1(new_n481), .A2(new_n719), .A3(new_n461), .ZN(new_n1014));
  XNOR2_X1  g813(.A(new_n1014), .B(KEYINPUT125), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n791), .A2(G197gat), .ZN(new_n1016));
  NOR3_X1   g815(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g816(.A1(new_n922), .A2(new_n796), .ZN(new_n1018));
  OAI211_X1 g817(.A(new_n718), .B(new_n1018), .C1(new_n872), .C2(new_n898), .ZN(new_n1019));
  XNOR2_X1  g818(.A(new_n1019), .B(KEYINPUT124), .ZN(new_n1020));
  AOI21_X1  g819(.A(G197gat), .B1(new_n1020), .B2(new_n791), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1022));
  OR3_X1    g821(.A1(new_n1017), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1022), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1023), .A2(new_n1024), .ZN(G1352gat));
  OR2_X1    g824(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1026));
  OAI21_X1  g825(.A(G204gat), .B1(new_n1026), .B2(new_n792), .ZN(new_n1027));
  NOR3_X1   g826(.A1(new_n1019), .A2(G204gat), .A3(new_n792), .ZN(new_n1028));
  XNOR2_X1  g827(.A(new_n1028), .B(KEYINPUT62), .ZN(new_n1029));
  NAND2_X1  g828(.A1(new_n1027), .A2(new_n1029), .ZN(G1353gat));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n659), .ZN(new_n1031));
  OAI211_X1 g830(.A(KEYINPUT63), .B(G211gat), .C1(new_n1013), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1032), .A2(KEYINPUT127), .ZN(new_n1033));
  INV_X1    g832(.A(new_n1031), .ZN(new_n1034));
  NAND2_X1  g833(.A1(new_n947), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1036));
  NAND4_X1  g835(.A1(new_n1035), .A2(new_n1036), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1037));
  OAI21_X1  g836(.A(G211gat), .B1(new_n1013), .B2(new_n1031), .ZN(new_n1038));
  INV_X1    g837(.A(KEYINPUT63), .ZN(new_n1039));
  NAND2_X1  g838(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g839(.A1(new_n1033), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NAND4_X1  g840(.A1(new_n1020), .A2(new_n271), .A3(new_n272), .A4(new_n659), .ZN(new_n1042));
  NAND2_X1  g841(.A1(new_n1041), .A2(new_n1042), .ZN(G1354gat));
  OAI21_X1  g842(.A(G218gat), .B1(new_n1026), .B2(new_n614), .ZN(new_n1044));
  NAND3_X1  g843(.A1(new_n1020), .A2(new_n280), .A3(new_n613), .ZN(new_n1045));
  NAND2_X1  g844(.A1(new_n1044), .A2(new_n1045), .ZN(G1355gat));
endmodule


