//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(G122), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT92), .B1(new_n187), .B2(G116), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT92), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(new_n190), .A3(G122), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT14), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n187), .A2(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n192), .A2(KEYINPUT14), .ZN(new_n196));
  OAI21_X1  g010(.A(G107), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n198), .A3(new_n194), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT93), .B1(new_n200), .B2(G143), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT93), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G128), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(G143), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G134), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n209), .A3(new_n206), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n197), .A2(new_n199), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n192), .A2(new_n194), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n199), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT13), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n205), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n201), .A2(new_n204), .A3(KEYINPUT13), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n217), .A2(new_n218), .A3(new_n206), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n215), .B(new_n210), .C1(new_n219), .C2(new_n209), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT9), .B(G234), .ZN(new_n222));
  INV_X1    g036(.A(G217), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n222), .A2(new_n223), .A3(G953), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n221), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n212), .A2(new_n220), .A3(new_n224), .ZN(new_n227));
  AOI21_X1  g041(.A(G902), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G478), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT15), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n228), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(G113), .B(G122), .ZN(new_n233));
  INV_X1    g047(.A(G104), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G140), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G125), .ZN(new_n237));
  INV_X1    g051(.A(G125), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G140), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(G146), .ZN(new_n241));
  NOR2_X1   g055(.A1(G237), .A2(G953), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(G143), .A3(G214), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(G143), .B1(new_n242), .B2(G214), .ZN(new_n245));
  OAI211_X1 g059(.A(KEYINPUT18), .B(G131), .C1(new_n244), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT18), .A2(G131), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n243), .A3(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n241), .A2(new_n246), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n244), .B2(new_n245), .ZN(new_n251));
  INV_X1    g065(.A(G131), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n252), .A3(new_n243), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT17), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT16), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n236), .A3(G125), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n240), .B2(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(G146), .B(new_n257), .C1(new_n240), .C2(new_n256), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT17), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n260), .B(new_n261), .C1(new_n262), .C2(new_n251), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n235), .B(new_n250), .C1(new_n255), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n250), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n261), .B(KEYINPUT72), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT19), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n240), .B(new_n267), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n268), .A2(new_n259), .B1(new_n251), .B2(new_n253), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n265), .B1(new_n266), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n264), .B1(new_n270), .B2(new_n235), .ZN(new_n271));
  NOR2_X1   g085(.A1(G475), .A2(G902), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(KEYINPUT20), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT20), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n271), .B2(new_n272), .ZN(new_n276));
  INV_X1    g090(.A(G475), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n250), .B1(new_n255), .B2(new_n263), .ZN(new_n278));
  INV_X1    g092(.A(new_n235), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n280), .B2(new_n264), .ZN(new_n281));
  OAI22_X1  g095(.A1(new_n274), .A2(new_n276), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n232), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(G952), .ZN(new_n285));
  NAND2_X1  g099(.A1(G234), .A2(G237), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(G902), .A3(G953), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT21), .B(G898), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT91), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n203), .A2(G146), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT64), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n300), .B1(new_n259), .B2(G143), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT0), .A2(G128), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT0), .A2(G128), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n259), .A2(G143), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n203), .A2(G146), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n303), .A2(new_n305), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(KEYINPUT86), .B1(new_n311), .B2(new_n238), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n303), .A2(new_n305), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n307), .A2(new_n310), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT86), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G125), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n203), .A2(KEYINPUT64), .A3(G146), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT64), .B1(new_n203), .B2(G146), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n308), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT1), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(G143), .B2(new_n259), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n310), .B1(new_n323), .B2(new_n200), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n325), .A2(new_n326), .A3(G125), .ZN(new_n327));
  OAI21_X1  g141(.A(G128), .B1(new_n299), .B2(new_n322), .ZN(new_n328));
  AOI22_X1  g142(.A1(new_n303), .A2(new_n318), .B1(new_n328), .B2(new_n310), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT87), .B1(new_n329), .B2(new_n238), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n312), .B(new_n317), .C1(new_n327), .C2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G224), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G953), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n190), .A2(G119), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT5), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT83), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT5), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT84), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n336), .A2(new_n338), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G113), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(new_n336), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G119), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G116), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n190), .A2(G119), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT66), .ZN(new_n351));
  XNOR2_X1  g165(.A(G116), .B(G119), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n346), .B1(new_n355), .B2(new_n344), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT2), .B(G113), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n198), .A2(G104), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n234), .A2(G107), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n360), .B2(KEYINPUT76), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(new_n198), .A3(KEYINPUT3), .A4(G104), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n359), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n362), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n356), .A2(new_n358), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G110), .B(G122), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n351), .A2(new_n354), .A3(new_n357), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n234), .A2(G107), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT3), .B1(new_n374), .B2(new_n365), .ZN(new_n375));
  INV_X1    g189(.A(new_n366), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n361), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n373), .A2(new_n358), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n198), .A2(G104), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n364), .B2(new_n366), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(KEYINPUT4), .C1(new_n382), .C2(new_n359), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n379), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT82), .B1(new_n379), .B2(new_n383), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n371), .B(new_n372), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT6), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n371), .B1(new_n384), .B2(new_n385), .ZN(new_n388));
  XOR2_X1   g202(.A(new_n372), .B(KEYINPUT85), .Z(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n335), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n327), .A2(new_n330), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n317), .A2(new_n312), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  OAI22_X1  g210(.A1(new_n394), .A2(new_n395), .B1(new_n396), .B2(new_n333), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT7), .B1(new_n332), .B2(G953), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n331), .B(new_n398), .C1(new_n396), .C2(new_n333), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n372), .B(KEYINPUT8), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n370), .A2(new_n358), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n346), .A2(KEYINPUT89), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT88), .B1(new_n350), .B2(new_n337), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n352), .A2(new_n406), .A3(KEYINPUT5), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n346), .B2(KEYINPUT89), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n403), .B1(new_n404), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n370), .B1(new_n356), .B2(new_n358), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n402), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n400), .A2(new_n386), .A3(new_n401), .A4(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G902), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n298), .B1(new_n393), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n413), .A2(new_n414), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n386), .A2(KEYINPUT6), .B1(new_n388), .B2(new_n389), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n388), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n334), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n420), .A3(new_n297), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(G214), .B1(G237), .B2(G902), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n423), .B(KEYINPUT80), .Z(new_n424));
  XOR2_X1   g238(.A(new_n424), .B(KEYINPUT81), .Z(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n296), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  AOI211_X1 g241(.A(KEYINPUT91), .B(new_n425), .C1(new_n416), .C2(new_n421), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n295), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G221), .B1(new_n222), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT78), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n323), .A2(new_n200), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n321), .B1(new_n303), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n370), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n377), .A2(new_n378), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n359), .B1(new_n367), .B2(new_n361), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n311), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G137), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT11), .A3(G134), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n209), .A2(G137), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n209), .B2(G137), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n444), .A2(KEYINPUT65), .A3(new_n252), .A4(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n446), .A2(new_n442), .A3(new_n252), .A4(new_n443), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT65), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n446), .A2(new_n442), .A3(new_n443), .ZN(new_n451));
  AOI22_X1  g265(.A1(new_n447), .A2(new_n450), .B1(G131), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n370), .A2(KEYINPUT10), .A3(new_n325), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n436), .A2(new_n440), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G140), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n284), .A2(G227), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n455), .B(new_n456), .Z(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n436), .A2(new_n440), .A3(new_n453), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n451), .A2(G131), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n448), .A2(new_n449), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n448), .A2(new_n449), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT77), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n459), .A2(KEYINPUT77), .A3(new_n463), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XOR2_X1   g282(.A(new_n457), .B(KEYINPUT75), .Z(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n368), .B1(new_n364), .B2(new_n366), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n321), .B(new_n324), .C1(new_n471), .C2(new_n362), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n434), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n463), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(KEYINPUT12), .A3(new_n463), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n470), .B1(new_n478), .B2(new_n454), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n431), .B1(new_n468), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n458), .ZN(new_n481));
  INV_X1    g295(.A(new_n467), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT77), .B1(new_n459), .B2(new_n463), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n477), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT12), .B1(new_n473), .B2(new_n463), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n454), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n469), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n484), .A2(KEYINPUT78), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n489), .A3(new_n414), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(G469), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n458), .B1(new_n477), .B2(new_n476), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n454), .B1(new_n482), .B2(new_n483), .ZN(new_n494));
  INV_X1    g308(.A(new_n457), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n496), .A2(G469), .A3(G902), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n491), .B1(new_n490), .B2(G469), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n430), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n429), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n373), .A2(new_n358), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n463), .B2(new_n311), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n447), .A2(new_n450), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n441), .A2(G134), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n252), .B1(new_n506), .B2(new_n443), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n321), .B2(new_n324), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT67), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT67), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n504), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n242), .A2(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n513), .A2(KEYINPUT68), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT68), .B1(new_n513), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n373), .A2(new_n358), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n463), .A2(new_n311), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n510), .A2(new_n522), .A3(new_n512), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT30), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n525), .A3(new_n509), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n521), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n502), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT68), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n521), .B1(new_n452), .B2(new_n315), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n505), .A2(new_n511), .A3(new_n508), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n511), .B1(new_n505), .B2(new_n508), .ZN(new_n532));
  NOR3_X1   g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n517), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n513), .A2(KEYINPUT68), .A3(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n531), .A2(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n525), .B1(new_n538), .B2(new_n522), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n522), .A2(new_n525), .A3(new_n509), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n503), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n522), .A2(new_n509), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n503), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n504), .A2(new_n510), .A3(KEYINPUT28), .A4(new_n512), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n509), .B(new_n521), .C1(new_n452), .C2(new_n315), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n528), .A2(new_n542), .B1(new_n534), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G472), .A2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n550), .A2(KEYINPUT32), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT32), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n549), .A2(new_n534), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n541), .ZN(new_n556));
  AOI21_X1  g370(.A(KEYINPUT31), .B1(new_n537), .B2(new_n541), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n554), .B1(new_n558), .B2(new_n551), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT69), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n534), .A2(new_n561), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n503), .A2(new_n523), .B1(new_n538), .B2(new_n504), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n548), .B(new_n562), .C1(new_n563), .C2(new_n547), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n517), .B1(new_n541), .B2(new_n513), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n544), .A2(new_n545), .A3(new_n548), .A4(new_n517), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n561), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n414), .B(new_n564), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n560), .B1(new_n568), .B2(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n540), .B1(KEYINPUT30), .B2(new_n523), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n513), .B1(new_n570), .B2(new_n521), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n571), .B2(new_n534), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n414), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n560), .B(G472), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  OAI22_X1  g389(.A1(new_n553), .A2(new_n559), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT70), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n568), .A2(G472), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT69), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n574), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT32), .B1(new_n550), .B2(new_n552), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n558), .A2(new_n554), .A3(new_n551), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT70), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT25), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n284), .A2(G221), .A3(G234), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(KEYINPUT73), .ZN(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT22), .B(G137), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n588), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT74), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n240), .A2(G146), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n347), .A2(G128), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n347), .A2(G128), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(KEYINPUT23), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n600), .A2(G110), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n200), .A2(G119), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT24), .B(G110), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n596), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n266), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(G110), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT71), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n260), .A2(new_n261), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n603), .B2(new_n604), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n607), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n595), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n607), .B(new_n593), .C1(new_n609), .C2(new_n611), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n586), .B1(new_n615), .B2(G902), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n613), .A2(KEYINPUT25), .A3(new_n414), .A4(new_n614), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n223), .B1(G234), .B2(new_n414), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n615), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n619), .A2(G902), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n501), .A2(new_n578), .A3(new_n585), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  OAI21_X1  g441(.A(G472), .B1(new_n550), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n558), .A2(new_n551), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n500), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n282), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n225), .B2(KEYINPUT94), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n226), .A2(new_n227), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n634), .B1(new_n226), .B2(new_n227), .ZN(new_n636));
  OAI21_X1  g450(.A(G478), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n229), .A2(new_n414), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n228), .B2(new_n229), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OR3_X1    g454(.A1(new_n632), .A2(KEYINPUT95), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n640), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n282), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT95), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n424), .B1(new_n416), .B2(new_n421), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n645), .A2(new_n293), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n631), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  INV_X1    g464(.A(new_n646), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n281), .A2(new_n277), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT96), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n274), .A2(new_n276), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR4_X1   g470(.A1(new_n651), .A2(new_n292), .A3(new_n231), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT35), .B(G107), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  NOR3_X1   g474(.A1(new_n393), .A2(new_n298), .A3(new_n415), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n297), .B1(new_n417), .B2(new_n420), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n426), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT91), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n422), .A2(new_n296), .A3(new_n426), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n294), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n430), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n492), .A2(new_n497), .ZN(new_n668));
  INV_X1    g482(.A(new_n499), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n628), .A2(new_n629), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(new_n612), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n618), .A2(new_n619), .B1(new_n622), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n670), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  XNOR2_X1  g492(.A(KEYINPUT97), .B(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n288), .B1(new_n679), .B2(new_n290), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n653), .A2(new_n655), .A3(new_n232), .A4(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n651), .A2(new_n674), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n578), .A2(new_n585), .A3(new_n670), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G128), .ZN(G30));
  XOR2_X1   g499(.A(new_n680), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n670), .A2(new_n686), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n520), .A2(new_n527), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n523), .A2(new_n503), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n513), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n690), .B1(new_n534), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(G472), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n584), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n422), .B(KEYINPUT38), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n632), .A2(new_n424), .A3(new_n231), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n674), .A2(new_n695), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n688), .A2(new_n689), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G143), .ZN(G45));
  NAND3_X1  g514(.A1(new_n642), .A2(new_n282), .A3(new_n681), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n674), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n646), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n578), .A2(new_n585), .A3(new_n670), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT98), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n500), .A2(new_n704), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT98), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n708), .A2(new_n709), .A3(new_n578), .A4(new_n585), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT99), .B(G146), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G48));
  OAI21_X1  g527(.A(G469), .B1(new_n496), .B2(G902), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n497), .A2(new_n430), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n624), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n647), .A2(new_n578), .A3(new_n585), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND4_X1  g533(.A1(new_n578), .A2(new_n657), .A3(new_n585), .A4(new_n716), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G116), .ZN(G18));
  NOR2_X1   g535(.A1(new_n651), .A2(new_n715), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n294), .A2(new_n674), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n578), .A2(new_n585), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G119), .ZN(G21));
  NAND2_X1  g539(.A1(new_n697), .A2(new_n422), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n726), .A2(new_n715), .A3(new_n292), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n692), .A2(KEYINPUT28), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n517), .B1(new_n728), .B2(new_n548), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n528), .B2(new_n542), .ZN(new_n730));
  OAI21_X1  g544(.A(KEYINPUT100), .B1(new_n730), .B2(new_n552), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n728), .A2(new_n548), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n534), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n556), .B2(new_n557), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n551), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n625), .A2(new_n628), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n727), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NOR3_X1   g553(.A1(new_n651), .A2(new_n715), .A3(new_n701), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n628), .A2(new_n731), .A3(new_n736), .A4(new_n703), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT101), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n741), .A2(new_n742), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  AOI21_X1  g560(.A(new_n624), .B1(new_n581), .B2(new_n584), .ZN(new_n747));
  INV_X1    g561(.A(G469), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n488), .A2(KEYINPUT102), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT102), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n479), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n751), .A3(new_n484), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n748), .B1(new_n752), .B2(new_n414), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n496), .A2(G469), .A3(G902), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n430), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n424), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n416), .A2(new_n421), .A3(new_n756), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n755), .A2(new_n701), .A3(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n747), .A2(KEYINPUT42), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n578), .A2(new_n585), .A3(new_n625), .A4(new_n758), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n760), .A2(KEYINPUT103), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT103), .B1(new_n760), .B2(new_n761), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(KEYINPUT104), .B(G131), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G33));
  NOR3_X1   g580(.A1(new_n755), .A2(new_n682), .A3(new_n757), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n578), .A2(new_n585), .A3(new_n625), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  INV_X1    g583(.A(KEYINPUT106), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT43), .B1(new_n632), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n632), .A2(new_n642), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT107), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n671), .A3(new_n703), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT108), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n757), .B1(new_n775), .B2(new_n776), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n752), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n480), .A2(new_n489), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n782), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n748), .A2(new_n414), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(KEYINPUT46), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n497), .A3(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(new_n430), .A3(new_n686), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT105), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n780), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n430), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n702), .A2(new_n624), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n757), .B(new_n797), .C1(new_n578), .C2(new_n585), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  NOR4_X1   g614(.A1(new_n624), .A2(new_n772), .A3(new_n667), .A4(new_n425), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT110), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n497), .A2(new_n714), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n802), .B1(KEYINPUT49), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n695), .ZN(new_n806));
  INV_X1    g620(.A(new_n696), .ZN(new_n807));
  OR2_X1    g621(.A1(new_n804), .A2(KEYINPUT49), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n758), .B1(new_n743), .B2(new_n744), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n231), .A2(new_n681), .ZN(new_n811));
  NOR4_X1   g625(.A1(new_n757), .A2(new_n656), .A3(new_n674), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n578), .A2(new_n670), .A3(new_n812), .A4(new_n585), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n768), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n764), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n717), .A2(new_n720), .A3(new_n724), .A4(new_n738), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n578), .A2(new_n585), .A3(new_n625), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n666), .A2(new_n670), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n283), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n282), .A2(new_n640), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n293), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n824), .B1(new_n664), .B2(new_n665), .ZN(new_n825));
  INV_X1    g639(.A(new_n630), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n825), .A2(new_n670), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n676), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n821), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n501), .A2(new_n675), .B1(new_n631), .B2(new_n825), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT111), .B1(new_n831), .B2(new_n626), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n818), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n816), .A2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n726), .A2(new_n755), .A3(new_n680), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n674), .A3(new_n695), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n745), .A2(new_n684), .A3(new_n836), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n837), .A2(new_n711), .A3(KEYINPUT52), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(new_n837), .B2(new_n711), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT112), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n711), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n837), .A2(new_n711), .A3(KEYINPUT52), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n834), .A2(new_n840), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n745), .A2(new_n684), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n711), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n764), .B1(new_n853), .B2(new_n839), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n817), .A2(new_n814), .A3(new_n848), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n829), .B1(new_n821), .B2(new_n828), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n831), .A2(new_n626), .A3(KEYINPUT111), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n850), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n855), .A2(new_n858), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n711), .A2(new_n851), .A3(new_n852), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n745), .A2(new_n684), .A3(new_n836), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n710), .B2(new_n707), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n864), .B2(KEYINPUT52), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n861), .A2(KEYINPUT114), .A3(new_n865), .A4(new_n764), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n860), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n849), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n847), .A2(new_n848), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT53), .B1(new_n834), .B2(new_n865), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n874), .B1(new_n871), .B2(new_n870), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n869), .B1(new_n875), .B2(KEYINPUT54), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n773), .A2(new_n288), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT115), .Z(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n737), .ZN(new_n880));
  NOR4_X1   g694(.A1(new_n880), .A2(new_n756), .A3(new_n696), .A4(new_n715), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT50), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n715), .A2(new_n757), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n806), .A2(new_n625), .A3(new_n288), .A4(new_n883), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n282), .A3(new_n642), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n879), .A2(new_n883), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n743), .A2(new_n744), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(new_n796), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n804), .A2(new_n430), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT116), .Z(new_n892));
  AOI211_X1 g706(.A(new_n757), .B(new_n880), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n877), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n880), .A2(new_n757), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n895), .B1(new_n796), .B2(new_n891), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n882), .A2(KEYINPUT51), .A3(new_n888), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n645), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n285), .B1(new_n884), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n886), .A2(new_n747), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT48), .Z(new_n901));
  INV_X1    g715(.A(new_n880), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n899), .B(new_n901), .C1(new_n722), .C2(new_n902), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n876), .A2(new_n894), .A3(new_n897), .A4(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(G952), .A2(G953), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n809), .B1(new_n904), .B2(new_n905), .ZN(G75));
  NOR2_X1   g720(.A1(new_n284), .A2(G952), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n414), .B1(new_n849), .B2(new_n867), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT56), .B1(new_n908), .B2(G210), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n418), .A2(new_n419), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n335), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(new_n420), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT55), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT117), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n908), .B(KEYINPUT118), .Z(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n298), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n914), .A2(KEYINPUT119), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n914), .A2(KEYINPUT119), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT56), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n907), .B(new_n916), .C1(new_n918), .C2(new_n921), .ZN(G51));
  NAND2_X1  g736(.A1(new_n917), .A2(new_n784), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT121), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n868), .B(KEYINPUT54), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n785), .B(KEYINPUT57), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n496), .B1(new_n927), .B2(KEYINPUT120), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(KEYINPUT120), .B2(new_n927), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n907), .B1(new_n924), .B2(new_n929), .ZN(G54));
  NAND3_X1  g744(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n931));
  INV_X1    g745(.A(new_n271), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n907), .ZN(G60));
  OR2_X1    g749(.A1(new_n635), .A2(new_n636), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n638), .B(KEYINPUT59), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n876), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n907), .B1(new_n925), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(G63));
  INV_X1    g755(.A(new_n907), .ZN(new_n942));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n849), .B2(new_n867), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(new_n621), .ZN(new_n946));
  INV_X1    g760(.A(new_n944), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n868), .A2(new_n673), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n949));
  OR3_X1    g763(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n948), .B1(new_n946), .B2(KEYINPUT122), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n953), .B(new_n942), .C1(new_n945), .C2(new_n621), .ZN(new_n954));
  AOI211_X1 g768(.A(new_n951), .B(KEYINPUT61), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n621), .B1(new_n868), .B2(new_n947), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT122), .B1(new_n956), .B2(new_n907), .ZN(new_n957));
  INV_X1    g771(.A(new_n948), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT123), .B1(new_n959), .B2(new_n949), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n950), .B1(new_n955), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT124), .B(new_n950), .C1(new_n955), .C2(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(G66));
  OAI21_X1  g779(.A(G953), .B1(new_n291), .B2(new_n332), .ZN(new_n966));
  INV_X1    g780(.A(new_n833), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(G953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n910), .B1(G898), .B2(new_n284), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT125), .Z(new_n970));
  XNOR2_X1  g784(.A(new_n968), .B(new_n970), .ZN(G69));
  NAND4_X1  g785(.A1(new_n791), .A2(new_n422), .A3(new_n697), .A4(new_n747), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n711), .A2(new_n851), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n799), .A2(new_n768), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n972), .A2(new_n792), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n764), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n284), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n284), .A2(G900), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n570), .B(new_n268), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n973), .A2(new_n699), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n991));
  INV_X1    g805(.A(new_n799), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n822), .A2(new_n823), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT126), .Z(new_n994));
  NOR4_X1   g808(.A1(new_n819), .A2(new_n994), .A3(new_n687), .A4(new_n757), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n792), .A2(new_n990), .A3(new_n991), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n985), .B1(new_n997), .B2(new_n284), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n986), .A2(new_n988), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n984), .B1(new_n981), .B2(new_n982), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n987), .B1(new_n1001), .B2(new_n998), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1000), .A2(new_n1002), .ZN(G72));
  NOR2_X1   g817(.A1(new_n571), .A2(new_n517), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n975), .A2(new_n976), .A3(new_n833), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G472), .A2(G902), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT63), .Z(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1004), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1007), .B1(new_n997), .B2(new_n833), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n517), .A3(new_n571), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1009), .A2(new_n1011), .A3(new_n942), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n690), .A2(new_n565), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1012), .B1(new_n875), .B2(new_n1014), .ZN(G57));
endmodule


