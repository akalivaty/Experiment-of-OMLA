//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n833, new_n834,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953;
  XNOR2_X1  g000(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n202));
  INV_X1    g001(.A(G127gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G134gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT68), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT67), .B(G134gat), .Z(new_n206));
  OAI21_X1  g005(.A(new_n205), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n207), .B1(KEYINPUT1), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT2), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g013(.A(KEYINPUT76), .B(G148gat), .Z(new_n215));
  AND2_X1   g014(.A1(new_n215), .A2(G141gat), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n217), .A2(G148gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n210), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(new_n213), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G113gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(KEYINPUT69), .A3(G120gat), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n203), .A2(G134gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT1), .B1(new_n203), .B2(G134gat), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n226), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n209), .A2(new_n219), .A3(new_n224), .A4(new_n231), .ZN(new_n232));
  MUX2_X1   g031(.A(new_n202), .B(KEYINPUT4), .S(new_n232), .Z(new_n233));
  NAND2_X1  g032(.A1(new_n219), .A2(new_n224), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT77), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT77), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n238), .B1(new_n234), .B2(KEYINPUT3), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n209), .A2(new_n231), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(KEYINPUT3), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT5), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n233), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n234), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n232), .ZN(new_n249));
  AND3_X1   g048(.A1(new_n249), .A2(KEYINPUT79), .A3(new_n245), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT79), .B1(new_n249), .B2(new_n245), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n209), .A2(new_n231), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n235), .ZN(new_n254));
  INV_X1    g053(.A(new_n232), .ZN(new_n255));
  INV_X1    g054(.A(new_n202), .ZN(new_n256));
  OAI211_X1 g055(.A(new_n254), .B(new_n244), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n241), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n239), .B2(new_n237), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT5), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n247), .B1(new_n252), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G1gat), .B(G29gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT0), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n263), .B(new_n264), .Z(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n261), .A2(KEYINPUT6), .A3(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n261), .B2(new_n266), .ZN(new_n269));
  OAI221_X1 g068(.A(KEYINPUT5), .B1(new_n257), .B2(new_n259), .C1(new_n250), .C2(new_n251), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n265), .B1(new_n270), .B2(new_n247), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n267), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT30), .ZN(new_n273));
  NOR2_X1   g072(.A1(G169gat), .A2(G176gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT26), .ZN(new_n276));
  INV_X1    g075(.A(G169gat), .ZN(new_n277));
  INV_X1    g076(.A(G176gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n275), .B1(new_n279), .B2(KEYINPUT26), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n281), .B2(new_n280), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT65), .B(KEYINPUT28), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT27), .B(G183gat), .Z(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT64), .ZN(new_n287));
  INV_X1    g086(.A(G183gat), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT64), .B1(new_n288), .B2(KEYINPUT27), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(G190gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n285), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n286), .A2(new_n292), .A3(G190gat), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n283), .B(new_n284), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT23), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n274), .B(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n284), .A2(KEYINPUT24), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(new_n279), .ZN(new_n298));
  OR2_X1    g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n299), .A2(KEYINPUT24), .A3(new_n284), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G226gat), .A2(G233gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n294), .B2(new_n303), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(KEYINPUT22), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G211gat), .B(G218gat), .ZN(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n315), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n306), .B(new_n317), .C1(new_n305), .C2(new_n307), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G8gat), .B(G36gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(G64gat), .B(G92gat), .ZN(new_n321));
  XOR2_X1   g120(.A(new_n320), .B(new_n321), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n273), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(new_n322), .B(KEYINPUT72), .Z(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n316), .B2(new_n318), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n319), .A2(new_n323), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n330), .A2(new_n331), .B1(KEYINPUT30), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n272), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n236), .B1(new_n315), .B2(KEYINPUT29), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n234), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT29), .B1(new_n237), .B2(new_n239), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n317), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G22gat), .ZN(new_n339));
  INV_X1    g138(.A(G22gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(new_n336), .C1(new_n337), .C2(new_n317), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n336), .A2(new_n343), .B1(G228gat), .B2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT80), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n339), .A2(new_n344), .A3(new_n341), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT31), .B(G50gat), .ZN(new_n351));
  INV_X1    g150(.A(new_n349), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n346), .A2(new_n352), .A3(new_n347), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n351), .ZN(new_n355));
  INV_X1    g154(.A(new_n353), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n346), .B2(new_n347), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n334), .B1(new_n354), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT36), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n294), .A2(new_n241), .A3(new_n303), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n241), .B1(new_n294), .B2(new_n303), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G227gat), .ZN(new_n365));
  INV_X1    g164(.A(G233gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n364), .A2(KEYINPUT34), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT34), .ZN(new_n369));
  INV_X1    g168(.A(new_n363), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  INV_X1    g170(.A(new_n367), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n369), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n364), .A2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT70), .B(G71gat), .ZN(new_n378));
  INV_X1    g177(.A(G99gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n378), .B(new_n379), .ZN(new_n380));
  XOR2_X1   g179(.A(G15gat), .B(G43gat), .Z(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NAND2_X1  g181(.A1(new_n377), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n374), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n377), .B(new_n382), .C1(new_n368), .C2(new_n373), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n375), .A2(KEYINPUT32), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n387), .B1(new_n384), .B2(new_n385), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n360), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI211_X1 g192(.A(KEYINPUT71), .B(KEYINPUT36), .C1(new_n389), .C2(new_n390), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n359), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(new_n265), .B(KEYINPUT82), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(new_n270), .B2(new_n247), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n255), .A2(new_n256), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(KEYINPUT4), .B2(new_n255), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n245), .B1(new_n400), .B2(new_n259), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT83), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT83), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n403), .B(new_n245), .C1(new_n400), .C2(new_n259), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT39), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n248), .A2(new_n244), .A3(new_n232), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n402), .A2(new_n404), .A3(KEYINPUT39), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n397), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT40), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n398), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n326), .A2(new_n333), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n407), .A2(KEYINPUT40), .A3(new_n409), .A4(new_n397), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n269), .A2(new_n398), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n319), .A2(KEYINPUT37), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n417), .A2(KEYINPUT38), .A3(new_n328), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n319), .A2(KEYINPUT37), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n332), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n419), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n323), .B1(new_n319), .B2(KEYINPUT37), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT38), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n416), .A2(new_n420), .A3(new_n267), .A4(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n415), .A2(new_n354), .A3(new_n358), .A4(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n267), .B1(new_n269), .B2(new_n398), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n426), .A2(new_n326), .A3(new_n333), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT84), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n426), .A2(new_n326), .A3(KEYINPUT84), .A4(new_n333), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n358), .A2(new_n354), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT85), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n389), .B2(new_n390), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n384), .A2(new_n385), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n386), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n436), .A2(KEYINPUT85), .A3(new_n388), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT35), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n431), .A2(new_n432), .A3(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n334), .A2(new_n358), .A3(new_n354), .A4(new_n391), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT35), .ZN(new_n442));
  AOI22_X1  g241(.A1(new_n396), .A2(new_n425), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444));
  OR2_X1    g243(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n446));
  AOI21_X1  g245(.A(G36gat), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(G29gat), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n448), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n444), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(G43gat), .A2(G50gat), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT15), .ZN(new_n452));
  NAND2_X1  g251(.A1(G43gat), .A2(G50gat), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n447), .B2(new_n449), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI221_X1 g257(.A(new_n454), .B1(new_n456), .B2(new_n444), .C1(new_n447), .C2(new_n449), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(KEYINPUT89), .A2(G1gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(KEYINPUT89), .A2(G1gat), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT16), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT90), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n467), .B(KEYINPUT16), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n469), .A2(KEYINPUT88), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n466), .B(new_n468), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G8gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n472), .ZN(new_n475));
  INV_X1    g274(.A(G1gat), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n470), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n473), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n474), .B1(new_n473), .B2(new_n477), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n461), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(new_n460), .A3(new_n478), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT93), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT93), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n461), .B(new_n485), .C1(new_n479), .C2(new_n480), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n488), .B(KEYINPUT92), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT13), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT91), .B1(new_n479), .B2(new_n480), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n482), .A2(new_n492), .A3(new_n478), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n460), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT17), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n491), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n489), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n481), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT18), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n487), .A2(new_n490), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n498), .A2(KEYINPUT18), .A3(new_n499), .A4(new_n481), .ZN(new_n503));
  XNOR2_X1  g302(.A(G113gat), .B(G141gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G169gat), .B(G197gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(KEYINPUT12), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n502), .A2(KEYINPUT94), .A3(new_n503), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n500), .A2(new_n501), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n484), .A2(new_n490), .A3(new_n486), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n511), .A2(new_n503), .A3(new_n512), .A4(new_n509), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT94), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n502), .A2(new_n503), .ZN(new_n516));
  INV_X1    g315(.A(new_n509), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n510), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G230gat), .A2(G233gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT95), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G71gat), .B2(G78gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n527), .ZN(new_n529));
  OR2_X1    g328(.A1(G57gat), .A2(G64gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G57gat), .A2(G64gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n530), .B(new_n531), .C1(new_n525), .C2(KEYINPUT9), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n532), .A3(new_n521), .ZN(new_n533));
  AND2_X1   g332(.A1(new_n528), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT7), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(KEYINPUT99), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT8), .ZN(new_n541));
  INV_X1    g340(.A(G85gat), .ZN(new_n542));
  INV_X1    g341(.A(G92gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n537), .A2(new_n539), .A3(new_n541), .A4(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G99gat), .B(G106gat), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(KEYINPUT102), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT102), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n545), .B2(new_n547), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n537), .A2(new_n539), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT100), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n546), .A4(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT100), .B1(new_n545), .B2(new_n547), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT101), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n556), .B2(new_n557), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n534), .B(new_n552), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n556), .A2(new_n557), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT103), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n545), .A2(new_n563), .A3(new_n547), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n548), .A2(KEYINPUT103), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n562), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n528), .A2(new_n533), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT10), .B1(new_n561), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n552), .B1(new_n559), .B2(new_n560), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n528), .A2(new_n533), .A3(KEYINPUT96), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n519), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT104), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(KEYINPUT104), .B(new_n519), .C1(new_n569), .C2(new_n575), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n561), .A2(new_n568), .ZN(new_n581));
  INV_X1    g380(.A(new_n519), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G120gat), .B(G148gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n576), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n587), .B1(new_n590), .B2(new_n583), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  INV_X1    g396(.A(G231gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n534), .B(new_n597), .C1(new_n598), .C2(new_n366), .ZN(new_n599));
  OAI211_X1 g398(.A(G231gat), .B(G233gat), .C1(new_n567), .C2(KEYINPUT21), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n203), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n203), .B1(new_n599), .B2(new_n600), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n596), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  INV_X1    g404(.A(new_n596), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(new_n606), .A3(new_n601), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  INV_X1    g407(.A(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n604), .B2(new_n607), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n572), .A2(new_n573), .ZN(new_n614));
  AOI211_X1 g413(.A(new_n480), .B(new_n479), .C1(new_n614), .C2(KEYINPUT21), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n604), .A2(new_n607), .ZN(new_n618));
  INV_X1    g417(.A(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n620), .B2(new_n611), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n595), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n615), .B1(new_n612), .B2(new_n613), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n617), .A3(new_n611), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n623), .A2(new_n594), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n570), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n461), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n497), .A2(new_n570), .ZN(new_n628));
  AND2_X1   g427(.A1(G232gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n627), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n629), .A2(KEYINPUT41), .ZN(new_n634));
  XNOR2_X1  g433(.A(G134gat), .B(G162gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n633), .B(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n593), .A2(new_n622), .A3(new_n625), .A4(new_n638), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n443), .A2(new_n518), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n272), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n413), .ZN(new_n644));
  OR2_X1    g443(.A1(new_n644), .A2(KEYINPUT105), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(KEYINPUT105), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(G8gat), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT42), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT16), .B(G8gat), .ZN(new_n649));
  OR3_X1    g448(.A1(new_n644), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n649), .B1(new_n645), .B2(new_n646), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n647), .B(new_n650), .C1(new_n651), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g451(.A(G15gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n434), .A2(new_n437), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n640), .A2(new_n395), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n653), .ZN(G1326gat));
  NAND2_X1  g457(.A1(new_n358), .A2(new_n354), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n640), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT43), .B(G22gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(G1327gat));
  NOR2_X1   g461(.A1(new_n443), .A2(new_n518), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n622), .A2(new_n625), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n638), .A3(new_n592), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n641), .A2(new_n448), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n667), .A2(KEYINPUT106), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(KEYINPUT106), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n669), .A2(KEYINPUT45), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT45), .B1(new_n669), .B2(new_n670), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT44), .B1(new_n443), .B2(new_n638), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n440), .A2(new_n442), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n393), .A2(new_n394), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n659), .B1(new_n641), .B2(new_n413), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n425), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n680));
  INV_X1    g479(.A(new_n638), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n674), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n638), .B1(new_n675), .B2(new_n678), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n680), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n665), .A2(new_n518), .A3(new_n592), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n641), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G29gat), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n690), .ZN(G1328gat));
  INV_X1    g490(.A(new_n667), .ZN(new_n692));
  AOI21_X1  g491(.A(G36gat), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n413), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n413), .B(new_n688), .C1(new_n684), .C2(new_n686), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(G36gat), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n697), .A2(KEYINPUT110), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(G1329gat));
  OAI211_X1 g500(.A(new_n395), .B(new_n688), .C1(new_n684), .C2(new_n686), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(G43gat), .ZN(new_n703));
  OR3_X1    g502(.A1(new_n667), .A2(G43gat), .A3(new_n654), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n703), .A2(KEYINPUT47), .A3(new_n704), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(G1330gat));
  OAI211_X1 g508(.A(new_n659), .B(new_n688), .C1(new_n684), .C2(new_n686), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(G50gat), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT48), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT111), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n432), .A2(G50gat), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n692), .A2(new_n714), .B1(KEYINPUT111), .B2(new_n712), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n711), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n711), .B2(new_n715), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n516), .A2(new_n517), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n513), .A2(new_n514), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n513), .A2(new_n514), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n719), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR4_X1   g521(.A1(new_n664), .A2(new_n722), .A3(new_n681), .A4(new_n593), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n679), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n641), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(G57gat), .ZN(G1332gat));
  INV_X1    g525(.A(KEYINPUT112), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n679), .A2(new_n723), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT112), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT113), .ZN(new_n733));
  INV_X1    g532(.A(new_n413), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n734), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n732), .B2(new_n735), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n736), .A2(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT113), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n743), .ZN(G1333gat));
  OAI21_X1  g543(.A(G71gat), .B1(new_n731), .B2(new_n676), .ZN(new_n745));
  OR3_X1    g544(.A1(new_n729), .A2(G71gat), .A3(new_n654), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1334gat));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n659), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g550(.A1(new_n665), .A2(new_n722), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n593), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n687), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(G85gat), .B1(new_n755), .B2(new_n272), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n685), .A2(KEYINPUT51), .A3(new_n752), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT51), .B1(new_n685), .B2(new_n752), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n592), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n641), .A2(new_n542), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n756), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  OAI211_X1 g560(.A(new_n413), .B(new_n754), .C1(new_n684), .C2(new_n686), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G92gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n734), .A2(G92gat), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n763), .B(new_n768), .C1(new_n759), .C2(new_n765), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n755), .B2(new_n676), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n655), .A2(new_n379), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n759), .B2(new_n772), .ZN(G1338gat));
  OAI211_X1 g572(.A(new_n659), .B(new_n754), .C1(new_n684), .C2(new_n686), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G106gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT114), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n432), .A2(G106gat), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n592), .B(new_n777), .C1(new_n757), .C2(new_n758), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n779), .A3(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n775), .B(new_n778), .C1(KEYINPUT114), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1339gat));
  OAI21_X1  g582(.A(new_n587), .B1(new_n576), .B2(KEYINPUT54), .ZN(new_n784));
  AND3_X1   g583(.A1(new_n578), .A2(KEYINPUT54), .A3(new_n579), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n569), .A2(new_n575), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n582), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT116), .ZN(new_n788));
  NOR4_X1   g587(.A1(new_n569), .A2(new_n575), .A3(KEYINPUT116), .A4(new_n519), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n785), .A2(new_n791), .A3(KEYINPUT117), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n786), .B2(new_n582), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n789), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n578), .A2(KEYINPUT54), .A3(new_n579), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n793), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n784), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n799), .A2(KEYINPUT55), .B1(new_n580), .B2(new_n588), .ZN(new_n800));
  INV_X1    g599(.A(new_n784), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT117), .B1(new_n785), .B2(new_n791), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n796), .A2(new_n797), .A3(new_n793), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n487), .A2(new_n490), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n498), .A2(new_n481), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n489), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n510), .A2(new_n515), .B1(new_n508), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n800), .A2(new_n806), .A3(new_n681), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n811), .A2(new_n592), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n518), .B1(new_n804), .B2(new_n805), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n800), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n812), .B1(new_n815), .B2(new_n681), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n664), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n622), .A2(new_n625), .A3(new_n638), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n818), .A2(new_n819), .A3(new_n518), .A4(new_n593), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT115), .B1(new_n639), .B2(new_n722), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n817), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n659), .A2(new_n389), .A3(new_n390), .ZN(new_n824));
  AND4_X1   g623(.A1(new_n641), .A2(new_n823), .A3(new_n734), .A4(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825), .B2(new_n722), .ZN(new_n826));
  INV_X1    g625(.A(new_n822), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n816), .B2(new_n664), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n734), .A2(new_n641), .ZN(new_n829));
  NOR4_X1   g628(.A1(new_n828), .A2(new_n659), .A3(new_n654), .A4(new_n829), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n518), .A2(new_n227), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n826), .B1(new_n830), .B2(new_n831), .ZN(G1340gat));
  AOI21_X1  g631(.A(G120gat), .B1(new_n825), .B2(new_n592), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n592), .A2(G120gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n830), .B2(new_n834), .ZN(G1341gat));
  NAND3_X1  g634(.A1(new_n825), .A2(new_n203), .A3(new_n665), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n830), .A2(new_n665), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n203), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT118), .ZN(G1342gat));
  INV_X1    g638(.A(new_n206), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n840), .A3(new_n681), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n830), .A2(new_n681), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(G134gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n842), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NOR2_X1   g645(.A1(new_n395), .A2(new_n829), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n659), .A2(KEYINPUT57), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n815), .B2(new_n681), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n811), .A2(new_n592), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n589), .B1(new_n804), .B2(new_n805), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n722), .B1(new_n799), .B2(KEYINPUT55), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(KEYINPUT119), .A3(new_n638), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n850), .A2(new_n812), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n664), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n848), .B1(new_n857), .B2(new_n822), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n823), .B2(new_n659), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n847), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G141gat), .B1(new_n860), .B2(new_n518), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n676), .A2(new_n659), .ZN(new_n862));
  NOR4_X1   g661(.A1(new_n828), .A2(new_n272), .A3(new_n413), .A4(new_n862), .ZN(new_n863));
  AND3_X1   g662(.A1(new_n863), .A2(new_n217), .A3(new_n722), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n864), .A2(KEYINPUT58), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n860), .A2(KEYINPUT120), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n828), .B2(new_n432), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n827), .B1(new_n856), .B2(new_n664), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n869), .B1(new_n870), .B2(new_n848), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n847), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n867), .A2(new_n722), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n864), .B1(new_n874), .B2(G141gat), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n866), .B1(new_n875), .B2(new_n876), .ZN(G1344gat));
  NAND3_X1  g676(.A1(new_n818), .A2(new_n518), .A3(new_n593), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n432), .B1(new_n817), .B2(new_n878), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n879), .A2(KEYINPUT57), .B1(new_n828), .B2(new_n848), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n395), .A2(new_n593), .A3(new_n829), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n880), .A2(KEYINPUT121), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(G148gat), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT121), .B1(new_n880), .B2(new_n881), .ZN(new_n884));
  OAI21_X1  g683(.A(KEYINPUT59), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g684(.A1(new_n871), .A2(new_n872), .A3(new_n847), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n872), .B1(new_n871), .B2(new_n847), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n886), .A2(new_n887), .A3(new_n593), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n215), .A2(KEYINPUT59), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n885), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n863), .A2(new_n215), .A3(new_n592), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1345gat));
  NAND3_X1  g691(.A1(new_n863), .A2(new_n609), .A3(new_n665), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n886), .A2(new_n887), .A3(new_n664), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n609), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n863), .B2(new_n681), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n886), .A2(new_n887), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n681), .A2(G162gat), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n734), .A2(new_n641), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n823), .A2(new_n432), .A3(new_n655), .A4(new_n900), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n901), .A2(new_n277), .A3(new_n518), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n824), .A2(new_n413), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n823), .A2(KEYINPUT122), .A3(new_n272), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT122), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n828), .B2(new_n641), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n722), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n908), .B2(new_n277), .ZN(G1348gat));
  NAND3_X1  g708(.A1(new_n907), .A2(new_n278), .A3(new_n592), .ZN(new_n910));
  OAI21_X1  g709(.A(G176gat), .B1(new_n901), .B2(new_n593), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT123), .ZN(G1349gat));
  OAI21_X1  g712(.A(G183gat), .B1(new_n901), .B2(new_n664), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n664), .A2(new_n286), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n907), .A2(KEYINPUT124), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(KEYINPUT124), .B1(new_n907), .B2(new_n915), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT60), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n920));
  OAI211_X1 g719(.A(new_n920), .B(new_n914), .C1(new_n916), .C2(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1350gat));
  INV_X1    g721(.A(G190gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n923), .A3(new_n681), .ZN(new_n924));
  OAI21_X1  g723(.A(G190gat), .B1(new_n901), .B2(new_n638), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(KEYINPUT61), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  AOI211_X1 g727(.A(new_n734), .B(new_n862), .C1(new_n904), .C2(new_n906), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT125), .ZN(new_n930));
  XNOR2_X1  g729(.A(KEYINPUT126), .B(G197gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(KEYINPUT125), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n930), .A2(new_n722), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n880), .A2(new_n676), .A3(new_n900), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(new_n518), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(new_n931), .ZN(G1352gat));
  INV_X1    g735(.A(G204gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n929), .A2(new_n937), .A3(new_n592), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n939));
  OAI21_X1  g738(.A(G204gat), .B1(new_n934), .B2(new_n593), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(G1353gat));
  NAND4_X1  g741(.A1(new_n930), .A2(new_n310), .A3(new_n665), .A4(new_n932), .ZN(new_n943));
  OAI21_X1  g742(.A(G211gat), .B1(new_n934), .B2(new_n664), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n944), .A2(new_n945), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1354gat));
  NAND4_X1  g747(.A1(new_n930), .A2(new_n311), .A3(new_n681), .A4(new_n932), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n681), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n952));
  OAI21_X1  g751(.A(G218gat), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n949), .A2(new_n953), .ZN(G1355gat));
endmodule


