//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT75), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n204), .B2(new_n206), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n203), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT76), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  INV_X1    g010(.A(KEYINPUT76), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n212), .B(new_n203), .C1(new_n207), .C2(new_n208), .ZN(new_n213));
  AND3_X1   g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(new_n210), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n202), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n211), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n218), .B(new_n205), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n212), .B1(new_n219), .B2(new_n203), .ZN(new_n220));
  INV_X1    g019(.A(new_n213), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT77), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n216), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G226gat), .A2(G233gat), .ZN(new_n227));
  XOR2_X1   g026(.A(new_n227), .B(KEYINPUT78), .Z(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n231), .B1(KEYINPUT23), .B2(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT65), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n232), .A2(new_n237), .A3(KEYINPUT23), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT66), .ZN(new_n240));
  NOR2_X1   g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(G183gat), .A2(G190gat), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT24), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n241), .B1(new_n244), .B2(KEYINPUT64), .ZN(new_n245));
  NAND3_X1  g044(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n245), .B(new_n246), .C1(KEYINPUT64), .C2(new_n244), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n233), .B(new_n248), .C1(new_n236), .C2(new_n238), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n240), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n230), .C1(new_n234), .C2(new_n235), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT25), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n230), .B1(new_n234), .B2(new_n235), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n234), .A2(KEYINPUT65), .A3(new_n235), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n237), .B1(new_n232), .B2(KEYINPUT23), .ZN(new_n259));
  AOI22_X1  g058(.A1(KEYINPUT67), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(G183gat), .B2(G190gat), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n244), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  AOI22_X1  g064(.A1(KEYINPUT24), .A2(new_n265), .B1(new_n241), .B2(KEYINPUT68), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n261), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  INV_X1    g067(.A(G190gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT68), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n244), .A2(new_n270), .A3(new_n263), .A4(new_n246), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n256), .B(new_n260), .C1(new_n267), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n264), .A2(new_n266), .A3(new_n261), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(KEYINPUT69), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n255), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT70), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n278), .A3(new_n260), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n252), .A2(new_n274), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT28), .ZN(new_n281));
  XNOR2_X1  g080(.A(KEYINPUT27), .B(G183gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(KEYINPUT72), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n283), .B2(new_n269), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n234), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n287));
  OR3_X1    g086(.A1(new_n287), .A2(new_n268), .A3(KEYINPUT27), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT27), .B1(new_n287), .B2(new_n268), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n288), .A2(new_n281), .A3(new_n269), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n234), .A2(new_n285), .A3(new_n230), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n242), .A3(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n284), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n229), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n227), .B1(new_n280), .B2(new_n294), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n226), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n229), .ZN(new_n300));
  INV_X1    g099(.A(new_n227), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n280), .B2(new_n294), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n300), .B(new_n225), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT79), .B(G64gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n304), .B(G92gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G8gat), .B(G36gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n303), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT80), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n299), .A2(KEYINPUT80), .A3(new_n303), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT30), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n308), .B1(new_n299), .B2(new_n303), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n309), .A2(new_n314), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT90), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G148gat), .ZN(new_n324));
  INV_X1    g123(.A(G148gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n325), .A2(G141gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n327), .B1(KEYINPUT83), .B2(KEYINPUT2), .ZN(new_n328));
  AND2_X1   g127(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n324), .A2(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(new_n327), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n330), .A2(new_n332), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT84), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n330), .A2(new_n336), .A3(new_n332), .A4(KEYINPUT84), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n324), .A2(new_n326), .ZN(new_n342));
  OR3_X1    g141(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n342), .B1(new_n331), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT3), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n341), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G127gat), .B(G134gat), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n347), .A2(new_n349), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n344), .B1(new_n339), .B2(new_n340), .ZN(new_n361));
  INV_X1    g160(.A(new_n357), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT86), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n346), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n360), .B(new_n363), .C1(new_n367), .C2(KEYINPUT4), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n361), .A2(new_n362), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT85), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n361), .ZN(new_n374));
  OR3_X1    g173(.A1(new_n374), .A2(KEYINPUT91), .A3(new_n370), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT91), .B1(new_n374), .B2(new_n370), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(KEYINPUT39), .A3(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n371), .A2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G1gat), .B(G29gat), .Z(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(G85gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT0), .B(G57gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n370), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(KEYINPUT39), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n378), .A2(new_n385), .A3(KEYINPUT40), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n378), .A2(new_n385), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n388));
  AOI211_X1 g187(.A(new_n364), .B(new_n344), .C1(new_n339), .C2(new_n340), .ZN(new_n389));
  OAI211_X1 g188(.A(KEYINPUT4), .B(new_n362), .C1(new_n388), .C2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n372), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n390), .A2(new_n360), .A3(new_n369), .A4(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT5), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n374), .B2(new_n370), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n362), .B1(new_n388), .B2(new_n389), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n391), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n370), .A2(KEYINPUT5), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n360), .A3(new_n363), .A4(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n383), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n387), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n386), .B1(new_n402), .B2(KEYINPUT40), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT30), .B1(new_n311), .B2(new_n312), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n405), .A2(new_n316), .A3(new_n318), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT90), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n322), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n396), .A2(new_n400), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n382), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n400), .A3(new_n383), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n410), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(KEYINPUT6), .A3(new_n382), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n299), .A2(KEYINPUT37), .A3(new_n303), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT37), .B1(new_n299), .B2(new_n303), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n307), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT93), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(KEYINPUT38), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT37), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n275), .A2(new_n276), .ZN(new_n424));
  AND4_X1   g223(.A1(new_n278), .A2(new_n424), .A3(new_n256), .A4(new_n260), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n278), .B1(new_n277), .B2(new_n260), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n293), .B1(new_n427), .B2(new_n252), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n228), .B1(new_n428), .B2(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n295), .A2(new_n301), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n225), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n301), .B1(new_n295), .B2(new_n296), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n228), .B1(new_n280), .B2(new_n294), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n432), .A2(new_n226), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n423), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n299), .A2(KEYINPUT37), .A3(new_n303), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n308), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT93), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT92), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(new_n226), .C1(new_n432), .C2(new_n433), .ZN(new_n441));
  INV_X1    g240(.A(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n440), .B1(new_n443), .B2(new_n226), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n430), .B(new_n225), .C1(new_n229), .C2(new_n302), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT37), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n442), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n438), .B(new_n307), .C1(new_n447), .C2(new_n418), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n422), .A2(new_n439), .A3(new_n313), .A4(new_n448), .ZN(new_n449));
  XNOR2_X1  g248(.A(KEYINPUT88), .B(G22gat), .ZN(new_n450));
  AOI211_X1 g249(.A(KEYINPUT3), .B(new_n344), .C1(new_n339), .C2(new_n340), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n216), .B(new_n224), .C1(new_n451), .C2(KEYINPUT29), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT29), .B1(new_n222), .B2(new_n223), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n346), .B1(new_n453), .B2(KEYINPUT3), .ZN(new_n454));
  NAND2_X1  g253(.A1(G228gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT87), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT29), .B1(new_n361), .B2(new_n348), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n225), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n365), .B(new_n366), .C1(KEYINPUT3), .C2(new_n453), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n349), .A2(new_n296), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n462), .A2(KEYINPUT87), .A3(new_n224), .A4(new_n216), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  AOI211_X1 g263(.A(new_n450), .B(new_n457), .C1(new_n455), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n455), .ZN(new_n466));
  INV_X1    g265(.A(new_n457), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n465), .B1(G22gat), .B2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(G78gat), .B(G106gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(KEYINPUT31), .B(G50gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n468), .A2(new_n450), .ZN(new_n475));
  INV_X1    g274(.A(new_n450), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n466), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n472), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n476), .B1(new_n466), .B2(new_n467), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n474), .B(new_n479), .C1(new_n465), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n473), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n408), .A2(new_n449), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n479), .B1(new_n465), .B2(new_n481), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT89), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n487), .A2(new_n482), .B1(new_n472), .B2(new_n469), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n320), .B2(new_n416), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT73), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n295), .A2(new_n357), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n280), .A2(new_n362), .A3(new_n294), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G227gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT34), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n280), .A2(new_n362), .A3(new_n294), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n362), .B1(new_n280), .B2(new_n294), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT34), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n494), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n490), .B1(new_n496), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  XOR2_X1   g302(.A(G15gat), .B(G43gat), .Z(new_n504));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n494), .B1(new_n491), .B2(new_n492), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(KEYINPUT33), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AOI221_X4 g310(.A(new_n509), .B1(KEYINPUT33), .B2(new_n506), .C1(new_n493), .C2(new_n495), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n503), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT32), .B1(new_n499), .B2(new_n494), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n514), .B(new_n506), .C1(KEYINPUT33), .C2(new_n507), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n508), .A2(new_n510), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n502), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n513), .A2(KEYINPUT36), .A3(new_n517), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n493), .A2(KEYINPUT34), .A3(new_n495), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n500), .B1(new_n499), .B2(new_n494), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT74), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT74), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n496), .A2(new_n501), .A3(new_n522), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n521), .B(new_n523), .C1(new_n511), .C2(new_n512), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n496), .A2(new_n501), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT74), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT36), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n518), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n489), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n517), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n484), .A2(new_n415), .A3(new_n406), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT35), .ZN(new_n532));
  AOI221_X4 g331(.A(KEYINPUT35), .B1(new_n413), .B2(new_n414), .C1(new_n524), .C2(new_n526), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n316), .B1(new_n313), .B2(new_n314), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT90), .B1(new_n534), .B2(new_n319), .ZN(new_n535));
  NOR4_X1   g334(.A1(new_n405), .A2(new_n321), .A3(new_n316), .A4(new_n318), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n533), .B(new_n484), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n485), .A2(new_n529), .B1(new_n532), .B2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT95), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT15), .B1(new_n539), .B2(KEYINPUT97), .ZN(new_n543));
  INV_X1    g342(.A(G50gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G43gat), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(KEYINPUT97), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(G29gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(G36gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(G29gat), .A2(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n547), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT17), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n542), .A2(new_n553), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n553), .B1(new_n542), .B2(new_n546), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n554), .B1(KEYINPUT15), .B2(new_n541), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT17), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  INV_X1    g361(.A(G1gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT16), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G1gat), .B2(new_n562), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(G8gat), .Z(new_n567));
  NAND3_X1  g366(.A1(new_n558), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  OR3_X1    g367(.A1(new_n567), .A2(new_n559), .A3(new_n560), .ZN(new_n569));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n557), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n567), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n570), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT18), .A4(new_n570), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n573), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT94), .B(KEYINPUT11), .Z(new_n581));
  XNOR2_X1  g380(.A(G113gat), .B(G141gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G169gat), .B(G197gat), .Z(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT12), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n580), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n573), .A2(new_n578), .A3(new_n579), .A4(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n538), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT104), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G57gat), .B(G64gat), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G71gat), .B(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n596), .A2(KEYINPUT100), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n594), .B(KEYINPUT98), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G57gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G64gat), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n599), .B1(new_n608), .B2(KEYINPUT99), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(KEYINPUT99), .B2(new_n597), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n606), .A2(KEYINPUT101), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT101), .B1(new_n606), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n601), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT21), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n593), .B1(new_n615), .B2(new_n567), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n615), .A2(new_n593), .A3(new_n567), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n617), .A2(G231gat), .A3(G233gat), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n618), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n616), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n619), .B2(new_n622), .ZN(new_n627));
  XOR2_X1   g426(.A(G127gat), .B(G155gat), .Z(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT103), .B(KEYINPUT19), .Z(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n613), .A2(new_n614), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G183gat), .B(G211gat), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n613), .B2(new_n614), .ZN(new_n636));
  NOR3_X1   g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n635), .B1(new_n633), .B2(new_n636), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n629), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n638), .A2(new_n629), .A3(new_n639), .ZN(new_n641));
  OAI22_X1  g440(.A1(new_n626), .A2(new_n627), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n619), .A2(new_n622), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n623), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n645), .A3(new_n625), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT106), .B(G85gat), .Z(new_n648));
  INV_X1    g447(.A(G92gat), .ZN(new_n649));
  NAND2_X1  g448(.A1(G99gat), .A2(G106gat), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n648), .A2(new_n649), .B1(KEYINPUT8), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT105), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(G85gat), .A3(G92gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT7), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AND2_X1   g454(.A1(G99gat), .A2(G106gat), .ZN(new_n656));
  NOR2_X1   g455(.A1(G99gat), .A2(G106gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n651), .B(new_n654), .C1(new_n656), .C2(new_n657), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n558), .A2(new_n561), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n664));
  NAND2_X1  g463(.A1(G232gat), .A2(G233gat), .ZN(new_n665));
  OAI221_X1 g464(.A(new_n663), .B1(new_n664), .B2(new_n665), .C1(new_n574), .C2(new_n662), .ZN(new_n666));
  XNOR2_X1  g465(.A(G134gat), .B(G162gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(KEYINPUT107), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n666), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g468(.A(G190gat), .B(G218gat), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n665), .A2(new_n664), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n669), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n647), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(G230gat), .A2(G233gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n613), .A2(new_n662), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT10), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n661), .B(new_n601), .C1(new_n611), .C2(new_n612), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n678), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n676), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n679), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n683), .B2(new_n676), .ZN(new_n684));
  XNOR2_X1  g483(.A(KEYINPUT108), .B(G176gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(G120gat), .B(G148gat), .Z(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n684), .A2(new_n688), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n674), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n592), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n415), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n563), .ZN(G1324gat));
  NOR2_X1   g495(.A1(new_n535), .A2(new_n536), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT16), .B(G8gat), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n592), .A2(new_n697), .A3(new_n693), .A4(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT42), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n700), .A2(new_n701), .ZN(new_n704));
  INV_X1    g503(.A(new_n697), .ZN(new_n705));
  OAI21_X1  g504(.A(G8gat), .B1(new_n694), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(KEYINPUT109), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .A4(new_n707), .ZN(G1325gat));
  INV_X1    g507(.A(new_n694), .ZN(new_n709));
  INV_X1    g508(.A(new_n528), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n709), .A2(G15gat), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n524), .A2(new_n526), .ZN(new_n712));
  AOI21_X1  g511(.A(G15gat), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(G1326gat));
  NOR2_X1   g513(.A1(new_n694), .A2(new_n484), .ZN(new_n715));
  XOR2_X1   g514(.A(KEYINPUT43), .B(G22gat), .Z(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1327gat));
  AND2_X1   g516(.A1(new_n642), .A2(new_n646), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n691), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n590), .A2(KEYINPUT110), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n588), .A2(new_n721), .A3(new_n589), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n719), .A2(new_n724), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n538), .A2(KEYINPUT44), .A3(new_n673), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n535), .A2(new_n536), .A3(new_n403), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n439), .A2(new_n313), .A3(new_n448), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n416), .A2(new_n421), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n484), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n489), .B(new_n528), .C1(new_n727), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n532), .A2(new_n537), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n673), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n416), .B(new_n725), .C1(new_n726), .C2(new_n735), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n736), .A2(KEYINPUT111), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(KEYINPUT111), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(new_n548), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n731), .A2(new_n732), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n719), .A2(new_n673), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n590), .A3(new_n741), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n742), .A2(new_n415), .A3(new_n548), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT45), .Z(new_n744));
  NAND2_X1  g543(.A1(new_n739), .A2(new_n744), .ZN(G1328gat));
  NOR3_X1   g544(.A1(new_n742), .A2(G36gat), .A3(new_n705), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT46), .ZN(new_n747));
  INV_X1    g546(.A(G36gat), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n538), .B2(new_n673), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n751), .A2(new_n697), .A3(new_n725), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n747), .B1(new_n748), .B2(new_n752), .ZN(G1329gat));
  NAND4_X1  g552(.A1(new_n751), .A2(G43gat), .A3(new_n710), .A4(new_n725), .ZN(new_n754));
  INV_X1    g553(.A(new_n712), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n742), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(G43gat), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT47), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n754), .B(new_n759), .C1(G43gat), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1330gat));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n751), .A2(G50gat), .A3(new_n488), .A4(new_n725), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n544), .B1(new_n742), .B2(new_n484), .ZN(new_n764));
  AOI211_X1 g563(.A(new_n762), .B(KEYINPUT48), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  OR2_X1    g564(.A1(new_n762), .A2(KEYINPUT48), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n762), .A2(KEYINPUT48), .ZN(new_n767));
  AND4_X1   g566(.A1(new_n766), .A2(new_n763), .A3(new_n767), .A4(new_n764), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n765), .A2(new_n768), .ZN(G1331gat));
  NOR2_X1   g568(.A1(new_n674), .A2(new_n723), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n740), .A2(new_n692), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n415), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n607), .ZN(G1332gat));
  NAND2_X1  g572(.A1(new_n771), .A2(KEYINPUT113), .ZN(new_n774));
  INV_X1    g573(.A(new_n770), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n731), .B2(new_n732), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n692), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n705), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n783));
  OAI22_X1  g582(.A1(new_n782), .A2(new_n783), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n779), .A2(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT114), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(G1333gat));
  INV_X1    g589(.A(KEYINPUT50), .ZN(new_n791));
  INV_X1    g590(.A(new_n778), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n777), .B1(new_n776), .B2(new_n692), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n710), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G71gat), .ZN(new_n795));
  INV_X1    g594(.A(G71gat), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n776), .A2(new_n796), .A3(new_n712), .A4(new_n692), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n791), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n528), .B1(new_n774), .B2(new_n778), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n791), .B(new_n797), .C1(new_n799), .C2(new_n796), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(G1334gat));
  NAND2_X1  g601(.A1(new_n779), .A2(new_n488), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g603(.A1(new_n718), .A2(new_n724), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT115), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n692), .B(new_n806), .C1(new_n726), .C2(new_n735), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(new_n415), .A3(new_n648), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n733), .A2(new_n806), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n806), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n691), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n416), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n808), .B1(new_n648), .B2(new_n814), .ZN(G1336gat));
  NAND4_X1  g614(.A1(new_n751), .A2(new_n697), .A3(new_n692), .A4(new_n806), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n705), .A2(G92gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n813), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n673), .ZN(new_n822));
  AND4_X1   g621(.A1(KEYINPUT51), .A2(new_n740), .A3(new_n822), .A4(new_n806), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT51), .B1(new_n733), .B2(new_n806), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT116), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n705), .A2(G92gat), .A3(new_n691), .ZN(new_n829));
  AOI22_X1  g628(.A1(new_n828), .A2(new_n829), .B1(G92gat), .B2(new_n816), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n821), .B1(new_n830), .B2(new_n818), .ZN(G1337gat));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n807), .B2(new_n528), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n691), .B1(new_n749), .B2(new_n750), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(KEYINPUT117), .A3(new_n710), .A4(new_n806), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(G99gat), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(new_n813), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n755), .A2(G99gat), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(G1338gat));
  NAND4_X1  g638(.A1(new_n751), .A2(new_n488), .A3(new_n692), .A4(new_n806), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(G106gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n811), .A2(new_n812), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n484), .A2(G106gat), .A3(new_n691), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT53), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n828), .A2(new_n843), .B1(G106gat), .B2(new_n840), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(G1339gat));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n688), .B1(new_n682), .B2(new_n849), .ZN(new_n850));
  AND3_X1   g649(.A1(new_n680), .A2(new_n681), .A3(new_n676), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n680), .A2(new_n681), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n675), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n680), .A2(new_n681), .A3(new_n676), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT54), .B1(new_n856), .B2(KEYINPUT118), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n850), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n689), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g659(.A(KEYINPUT55), .B(new_n850), .C1(new_n855), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT119), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n856), .B1(new_n682), .B2(KEYINPUT118), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n863), .B(KEYINPUT54), .C1(KEYINPUT118), .C2(new_n856), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT55), .A4(new_n850), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n860), .A2(new_n723), .A3(new_n862), .A4(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n576), .A2(new_n577), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n585), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n589), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n692), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n822), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n860), .A2(new_n862), .A3(new_n866), .A4(new_n871), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n673), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n718), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n770), .A2(new_n691), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n878), .A2(new_n416), .A3(new_n484), .A4(new_n705), .ZN(new_n879));
  INV_X1    g678(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n712), .ZN(new_n881));
  OAI21_X1  g680(.A(G113gat), .B1(new_n881), .B2(new_n591), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n530), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n883), .A2(G113gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n724), .ZN(G1340gat));
  OAI21_X1  g684(.A(G120gat), .B1(new_n881), .B2(new_n691), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n883), .A2(G120gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n691), .ZN(G1341gat));
  INV_X1    g687(.A(G127gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n881), .A2(new_n889), .A3(new_n718), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT120), .B1(new_n883), .B2(new_n718), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT120), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n880), .A2(new_n892), .A3(new_n530), .A4(new_n647), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n894), .B2(new_n889), .ZN(G1342gat));
  INV_X1    g694(.A(G134gat), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n896), .A3(new_n530), .A4(new_n822), .ZN(new_n897));
  OR3_X1    g696(.A1(new_n897), .A2(KEYINPUT121), .A3(KEYINPUT56), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT121), .B1(new_n897), .B2(KEYINPUT56), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n712), .A3(new_n822), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT56), .B1(new_n900), .B2(G134gat), .ZN(new_n901));
  INV_X1    g700(.A(new_n897), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n898), .B(new_n899), .C1(new_n901), .C2(new_n902), .ZN(G1343gat));
  NOR3_X1   g702(.A1(new_n710), .A2(new_n697), .A3(new_n415), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n878), .B2(new_n488), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT57), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n860), .A2(new_n862), .A3(new_n590), .A4(new_n866), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n822), .B1(new_n907), .B2(new_n872), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n718), .B1(new_n908), .B2(new_n875), .ZN(new_n909));
  AOI211_X1 g708(.A(new_n906), .B(new_n484), .C1(new_n909), .C2(new_n877), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n904), .B1(new_n905), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G141gat), .B1(new_n911), .B2(new_n591), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n878), .A2(new_n488), .ZN(new_n914));
  INV_X1    g713(.A(new_n904), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n323), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n912), .B(new_n913), .C1(new_n591), .C2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n917), .A2(new_n591), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n723), .B(new_n904), .C1(new_n905), .C2(new_n910), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(G141gat), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n918), .B1(new_n921), .B2(new_n913), .ZN(G1344gat));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n872), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n673), .ZN(new_n924));
  INV_X1    g723(.A(new_n875), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n647), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n674), .A2(new_n590), .A3(new_n692), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n906), .B(new_n488), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n484), .B1(new_n876), .B2(new_n877), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n928), .B(new_n692), .C1(new_n906), .C2(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(G148gat), .B1(new_n930), .B2(new_n915), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT59), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n692), .B(new_n904), .C1(new_n905), .C2(new_n910), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n325), .A2(KEYINPUT59), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n916), .A2(new_n325), .A3(new_n692), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1345gat));
  NAND2_X1  g739(.A1(new_n647), .A2(G155gat), .ZN(new_n941));
  NOR3_X1   g740(.A1(new_n914), .A2(new_n718), .A3(new_n915), .ZN(new_n942));
  OAI22_X1  g741(.A1(new_n911), .A2(new_n941), .B1(new_n942), .B2(G155gat), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT123), .ZN(G1346gat));
  NAND2_X1  g743(.A1(new_n822), .A2(G162gat), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n914), .A2(new_n673), .A3(new_n915), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n911), .A2(new_n945), .B1(new_n946), .B2(G162gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT124), .ZN(G1347gat));
  AOI21_X1  g747(.A(new_n488), .B1(new_n876), .B2(new_n877), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n697), .A2(new_n415), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n952), .A2(new_n755), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n590), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G169gat), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n949), .A2(new_n530), .A3(new_n951), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n956), .A2(G169gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n724), .B2(new_n957), .ZN(G1348gat));
  INV_X1    g757(.A(new_n956), .ZN(new_n959));
  AOI21_X1  g758(.A(G176gat), .B1(new_n959), .B2(new_n692), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n952), .A2(new_n755), .A3(new_n691), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(G176gat), .B2(new_n961), .ZN(G1349gat));
  AND2_X1   g761(.A1(new_n647), .A2(new_n283), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n949), .A2(new_n712), .A3(new_n647), .A4(new_n951), .ZN(new_n964));
  AOI22_X1  g763(.A1(new_n959), .A2(new_n963), .B1(new_n964), .B2(G183gat), .ZN(new_n965));
  XNOR2_X1  g764(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n965), .B(new_n966), .ZN(G1350gat));
  NAND3_X1  g766(.A1(new_n959), .A2(new_n269), .A3(new_n822), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT61), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n822), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(G190gat), .ZN(new_n971));
  AOI211_X1 g770(.A(KEYINPUT61), .B(new_n269), .C1(new_n953), .C2(new_n822), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1351gat));
  NAND2_X1  g772(.A1(new_n914), .A2(KEYINPUT57), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n950), .A2(new_n710), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n974), .A2(new_n928), .A3(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n977), .A2(KEYINPUT126), .A3(new_n590), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n979), .B1(new_n976), .B2(new_n591), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n978), .A2(G197gat), .A3(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(new_n975), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n914), .A2(new_n982), .ZN(new_n983));
  INV_X1    g782(.A(G197gat), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n983), .A2(new_n984), .A3(new_n723), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n981), .A2(new_n985), .ZN(G1352gat));
  NOR4_X1   g785(.A1(new_n914), .A2(G204gat), .A3(new_n691), .A4(new_n982), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT62), .ZN(new_n988));
  OAI21_X1  g787(.A(G204gat), .B1(new_n930), .B2(new_n982), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(G1353gat));
  INV_X1    g789(.A(G211gat), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n983), .A2(new_n991), .A3(new_n647), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n974), .A2(new_n647), .A3(new_n928), .A4(new_n975), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n983), .B2(new_n822), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n822), .A2(G218gat), .ZN(new_n998));
  XOR2_X1   g797(.A(new_n998), .B(KEYINPUT127), .Z(new_n999));
  AOI21_X1  g798(.A(new_n997), .B1(new_n977), .B2(new_n999), .ZN(G1355gat));
endmodule


