//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT78), .ZN(new_n203));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  NOR3_X1   g009(.A1(new_n210), .A2(KEYINPUT26), .A3(new_n205), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT68), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT27), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT27), .ZN(new_n219));
  AOI21_X1  g018(.A(G190gat), .B1(new_n219), .B2(G183gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT28), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n224), .A3(new_n220), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n220), .A2(KEYINPUT28), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n213), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(KEYINPUT67), .B(G176gat), .ZN(new_n232));
  INV_X1    g031(.A(G169gat), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n233), .A2(KEYINPUT23), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n209), .A2(KEYINPUT23), .ZN(new_n235));
  AOI22_X1  g034(.A1(new_n232), .A2(new_n234), .B1(new_n206), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n204), .A2(KEYINPUT24), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G183gat), .A3(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n241));
  OR3_X1    g040(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n231), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G190gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n215), .A2(new_n217), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n240), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT69), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n240), .A3(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(G176gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n206), .A2(new_n235), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT25), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n244), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n203), .B1(new_n229), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n225), .A2(new_n223), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n224), .B1(new_n218), .B2(new_n220), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n228), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n212), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n246), .A2(new_n240), .A3(new_n249), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n249), .B1(new_n246), .B2(new_n240), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n236), .A2(new_n243), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n230), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n261), .A2(KEYINPUT78), .A3(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(KEYINPUT79), .B(KEYINPUT29), .Z(new_n269));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n257), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT22), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT76), .B(G218gat), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT77), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n276), .A2(new_n279), .A3(new_n277), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n279), .B1(new_n276), .B2(new_n277), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT77), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n270), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n261), .A2(new_n288), .A3(new_n267), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n272), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT37), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n261), .A2(KEYINPUT78), .A3(new_n267), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT78), .B1(new_n261), .B2(new_n267), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI211_X1 g093(.A(KEYINPUT29), .B(new_n288), .C1(new_n261), .C2(new_n267), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n287), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT80), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n270), .B1(new_n257), .B2(new_n268), .ZN(new_n300));
  OAI211_X1 g099(.A(KEYINPUT80), .B(new_n298), .C1(new_n300), .C2(new_n295), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n291), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT37), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(new_n297), .B2(new_n287), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n272), .A2(new_n298), .A3(new_n289), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT38), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G8gat), .B(G36gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(G64gat), .B(G92gat), .ZN(new_n309));
  XOR2_X1   g108(.A(new_n308), .B(new_n309), .Z(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND4_X1  g110(.A1(new_n303), .A2(new_n307), .A3(KEYINPUT90), .A4(new_n311), .ZN(new_n312));
  OR2_X1    g111(.A1(G113gat), .A2(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(G113gat), .A2(G120gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n313), .A2(KEYINPUT71), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT71), .ZN(new_n316));
  AND2_X1   g115(.A1(G113gat), .A2(G120gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(G113gat), .A2(G120gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  XNOR2_X1  g119(.A(G127gat), .B(G134gat), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n315), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT72), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G134gat), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n326), .A2(new_n328), .A3(new_n320), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n319), .A4(new_n315), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT82), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G155gat), .ZN(new_n335));
  INV_X1    g134(.A(G162gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT82), .ZN(new_n338));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n334), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(KEYINPUT2), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT83), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n332), .A2(new_n333), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT2), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n344), .A2(new_n347), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT1), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n352), .A2(new_n321), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n331), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n317), .A2(new_n318), .A3(new_n316), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n328), .A3(new_n320), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT72), .B1(new_n360), .B2(new_n319), .ZN(new_n361));
  INV_X1    g160(.A(new_n330), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n354), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n350), .A2(new_n348), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n345), .B(KEYINPUT83), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n334), .A2(new_n340), .A3(new_n343), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT3), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n364), .B(new_n369), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n363), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n353), .B1(new_n324), .B2(new_n330), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(KEYINPUT4), .A3(new_n351), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n357), .A2(new_n371), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n363), .A2(new_n367), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n372), .B1(new_n377), .B2(new_n355), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n375), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n380), .B(KEYINPUT0), .ZN(new_n381));
  XOR2_X1   g180(.A(G57gat), .B(G85gat), .Z(new_n382));
  XNOR2_X1  g181(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AND4_X1   g183(.A1(KEYINPUT4), .A2(new_n331), .A3(new_n351), .A4(new_n354), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT4), .B1(new_n373), .B2(new_n351), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n387), .A2(KEYINPUT5), .A3(new_n372), .A4(new_n371), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n379), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n384), .B1(new_n379), .B2(new_n388), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT6), .ZN(new_n391));
  AND4_X1   g190(.A1(KEYINPUT6), .A2(new_n379), .A3(new_n384), .A4(new_n388), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT80), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n257), .A2(new_n268), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n295), .B1(new_n395), .B2(new_n288), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n394), .B1(new_n396), .B2(new_n287), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n301), .ZN(new_n398));
  INV_X1    g197(.A(new_n290), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n310), .A3(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n312), .A2(new_n393), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n310), .B1(new_n398), .B2(new_n291), .ZN(new_n402));
  AOI21_X1  g201(.A(KEYINPUT90), .B1(new_n402), .B2(new_n307), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n202), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  OR3_X1    g203(.A1(new_n389), .A2(new_n390), .A3(KEYINPUT6), .ZN(new_n405));
  INV_X1    g204(.A(new_n392), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n405), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n303), .A2(new_n307), .A3(new_n311), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n407), .A2(new_n410), .A3(KEYINPUT91), .A4(new_n312), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT81), .B1(new_n398), .B2(new_n399), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n413));
  AOI211_X1 g212(.A(new_n413), .B(new_n290), .C1(new_n397), .C2(new_n301), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n412), .A2(new_n414), .A3(new_n304), .ZN(new_n415));
  INV_X1    g214(.A(new_n402), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT38), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n404), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  INV_X1    g218(.A(new_n283), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n269), .B1(new_n420), .B2(new_n285), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n351), .B1(new_n421), .B2(new_n369), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n284), .A2(new_n286), .B1(new_n370), .B2(new_n269), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  OR2_X1    g223(.A1(new_n423), .A2(new_n419), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n284), .A2(new_n426), .A3(new_n286), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n351), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(G22gat), .ZN(new_n431));
  INV_X1    g230(.A(G22gat), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n424), .B(new_n432), .C1(new_n425), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT87), .B1(new_n430), .B2(G22gat), .ZN(new_n435));
  XOR2_X1   g234(.A(G78gat), .B(G106gat), .Z(new_n436));
  XNOR2_X1  g235(.A(KEYINPUT86), .B(G50gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(KEYINPUT85), .B(KEYINPUT31), .Z(new_n439));
  XOR2_X1   g238(.A(new_n438), .B(new_n439), .Z(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n434), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n431), .A2(KEYINPUT87), .A3(new_n433), .A4(new_n440), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n399), .B1(new_n299), .B2(new_n302), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(new_n413), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n290), .B1(new_n397), .B2(new_n301), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT81), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n449), .A3(new_n311), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT30), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n400), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(KEYINPUT30), .A3(new_n310), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n372), .B1(new_n387), .B2(new_n371), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT39), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n384), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n377), .A2(new_n372), .A3(new_n355), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT39), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n457), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT40), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n462), .B1(new_n460), .B2(new_n461), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n463), .A2(new_n464), .A3(new_n389), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n445), .B1(new_n454), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n418), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n468), .A2(KEYINPUT75), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n471), .A2(KEYINPUT36), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n373), .B1(new_n229), .B2(new_n256), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n261), .A2(new_n363), .A3(new_n267), .ZN(new_n475));
  INV_X1    g274(.A(G227gat), .ZN(new_n476));
  INV_X1    g275(.A(G233gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(new_n478), .B(KEYINPUT64), .Z(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n480), .A2(KEYINPUT32), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G43gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G71gat), .B(G99gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(KEYINPUT33), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n486), .A2(KEYINPUT73), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n481), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n474), .A2(new_n475), .A3(new_n479), .A4(new_n485), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT73), .B1(new_n489), .B2(new_n486), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n488), .B1(new_n490), .B2(new_n481), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n475), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n479), .A2(KEYINPUT34), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n478), .B1(new_n474), .B2(new_n475), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n494), .B(KEYINPUT74), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT74), .ZN(new_n498));
  INV_X1    g297(.A(new_n494), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n496), .A2(new_n495), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n491), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n490), .A2(new_n481), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n499), .A2(new_n500), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT74), .A4(new_n488), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n470), .B(new_n473), .C1(new_n503), .C2(new_n507), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n502), .A2(new_n506), .A3(new_n471), .A4(KEYINPUT36), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n393), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n450), .A2(new_n511), .A3(new_n452), .A4(new_n453), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n442), .A2(KEYINPUT88), .A3(new_n443), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT88), .B1(new_n442), .B2(new_n443), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n510), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n452), .A2(new_n453), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n506), .A2(new_n502), .B1(new_n442), .B2(new_n443), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n517), .A2(new_n511), .A3(new_n450), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n520));
  INV_X1    g319(.A(new_n518), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n454), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT35), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n523), .A3(new_n511), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n467), .A2(new_n516), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n526), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT93), .B(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT14), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  NAND2_X1  g338(.A1(G43gat), .A2(G50gat), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT96), .B(G50gat), .Z(new_n541));
  OAI211_X1 g340(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(G43gat), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(G43gat), .A2(G50gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n539), .B1(new_n544), .B2(new_n540), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(KEYINPUT95), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  INV_X1    g347(.A(new_n545), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n538), .B2(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT94), .B(new_n545), .C1(new_n535), .C2(new_n537), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n547), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n532), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n543), .A2(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT17), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(G229gat), .A2(G233gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n553), .A2(new_n532), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n558), .A2(KEYINPUT18), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT97), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n555), .A2(new_n557), .B1(new_n553), .B2(new_n532), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n564), .A2(KEYINPUT97), .A3(KEYINPUT18), .A4(new_n559), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n559), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n556), .A2(new_n531), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n559), .B(KEYINPUT13), .Z(new_n571));
  AOI22_X1  g370(.A1(new_n567), .A2(new_n568), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n577), .B(KEYINPUT12), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n566), .A2(new_n572), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n579), .B1(new_n566), .B2(new_n572), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n525), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n553), .A2(new_n554), .ZN(new_n585));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT7), .ZN(new_n587));
  INV_X1    g386(.A(G99gat), .ZN(new_n588));
  INV_X1    g387(.A(G106gat), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT8), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT101), .B(G92gat), .Z(new_n591));
  OAI211_X1 g390(.A(new_n587), .B(new_n590), .C1(G85gat), .C2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n585), .A2(new_n557), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n593), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n592), .B(new_n596), .ZN(new_n597));
  AND2_X1   g396(.A1(G232gat), .A2(G233gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n553), .A2(new_n597), .B1(KEYINPUT41), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT102), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G134gat), .B(G162gat), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n601), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n598), .A2(KEYINPUT41), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  OR3_X1    g409(.A1(new_n605), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n610), .B1(new_n605), .B2(new_n606), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G57gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(G64gat), .ZN(new_n615));
  INV_X1    g414(.A(G64gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G57gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT98), .B2(KEYINPUT9), .ZN(new_n619));
  INV_X1    g418(.A(G71gat), .ZN(new_n620));
  INV_X1    g419(.A(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR3_X1    g421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT98), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT98), .B1(new_n620), .B2(new_n621), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT9), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n620), .B2(new_n621), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n615), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n617), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n625), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT21), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(G231gat), .A2(G233gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(new_n327), .ZN(new_n638));
  XNOR2_X1  g437(.A(G183gat), .B(G211gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n531), .B1(new_n634), .B2(new_n633), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT100), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n335), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n640), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT10), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n594), .A2(new_n647), .A3(new_n633), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT103), .ZN(new_n649));
  INV_X1    g448(.A(new_n633), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n649), .B1(new_n597), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n594), .A2(KEYINPUT103), .A3(new_n633), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT104), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n592), .A2(new_n653), .A3(new_n593), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n593), .B1(new_n592), .B2(new_n653), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n633), .ZN(new_n656));
  AOI22_X1  g455(.A1(new_n651), .A2(new_n652), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n648), .B1(new_n657), .B2(new_n647), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT105), .Z(new_n660));
  OR2_X1    g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n657), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  XOR2_X1   g463(.A(G120gat), .B(G148gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT106), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n661), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n670));
  INV_X1    g469(.A(new_n668), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n658), .A2(new_n660), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n671), .B1(new_n672), .B2(new_n663), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  OAI211_X1 g473(.A(KEYINPUT107), .B(new_n671), .C1(new_n672), .C2(new_n663), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n613), .A2(new_n646), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n584), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n511), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(G1gat), .Z(G1324gat));
  NAND2_X1  g480(.A1(new_n584), .A2(new_n454), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n677), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT16), .B(G8gat), .Z(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n685), .B1(new_n530), .B2(new_n683), .ZN(new_n686));
  MUX2_X1   g485(.A(new_n685), .B(new_n686), .S(KEYINPUT42), .Z(G1325gat));
  AOI211_X1 g486(.A(new_n469), .B(new_n472), .C1(new_n502), .C2(new_n506), .ZN(new_n688));
  INV_X1    g487(.A(new_n509), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G15gat), .B1(new_n679), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n503), .A2(new_n507), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n584), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n677), .A2(G15gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g495(.A1(new_n584), .A2(new_n515), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n677), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT43), .B(G22gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n613), .ZN(new_n701));
  INV_X1    g500(.A(new_n646), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n676), .ZN(new_n703));
  INV_X1    g502(.A(new_n533), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(new_n511), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n584), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n525), .B2(new_n613), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n646), .B(KEYINPUT108), .ZN(new_n710));
  INV_X1    g509(.A(new_n582), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n580), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n710), .A2(new_n712), .A3(new_n676), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT109), .Z(new_n714));
  NAND2_X1  g513(.A1(new_n512), .A2(new_n515), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n690), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n418), .B2(new_n466), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n519), .B(new_n523), .ZN(new_n718));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n701), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n709), .A2(new_n714), .A3(new_n393), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n704), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n707), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT110), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1328gat));
  NOR3_X1   g523(.A1(new_n682), .A2(G36gat), .A3(new_n703), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT46), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n709), .A2(new_n719), .ZN(new_n727));
  AND3_X1   g526(.A1(new_n727), .A2(new_n454), .A3(new_n714), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n534), .B2(new_n728), .ZN(G1329gat));
  NAND3_X1  g528(.A1(new_n727), .A2(new_n510), .A3(new_n714), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G43gat), .ZN(new_n731));
  OR3_X1    g530(.A1(new_n694), .A2(G43gat), .A3(new_n703), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1330gat));
  NAND3_X1  g535(.A1(new_n727), .A2(new_n445), .A3(new_n714), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n737), .A2(new_n541), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n697), .A2(new_n541), .A3(new_n703), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n727), .A2(new_n515), .A3(new_n714), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(new_n541), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n738), .A2(new_n741), .B1(new_n743), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n467), .A2(new_n516), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n524), .A2(new_n520), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n676), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n701), .A2(new_n702), .A3(new_n712), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(new_n511), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n614), .ZN(G1332gat));
  XNOR2_X1  g551(.A(new_n750), .B(KEYINPUT112), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n753), .A2(new_n454), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NAND3_X1  g557(.A1(new_n753), .A2(G71gat), .A3(new_n510), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n620), .B1(new_n750), .B2(new_n692), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(KEYINPUT50), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT50), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n761), .A2(new_n762), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n753), .A2(new_n515), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G78gat), .ZN(G1335gat));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n525), .B2(new_n613), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n712), .A2(new_n646), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT114), .B(new_n701), .C1(new_n717), .C2(new_n718), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n767), .A2(KEYINPUT51), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT115), .ZN(new_n771));
  INV_X1    g570(.A(new_n768), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n613), .B1(new_n745), .B2(new_n746), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(KEYINPUT114), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n774), .A2(new_n775), .A3(KEYINPUT51), .A4(new_n767), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n768), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT114), .B1(new_n747), .B2(new_n701), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n771), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n676), .A2(new_n511), .A3(G85gat), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT116), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n772), .A2(new_n676), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n709), .A2(new_n719), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n709), .A2(KEYINPUT113), .A3(new_n719), .A4(new_n785), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n393), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G85gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n784), .A2(new_n791), .ZN(G1336gat));
  INV_X1    g591(.A(new_n454), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n793), .A2(G92gat), .A3(new_n676), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n781), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n591), .B1(new_n786), .B2(new_n793), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n788), .A2(new_n454), .A3(new_n789), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n780), .A2(new_n770), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n799), .A2(new_n591), .B1(new_n800), .B2(new_n794), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n795), .A2(new_n798), .B1(new_n801), .B2(new_n802), .ZN(G1337gat));
  NAND4_X1  g602(.A1(new_n781), .A2(new_n588), .A3(new_n693), .A4(new_n748), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n788), .A2(new_n510), .A3(new_n789), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n588), .B2(new_n805), .ZN(G1338gat));
  NOR3_X1   g605(.A1(new_n676), .A2(G106gat), .A3(new_n444), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n781), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g607(.A(KEYINPUT118), .B(G106gat), .Z(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n786), .B2(new_n444), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n788), .A2(new_n515), .A3(new_n789), .ZN(new_n813));
  AOI22_X1  g612(.A1(new_n813), .A2(new_n809), .B1(new_n800), .B2(new_n807), .ZN(new_n814));
  OAI22_X1  g613(.A1(new_n808), .A2(new_n812), .B1(new_n814), .B2(new_n811), .ZN(G1339gat));
  NOR2_X1   g614(.A1(new_n677), .A2(new_n712), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n658), .A2(new_n660), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n661), .A2(KEYINPUT54), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n668), .B1(new_n672), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n819), .A2(KEYINPUT55), .A3(new_n821), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n669), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n564), .A2(new_n559), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n570), .A2(new_n571), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n577), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n580), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n826), .A2(new_n613), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n674), .A2(new_n580), .A3(new_n675), .A4(new_n829), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n826), .B2(new_n583), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n831), .B1(new_n613), .B2(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n646), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n817), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  AND3_X1   g636(.A1(new_n837), .A2(new_n393), .A3(new_n522), .ZN(new_n838));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838), .B2(new_n712), .ZN(new_n839));
  INV_X1    g638(.A(new_n515), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT119), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n837), .A2(KEYINPUT119), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n793), .A2(new_n393), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n692), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n712), .A2(G113gat), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n839), .B1(new_n847), .B2(new_n848), .ZN(G1340gat));
  AOI21_X1  g648(.A(G120gat), .B1(new_n838), .B2(new_n748), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n748), .A2(G120gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n847), .B2(new_n851), .ZN(G1341gat));
  NAND3_X1  g651(.A1(new_n838), .A2(new_n327), .A3(new_n646), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n847), .A2(new_n836), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(new_n327), .ZN(G1342gat));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n325), .A3(new_n701), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n844), .A2(new_n701), .A3(new_n846), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n859), .A2(KEYINPUT120), .A3(G134gat), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT120), .B1(new_n859), .B2(G134gat), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n857), .B(new_n858), .C1(new_n860), .C2(new_n861), .ZN(G1343gat));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n833), .A2(new_n613), .ZN(new_n864));
  OR3_X1    g663(.A1(new_n826), .A2(new_n613), .A3(new_n830), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n836), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g665(.A(new_n863), .B(new_n445), .C1(new_n866), .C2(new_n816), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n845), .A2(new_n510), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n822), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n819), .A2(KEYINPUT121), .A3(new_n821), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n823), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n825), .A2(new_n669), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n712), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n701), .B1(new_n875), .B2(new_n832), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n702), .B1(new_n876), .B2(new_n831), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n840), .B1(new_n877), .B2(new_n817), .ZN(new_n878));
  OAI211_X1 g677(.A(new_n867), .B(new_n868), .C1(new_n878), .C2(new_n863), .ZN(new_n879));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879), .B2(new_n583), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n510), .A2(new_n444), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n393), .A2(new_n837), .A3(new_n793), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n583), .A2(G141gat), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT58), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n832), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n583), .A2(new_n873), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(new_n872), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n865), .B1(new_n890), .B2(new_n701), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n816), .B1(new_n891), .B2(new_n702), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n840), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n893), .A2(KEYINPUT122), .A3(new_n867), .A4(new_n868), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n894), .A3(new_n712), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n895), .A2(G141gat), .B1(new_n882), .B2(new_n883), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n885), .B1(new_n896), .B2(new_n897), .ZN(G1344gat));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n899), .B(G148gat), .C1(new_n882), .C2(new_n748), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n887), .A2(new_n894), .A3(new_n748), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n899), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n863), .B1(new_n837), .B2(new_n445), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n863), .B2(new_n878), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(KEYINPUT59), .A3(new_n748), .A4(new_n868), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n900), .B1(new_n906), .B2(G148gat), .ZN(G1345gat));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n894), .ZN(new_n908));
  OAI21_X1  g707(.A(G155gat), .B1(new_n908), .B2(new_n710), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n882), .A2(new_n335), .A3(new_n646), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1346gat));
  NAND3_X1  g710(.A1(new_n882), .A2(new_n336), .A3(new_n701), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT123), .Z(new_n913));
  OAI21_X1  g712(.A(G162gat), .B1(new_n908), .B2(new_n613), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n866), .A2(new_n816), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(new_n393), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n793), .A2(new_n521), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(KEYINPUT124), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n712), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n793), .A2(new_n393), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n692), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n842), .B2(new_n843), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n583), .A2(new_n233), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n922), .A2(new_n233), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  NAND3_X1  g728(.A1(new_n920), .A2(new_n748), .A3(new_n921), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n676), .A2(new_n232), .ZN(new_n931));
  AOI22_X1  g730(.A1(new_n930), .A2(new_n252), .B1(new_n927), .B2(new_n931), .ZN(G1349gat));
  INV_X1    g731(.A(new_n919), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n219), .A2(G183gat), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n933), .A2(new_n934), .A3(new_n227), .A4(new_n646), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n927), .A2(new_n836), .B1(new_n215), .B2(new_n217), .ZN(new_n937));
  OAI21_X1  g736(.A(KEYINPUT60), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n927), .A2(new_n836), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n215), .A2(new_n217), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT60), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n941), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n938), .A2(new_n943), .ZN(G1350gat));
  INV_X1    g743(.A(new_n843), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n701), .B(new_n925), .C1(new_n945), .C2(new_n841), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(G190gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n946), .A2(new_n949), .A3(G190gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n948), .A2(KEYINPUT61), .A3(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(KEYINPUT125), .A3(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n920), .A2(new_n245), .A3(new_n701), .A4(new_n921), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n953), .A3(new_n954), .ZN(G1351gat));
  NOR2_X1   g754(.A1(new_n924), .A2(new_n510), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n904), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n957), .A2(new_n958), .A3(new_n583), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n917), .A2(new_n454), .A3(new_n881), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n960), .A2(new_n583), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n959), .B1(new_n958), .B2(new_n961), .ZN(G1352gat));
  NOR3_X1   g761(.A1(new_n793), .A2(G204gat), .A3(new_n676), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n917), .A2(new_n881), .A3(new_n963), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(KEYINPUT62), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n967));
  XOR2_X1   g766(.A(new_n966), .B(new_n967), .Z(new_n968));
  OAI21_X1  g767(.A(G204gat), .B1(new_n957), .B2(new_n676), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n968), .A2(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n904), .A2(new_n646), .A3(new_n956), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n971), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT63), .B1(new_n971), .B2(G211gat), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n646), .A2(new_n275), .ZN(new_n974));
  OAI22_X1  g773(.A1(new_n972), .A2(new_n973), .B1(new_n960), .B2(new_n974), .ZN(G1354gat));
  INV_X1    g774(.A(new_n957), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n613), .A2(new_n274), .ZN(new_n977));
  XOR2_X1   g776(.A(new_n977), .B(KEYINPUT127), .Z(new_n978));
  OR2_X1    g777(.A1(new_n960), .A2(new_n613), .ZN(new_n979));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  AOI22_X1  g779(.A1(new_n976), .A2(new_n978), .B1(new_n979), .B2(new_n980), .ZN(G1355gat));
endmodule


