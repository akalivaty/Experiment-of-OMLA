//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT74), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n203), .A2(new_n204), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G211gat), .B(G218gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT76), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT29), .ZN(new_n213));
  XOR2_X1   g012(.A(G155gat), .B(G162gat), .Z(new_n214));
  XOR2_X1   g013(.A(G141gat), .B(G148gat), .Z(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(KEYINPUT81), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT2), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n219), .B(new_n215), .C1(new_n214), .C2(KEYINPUT81), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XOR2_X1   g023(.A(KEYINPUT82), .B(KEYINPUT3), .Z(new_n225));
  OAI21_X1  g024(.A(new_n213), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n212), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n207), .A2(new_n210), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT29), .B1(new_n207), .B2(new_n210), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n225), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G228gat), .ZN(new_n232));
  INV_X1    g031(.A(G233gat), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n231), .A2(new_n223), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n211), .A2(new_n213), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n235), .B2(KEYINPUT3), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G228gat), .A2(G233gat), .ZN(new_n238));
  OAI221_X1 g037(.A(G22gat), .B1(new_n228), .B2(new_n234), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  AOI211_X1 g039(.A(new_n232), .B(new_n233), .C1(new_n227), .C2(new_n236), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n228), .A2(new_n234), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G78gat), .B(G106gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT31), .B(G50gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(KEYINPUT84), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n239), .A2(new_n243), .A3(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n239), .A2(new_n243), .B1(KEYINPUT84), .B2(new_n246), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT72), .ZN(new_n251));
  XNOR2_X1  g050(.A(G15gat), .B(G43gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(G71gat), .B(G99gat), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n252), .B(new_n253), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G227gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(new_n233), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(G113gat), .B2(G120gat), .ZN(new_n260));
  AND2_X1   g059(.A1(G113gat), .A2(G120gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT68), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G127gat), .B(G134gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  INV_X1    g066(.A(G183gat), .ZN(new_n268));
  OAI211_X1 g067(.A(KEYINPUT65), .B(new_n267), .C1(new_n268), .C2(KEYINPUT27), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT28), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272));
  AOI21_X1  g071(.A(G190gat), .B1(new_n272), .B2(G183gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n268), .A2(KEYINPUT27), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n266), .B1(new_n271), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT66), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n277), .A2(new_n281), .A3(new_n278), .ZN(new_n282));
  OR2_X1    g081(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n283));
  INV_X1    g082(.A(G169gat), .ZN(new_n284));
  INV_X1    g083(.A(G176gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(KEYINPUT67), .A2(KEYINPUT26), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n283), .A2(new_n284), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n280), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n269), .A2(new_n273), .A3(new_n270), .A4(new_n274), .ZN(new_n289));
  AND3_X1   g088(.A1(new_n276), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT24), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n265), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n268), .A2(new_n267), .ZN(new_n293));
  NAND3_X1  g092(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(G169gat), .B2(G176gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT23), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n295), .A2(new_n297), .A3(new_n278), .A4(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n292), .A2(KEYINPUT64), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n265), .A2(new_n302), .A3(new_n291), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n301), .A2(new_n293), .A3(new_n294), .A4(new_n303), .ZN(new_n304));
  AND4_X1   g103(.A1(KEYINPUT25), .A2(new_n298), .A3(new_n297), .A4(new_n278), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n299), .A2(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI211_X1 g105(.A(new_n258), .B(new_n264), .C1(new_n290), .C2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n264), .ZN(new_n308));
  INV_X1    g107(.A(new_n295), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n298), .A2(new_n297), .A3(new_n278), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n300), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n305), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n276), .A2(new_n288), .A3(new_n289), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n313), .A2(new_n314), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n258), .B1(new_n317), .B2(new_n264), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n257), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n255), .B1(new_n319), .B2(KEYINPUT32), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT71), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT70), .B(KEYINPUT33), .Z(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n319), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n319), .B2(new_n323), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n251), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n326), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n324), .A4(new_n320), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n319), .B(KEYINPUT32), .C1(new_n323), .C2(new_n255), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT73), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT34), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n316), .A2(new_n318), .ZN(new_n337));
  INV_X1    g136(.A(new_n257), .ZN(new_n338));
  AOI22_X1  g137(.A1(new_n337), .A2(new_n338), .B1(new_n333), .B2(new_n334), .ZN(new_n339));
  INV_X1    g138(.A(new_n335), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n330), .A2(new_n340), .A3(new_n331), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n339), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n340), .B1(new_n330), .B2(new_n331), .ZN(new_n344));
  INV_X1    g143(.A(new_n331), .ZN(new_n345));
  AOI211_X1 g144(.A(new_n335), .B(new_n345), .C1(new_n327), .C2(new_n329), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n343), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n250), .B1(new_n342), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n223), .B(new_n264), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT5), .ZN(new_n350));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n223), .A2(new_n308), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(KEYINPUT4), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n357));
  INV_X1    g156(.A(new_n225), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n308), .B1(new_n223), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n351), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(new_n350), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n354), .A2(new_n355), .B1(new_n357), .B2(new_n359), .ZN(new_n365));
  INV_X1    g164(.A(new_n363), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n351), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n352), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  INV_X1    g168(.A(G85gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  NAND3_X1  g172(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n352), .ZN(new_n375));
  INV_X1    g174(.A(new_n367), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n366), .B1(new_n365), .B2(new_n351), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n373), .B(new_n375), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n368), .A2(new_n373), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n374), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n313), .B2(new_n314), .ZN(new_n383));
  AND2_X1   g182(.A1(G226gat), .A2(G233gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n317), .A2(new_n384), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n212), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n385), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n388), .B1(new_n391), .B2(new_n212), .ZN(new_n392));
  XNOR2_X1  g191(.A(G8gat), .B(G36gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(G92gat), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT78), .B(G64gat), .ZN(new_n395));
  XOR2_X1   g194(.A(new_n394), .B(new_n395), .Z(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(KEYINPUT30), .A3(new_n397), .ZN(new_n399));
  XOR2_X1   g198(.A(KEYINPUT79), .B(KEYINPUT30), .Z(new_n400));
  AOI21_X1  g199(.A(new_n400), .B1(new_n392), .B2(new_n397), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n398), .B(new_n399), .C1(new_n401), .C2(KEYINPUT80), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(KEYINPUT80), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n348), .A2(new_n382), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT6), .B1(new_n368), .B2(new_n373), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n407), .B(new_n408), .C1(new_n373), .C2(new_n368), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT86), .B1(new_n380), .B2(new_n381), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n374), .ZN(new_n411));
  XOR2_X1   g210(.A(KEYINPUT87), .B(KEYINPUT35), .Z(new_n412));
  AND3_X1   g211(.A1(new_n411), .A2(new_n405), .A3(new_n412), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n406), .A2(KEYINPUT35), .B1(new_n348), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT36), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n339), .B1(new_n336), .B2(new_n341), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n344), .A2(new_n346), .A3(new_n343), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n342), .A2(new_n347), .A3(KEYINPUT36), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n349), .A2(new_n351), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT39), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n356), .A2(new_n360), .ZN(new_n423));
  INV_X1    g222(.A(new_n351), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n373), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(KEYINPUT40), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  OR3_X1    g229(.A1(new_n365), .A2(KEYINPUT39), .A3(new_n351), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n426), .A2(new_n427), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n432), .A2(new_n378), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n423), .A2(new_n424), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n427), .B1(new_n434), .B2(KEYINPUT39), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n429), .B1(new_n435), .B2(new_n425), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n433), .B(new_n436), .C1(new_n402), .C2(new_n404), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n239), .A2(new_n243), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n246), .A2(KEYINPUT84), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n239), .A2(new_n243), .A3(new_n247), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT37), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n397), .B1(new_n392), .B2(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n443), .B2(new_n392), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT38), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n397), .A2(KEYINPUT38), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n212), .B1(new_n386), .B2(new_n387), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n448), .A2(new_n443), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n391), .A2(new_n212), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n392), .A2(new_n443), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n451), .A2(new_n452), .B1(new_n397), .B2(new_n392), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n437), .B(new_n442), .C1(new_n411), .C2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n401), .A2(KEYINPUT80), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n398), .A2(new_n399), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n382), .A2(new_n403), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n250), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n420), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n414), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G43gat), .B(G50gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT90), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(G29gat), .A2(G36gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT14), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT89), .B(G36gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G29gat), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n465), .A2(new_n468), .A3(KEYINPUT15), .A4(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n470), .ZN(new_n473));
  INV_X1    g272(.A(new_n463), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n464), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n471), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT17), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g278(.A(KEYINPUT17), .B(new_n471), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  XOR2_X1   g280(.A(G15gat), .B(G22gat), .Z(new_n482));
  INV_X1    g281(.A(G1gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n485), .B1(new_n486), .B2(G1gat), .ZN(new_n487));
  INV_X1    g286(.A(G8gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT93), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n489), .A2(new_n490), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT92), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(KEYINPUT91), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n482), .A2(KEYINPUT92), .A3(new_n483), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT91), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n485), .B(new_n497), .C1(new_n486), .C2(G1gat), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n498), .ZN(new_n499));
  AOI22_X1  g298(.A1(new_n491), .A2(new_n492), .B1(new_n499), .B2(G8gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n481), .A2(KEYINPUT94), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n491), .A2(new_n492), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(G8gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n505), .B1(new_n479), .B2(new_n480), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT94), .ZN(new_n507));
  INV_X1    g306(.A(new_n477), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n507), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n501), .B(new_n502), .C1(new_n506), .C2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT18), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n481), .A2(new_n500), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT94), .B1(new_n500), .B2(new_n477), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n515), .A2(KEYINPUT18), .A3(new_n502), .A4(new_n501), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n500), .B(new_n508), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT13), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n512), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n521));
  XNOR2_X1  g320(.A(G113gat), .B(G141gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n525), .B(KEYINPUT12), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n520), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n526), .A3(new_n519), .A4(new_n516), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n462), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G71gat), .A2(G78gat), .ZN(new_n533));
  OR2_X1    g332(.A1(G71gat), .A2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT9), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G64gat), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT95), .B1(new_n537), .B2(G57gat), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G64gat), .ZN(new_n540));
  NOR3_X1   g339(.A1(new_n537), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n537), .A2(G57gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n539), .A2(G64gat), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT9), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n545), .A2(new_n533), .A3(new_n534), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT21), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n500), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT96), .ZN(new_n550));
  AND2_X1   g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n547), .A2(KEYINPUT21), .ZN(new_n553));
  XNOR2_X1  g352(.A(G127gat), .B(G155gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n552), .A2(new_n555), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n561), .A3(new_n557), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  AOI22_X1  g366(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n370), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n569), .B1(new_n370), .B2(new_n567), .ZN(new_n570));
  NAND3_X1  g369(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n572), .B(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n575), .B1(new_n479), .B2(new_n480), .ZN(new_n576));
  XOR2_X1   g375(.A(G190gat), .B(G218gat), .Z(new_n577));
  NAND3_X1  g376(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n572), .B(new_n573), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n578), .B1(new_n477), .B2(new_n579), .ZN(new_n580));
  OR3_X1    g379(.A1(new_n576), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT97), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n577), .B1(new_n576), .B2(new_n580), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n585), .B1(new_n581), .B2(new_n586), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n572), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n547), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n592), .A2(new_n542), .A3(new_n546), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n575), .A2(new_n547), .A3(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(G230gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n600), .A2(new_n233), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n593), .A2(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n601), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G176gat), .B(G204gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(KEYINPUT99), .ZN(new_n608));
  XNOR2_X1  g407(.A(G120gat), .B(G148gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n605), .A3(new_n610), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT100), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT100), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n565), .A2(new_n590), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n532), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(new_n382), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n483), .ZN(G1324gat));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  INV_X1    g423(.A(new_n405), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT16), .B(G8gat), .Z(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(KEYINPUT42), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n625), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n630), .B2(G8gat), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n628), .B1(new_n627), .B2(new_n631), .ZN(G1325gat));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n342), .A2(new_n347), .A3(KEYINPUT36), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT36), .B1(new_n342), .B2(new_n347), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT101), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n418), .A2(new_n637), .A3(new_n419), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n621), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n342), .A2(new_n347), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n633), .B2(new_n642), .ZN(G1326gat));
  NOR2_X1   g442(.A1(new_n621), .A2(new_n442), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT43), .B(G22gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(G1327gat));
  NOR3_X1   g445(.A1(new_n565), .A2(new_n590), .A3(new_n617), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n532), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n382), .A2(G29gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT45), .Z(new_n651));
  INV_X1    g450(.A(new_n590), .ZN(new_n652));
  OAI211_X1 g451(.A(KEYINPUT44), .B(new_n652), .C1(new_n414), .C2(new_n461), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n617), .B(KEYINPUT102), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NOR3_X1   g454(.A1(new_n655), .A2(new_n531), .A3(new_n565), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT103), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n657), .B1(new_n588), .B2(new_n589), .ZN(new_n658));
  INV_X1    g457(.A(new_n589), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n659), .A2(KEYINPUT103), .A3(new_n587), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n455), .A2(new_n459), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n636), .A2(new_n638), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n413), .A2(new_n348), .ZN(new_n665));
  AOI211_X1 g464(.A(new_n250), .B(new_n458), .C1(new_n342), .C2(new_n347), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT35), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n662), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n653), .B(new_n656), .C1(new_n669), .C2(KEYINPUT44), .ZN(new_n670));
  OAI21_X1  g469(.A(G29gat), .B1(new_n670), .B2(new_n382), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n671), .ZN(G1328gat));
  NOR3_X1   g471(.A1(new_n648), .A2(new_n405), .A3(new_n469), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT46), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n469), .B1(new_n670), .B2(new_n405), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(G1329gat));
  OAI21_X1  g475(.A(G43gat), .B1(new_n670), .B2(new_n639), .ZN(new_n677));
  INV_X1    g476(.A(G43gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n641), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n648), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT47), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1330gat));
  NOR2_X1   g481(.A1(new_n648), .A2(new_n442), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n250), .A2(G50gat), .ZN(new_n684));
  OAI22_X1  g483(.A1(new_n683), .A2(G50gat), .B1(new_n670), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g485(.A1(new_n664), .A2(new_n668), .ZN(new_n687));
  INV_X1    g486(.A(new_n565), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n688), .A2(new_n654), .A3(new_n530), .A4(new_n652), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n382), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(new_n539), .ZN(G1332gat));
  INV_X1    g491(.A(new_n690), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n405), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT104), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n696), .B(new_n697), .Z(G1333gat));
  OAI21_X1  g497(.A(G71gat), .B1(new_n690), .B2(new_n639), .ZN(new_n699));
  INV_X1    g498(.A(G71gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n641), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n690), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g502(.A1(new_n693), .A2(new_n250), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n531), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(new_n590), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n687), .A2(KEYINPUT51), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(KEYINPUT51), .B1(new_n687), .B2(new_n707), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n618), .A2(new_n382), .A3(G85gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT105), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n706), .A2(new_n618), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n653), .B(new_n714), .C1(new_n669), .C2(KEYINPUT44), .ZN(new_n715));
  OAI21_X1  g514(.A(G85gat), .B1(new_n715), .B2(new_n382), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1336gat));
  OAI21_X1  g516(.A(G92gat), .B1(new_n715), .B2(new_n405), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n405), .A2(G92gat), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n655), .B(new_n719), .C1(new_n708), .C2(new_n709), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT52), .ZN(G1337gat));
  AOI211_X1 g521(.A(G99gat), .B(new_n618), .C1(new_n342), .C2(new_n347), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT106), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n710), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G99gat), .B1(new_n715), .B2(new_n639), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n725), .A2(KEYINPUT107), .A3(new_n726), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(G1338gat));
  OAI21_X1  g530(.A(G106gat), .B1(new_n715), .B2(new_n442), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(KEYINPUT108), .B(G106gat), .C1(new_n715), .C2(new_n442), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n442), .A2(G106gat), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n655), .B(new_n736), .C1(new_n708), .C2(new_n709), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT53), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT53), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT109), .B1(new_n715), .B2(new_n442), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G106gat), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n715), .A2(KEYINPUT109), .A3(new_n442), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n740), .B(new_n737), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n739), .A2(new_n744), .ZN(G1339gat));
  INV_X1    g544(.A(G113gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n620), .A2(new_n531), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n597), .A2(new_n601), .A3(new_n598), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n603), .A2(KEYINPUT54), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT110), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n603), .A2(new_n752), .A3(KEYINPUT54), .A4(new_n749), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n601), .B1(new_n597), .B2(new_n598), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n610), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n751), .A2(KEYINPUT55), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n613), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n611), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n750), .B2(KEYINPUT110), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT55), .B1(new_n761), .B2(new_n753), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n758), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n530), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n502), .B1(new_n515), .B2(new_n501), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n517), .A2(new_n518), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n525), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n529), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n617), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n661), .B1(new_n764), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n529), .A2(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT112), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n529), .A2(new_n767), .A3(new_n773), .ZN(new_n774));
  AND4_X1   g573(.A1(new_n661), .A2(new_n763), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n748), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n763), .A2(new_n772), .A3(new_n661), .A4(new_n774), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n763), .A2(new_n530), .B1(new_n617), .B2(new_n768), .ZN(new_n778));
  OAI211_X1 g577(.A(KEYINPUT113), .B(new_n777), .C1(new_n778), .C2(new_n661), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n688), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n747), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n625), .A2(new_n382), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n348), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n746), .B1(new_n784), .B2(new_n530), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT114), .Z(new_n786));
  XOR2_X1   g585(.A(new_n784), .B(KEYINPUT115), .Z(new_n787));
  NAND3_X1  g586(.A1(new_n787), .A2(new_n746), .A3(new_n530), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1340gat));
  NOR2_X1   g588(.A1(new_n618), .A2(G120gat), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n790), .B(KEYINPUT116), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n784), .ZN(new_n793));
  OAI21_X1  g592(.A(G120gat), .B1(new_n793), .B2(new_n654), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1341gat));
  NAND2_X1  g594(.A1(new_n784), .A2(new_n565), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT117), .B(G127gat), .Z(new_n797));
  XNOR2_X1  g596(.A(new_n796), .B(new_n797), .ZN(G1342gat));
  NAND2_X1  g597(.A1(new_n784), .A2(new_n652), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(G134gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(KEYINPUT56), .B2(new_n803), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(KEYINPUT56), .B2(new_n803), .ZN(G1343gat));
  AND2_X1   g604(.A1(new_n639), .A2(new_n782), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n778), .A2(new_n652), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n565), .B1(new_n807), .B2(new_n777), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n619), .A2(new_n530), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n250), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT57), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n781), .A2(new_n250), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(KEYINPUT57), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(G141gat), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n531), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n813), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n806), .A2(new_n818), .A3(new_n530), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n815), .A2(new_n817), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT118), .ZN(new_n821));
  OR3_X1    g620(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT58), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT58), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1344gat));
  INV_X1    g623(.A(G148gat), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n806), .A2(new_n818), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n618), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n763), .A2(new_n772), .A3(new_n652), .A4(new_n774), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n807), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(new_n688), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n747), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n250), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n813), .A2(KEYINPUT57), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n806), .A2(G148gat), .A3(new_n617), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n827), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n815), .A2(new_n617), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n825), .A2(KEYINPUT59), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n841), .ZN(G1345gat));
  NAND2_X1  g641(.A1(new_n565), .A2(G155gat), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT120), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n806), .A2(new_n818), .A3(new_n565), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n815), .A2(new_n844), .B1(new_n217), .B2(new_n845), .ZN(G1346gat));
  NOR3_X1   g645(.A1(new_n812), .A2(new_n662), .A3(new_n814), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n652), .A2(new_n218), .ZN(new_n848));
  OAI22_X1  g647(.A1(new_n847), .A2(new_n218), .B1(new_n826), .B2(new_n848), .ZN(G1347gat));
  OAI21_X1  g648(.A(new_n777), .B1(new_n778), .B2(new_n661), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n565), .B1(new_n850), .B2(new_n748), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n809), .B1(new_n779), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(new_n382), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n853), .A2(new_n405), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n348), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT121), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n857), .A2(new_n284), .A3(new_n530), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n852), .A2(new_n531), .A3(new_n855), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n284), .B2(new_n859), .ZN(G1348gat));
  AOI21_X1  g659(.A(new_n285), .B1(new_n856), .B2(new_n655), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n618), .A2(G176gat), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n861), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT122), .ZN(G1349gat));
  NAND2_X1  g663(.A1(new_n856), .A2(new_n565), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n272), .A2(G183gat), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n274), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n268), .B2(new_n865), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n868), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g668(.A(new_n267), .B1(new_n856), .B2(new_n652), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT61), .Z(new_n871));
  NOR2_X1   g670(.A1(new_n662), .A2(G190gat), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n857), .A2(KEYINPUT123), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT123), .B1(new_n857), .B2(new_n872), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n871), .B1(new_n873), .B2(new_n874), .ZN(G1351gat));
  AND3_X1   g674(.A1(new_n636), .A2(new_n638), .A3(new_n854), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n835), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G197gat), .B1(new_n877), .B2(new_n531), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n818), .A2(new_n876), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n879), .A2(G197gat), .A3(new_n531), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1352gat));
  OR2_X1    g680(.A1(new_n618), .A2(G204gat), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G204gat), .B1(new_n877), .B2(new_n654), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n885), .B(new_n886), .C1(new_n890), .C2(new_n891), .ZN(G1353gat));
  OAI21_X1  g691(.A(KEYINPUT57), .B1(new_n852), .B2(new_n442), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n831), .A2(new_n834), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n565), .A3(new_n894), .A4(new_n876), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n835), .A2(KEYINPUT125), .A3(new_n565), .A4(new_n876), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n897), .A2(new_n898), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT126), .ZN(new_n900));
  INV_X1    g699(.A(G211gat), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n895), .B2(new_n896), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n898), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n902), .A2(new_n906), .A3(KEYINPUT63), .A4(new_n898), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n900), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n818), .A2(new_n901), .A3(new_n565), .A4(new_n876), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(G1354gat));
  OR2_X1    g709(.A1(new_n877), .A2(KEYINPUT127), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n877), .A2(KEYINPUT127), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n911), .A2(new_n652), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G218gat), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n662), .A2(G218gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n879), .B2(new_n915), .ZN(G1355gat));
endmodule


