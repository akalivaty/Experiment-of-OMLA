

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593;

  XNOR2_X1 U321 ( .A(n375), .B(KEYINPUT48), .ZN(n547) );
  NOR2_X2 U322 ( .A1(n565), .A2(n564), .ZN(n573) );
  XNOR2_X1 U323 ( .A(n480), .B(KEYINPUT104), .ZN(n481) );
  XNOR2_X1 U324 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U325 ( .A(n388), .B(n387), .ZN(n389) );
  AND2_X1 U326 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  INV_X1 U327 ( .A(KEYINPUT110), .ZN(n361) );
  XNOR2_X1 U328 ( .A(n364), .B(KEYINPUT47), .ZN(n365) );
  INV_X1 U329 ( .A(G204GAT), .ZN(n387) );
  INV_X1 U330 ( .A(KEYINPUT88), .ZN(n379) );
  XNOR2_X1 U331 ( .A(n331), .B(n330), .ZN(n337) );
  XNOR2_X1 U332 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U333 ( .A(n337), .B(n336), .ZN(n342) );
  XNOR2_X1 U334 ( .A(n382), .B(n381), .ZN(n457) );
  XNOR2_X1 U335 ( .A(n482), .B(n481), .ZN(n521) );
  XOR2_X1 U336 ( .A(n393), .B(n392), .Z(n497) );
  INV_X1 U337 ( .A(G43GAT), .ZN(n485) );
  XNOR2_X1 U338 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U339 ( .A(n485), .B(KEYINPUT40), .ZN(n486) );
  XNOR2_X1 U340 ( .A(n462), .B(n461), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n487), .B(n486), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n291) );
  XNOR2_X1 U343 ( .A(G92GAT), .B(KEYINPUT76), .ZN(n290) );
  XNOR2_X1 U344 ( .A(n291), .B(n290), .ZN(n295) );
  XOR2_X1 U345 ( .A(G99GAT), .B(G85GAT), .Z(n332) );
  XOR2_X1 U346 ( .A(KEYINPUT10), .B(n332), .Z(n293) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  XNOR2_X1 U348 ( .A(G218GAT), .B(n424), .ZN(n292) );
  XNOR2_X1 U349 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U350 ( .A(n295), .B(n294), .Z(n297) );
  NAND2_X1 U351 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U352 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U353 ( .A(KEYINPUT77), .B(KEYINPUT11), .Z(n299) );
  XNOR2_X1 U354 ( .A(G134GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U356 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U357 ( .A(G29GAT), .B(G43GAT), .Z(n303) );
  XNOR2_X1 U358 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n317) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n304) );
  XNOR2_X1 U361 ( .A(n304), .B(KEYINPUT78), .ZN(n386) );
  XNOR2_X1 U362 ( .A(n317), .B(n386), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n560) );
  XOR2_X1 U364 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n308) );
  XNOR2_X1 U365 ( .A(G22GAT), .B(KEYINPUT29), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n325) );
  XOR2_X1 U367 ( .A(G8GAT), .B(G141GAT), .Z(n310) );
  XNOR2_X1 U368 ( .A(G50GAT), .B(G36GAT), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U370 ( .A(G15GAT), .B(KEYINPUT70), .Z(n312) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(G197GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U373 ( .A(n314), .B(n313), .Z(n323) );
  XOR2_X1 U374 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n316) );
  XNOR2_X1 U375 ( .A(KEYINPUT67), .B(KEYINPUT71), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n316), .B(n315), .ZN(n321) );
  XOR2_X1 U377 ( .A(G113GAT), .B(G1GAT), .Z(n412) );
  XOR2_X1 U378 ( .A(n317), .B(n412), .Z(n319) );
  NAND2_X1 U379 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U380 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U382 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U383 ( .A(n325), .B(n324), .ZN(n581) );
  INV_X1 U384 ( .A(n581), .ZN(n509) );
  XOR2_X1 U385 ( .A(G176GAT), .B(G92GAT), .Z(n326) );
  XOR2_X1 U386 ( .A(G64GAT), .B(n326), .Z(n392) );
  INV_X1 U387 ( .A(n392), .ZN(n327) );
  XOR2_X1 U388 ( .A(n327), .B(KEYINPUT31), .Z(n331) );
  XOR2_X1 U389 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n329) );
  XNOR2_X1 U390 ( .A(G120GAT), .B(KEYINPUT72), .ZN(n328) );
  XNOR2_X1 U391 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n332), .B(n289), .ZN(n334) );
  XNOR2_X1 U393 ( .A(G71GAT), .B(G57GAT), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n333), .B(KEYINPUT13), .ZN(n350) );
  XNOR2_X1 U395 ( .A(n334), .B(n350), .ZN(n335) );
  XOR2_X1 U396 ( .A(n335), .B(KEYINPUT32), .Z(n336) );
  XOR2_X1 U397 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n339) );
  XNOR2_X1 U398 ( .A(G204GAT), .B(G78GAT), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n339), .B(n338), .ZN(n341) );
  XOR2_X1 U400 ( .A(G148GAT), .B(G106GAT), .Z(n340) );
  XOR2_X1 U401 ( .A(n341), .B(n340), .Z(n427) );
  XOR2_X1 U402 ( .A(n342), .B(n427), .Z(n370) );
  XNOR2_X1 U403 ( .A(n370), .B(KEYINPUT41), .ZN(n553) );
  NOR2_X1 U404 ( .A1(n509), .A2(n553), .ZN(n343) );
  XNOR2_X1 U405 ( .A(n343), .B(KEYINPUT46), .ZN(n360) );
  XOR2_X1 U406 ( .A(KEYINPUT81), .B(G78GAT), .Z(n345) );
  XNOR2_X1 U407 ( .A(G211GAT), .B(KEYINPUT80), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n349) );
  XOR2_X1 U409 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n347) );
  XNOR2_X1 U410 ( .A(KEYINPUT70), .B(KEYINPUT14), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n359) );
  XOR2_X1 U413 ( .A(G15GAT), .B(G127GAT), .Z(n449) );
  XOR2_X1 U414 ( .A(n350), .B(KEYINPUT79), .Z(n352) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n449), .B(n353), .ZN(n357) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G155GAT), .Z(n423) );
  XOR2_X1 U419 ( .A(n423), .B(G64GAT), .Z(n355) );
  XOR2_X1 U420 ( .A(G8GAT), .B(G183GAT), .Z(n383) );
  XNOR2_X1 U421 ( .A(G1GAT), .B(n383), .ZN(n354) );
  XNOR2_X1 U422 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U423 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U424 ( .A(n359), .B(n358), .Z(n488) );
  INV_X1 U425 ( .A(n488), .ZN(n586) );
  NOR2_X1 U426 ( .A1(n360), .A2(n586), .ZN(n362) );
  XNOR2_X1 U427 ( .A(n362), .B(n361), .ZN(n363) );
  NOR2_X1 U428 ( .A1(n560), .A2(n363), .ZN(n366) );
  INV_X1 U429 ( .A(KEYINPUT111), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n374) );
  XOR2_X1 U431 ( .A(KEYINPUT36), .B(KEYINPUT102), .Z(n367) );
  XNOR2_X1 U432 ( .A(n560), .B(n367), .ZN(n591) );
  NOR2_X1 U433 ( .A1(n488), .A2(n591), .ZN(n368) );
  XOR2_X1 U434 ( .A(KEYINPUT45), .B(n368), .Z(n369) );
  NOR2_X1 U435 ( .A1(n581), .A2(n369), .ZN(n372) );
  INV_X1 U436 ( .A(n370), .ZN(n371) );
  NAND2_X1 U437 ( .A1(n372), .A2(n371), .ZN(n373) );
  NAND2_X1 U438 ( .A1(n374), .A2(n373), .ZN(n375) );
  XOR2_X1 U439 ( .A(G211GAT), .B(KEYINPUT21), .Z(n377) );
  XNOR2_X1 U440 ( .A(G197GAT), .B(G218GAT), .ZN(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n429) );
  XNOR2_X1 U442 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n378) );
  XNOR2_X1 U443 ( .A(n378), .B(KEYINPUT18), .ZN(n382) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(KEYINPUT87), .ZN(n380) );
  XOR2_X1 U445 ( .A(n457), .B(n383), .Z(n385) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n386), .B(KEYINPUT97), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n429), .B(n391), .ZN(n393) );
  NAND2_X1 U450 ( .A1(n547), .A2(n497), .ZN(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n420) );
  XOR2_X1 U453 ( .A(G120GAT), .B(KEYINPUT83), .Z(n397) );
  XNOR2_X1 U454 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n396) );
  XNOR2_X1 U455 ( .A(n397), .B(n396), .ZN(n448) );
  XOR2_X1 U456 ( .A(G127GAT), .B(n448), .Z(n399) );
  NAND2_X1 U457 ( .A1(G225GAT), .A2(G233GAT), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n419) );
  XOR2_X1 U459 ( .A(G57GAT), .B(KEYINPUT1), .Z(n401) );
  XNOR2_X1 U460 ( .A(KEYINPUT6), .B(KEYINPUT93), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n405) );
  XOR2_X1 U462 ( .A(G148GAT), .B(KEYINPUT5), .Z(n403) );
  XNOR2_X1 U463 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U465 ( .A(n405), .B(n404), .Z(n417) );
  XOR2_X1 U466 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n407) );
  XNOR2_X1 U467 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n406) );
  XNOR2_X1 U468 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U469 ( .A(G141GAT), .B(n408), .Z(n437) );
  XOR2_X1 U470 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n410) );
  XNOR2_X1 U471 ( .A(G162GAT), .B(G85GAT), .ZN(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U473 ( .A(n411), .B(G155GAT), .Z(n414) );
  XNOR2_X1 U474 ( .A(G29GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U475 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U476 ( .A(n437), .B(n415), .ZN(n416) );
  XNOR2_X1 U477 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U478 ( .A(n419), .B(n418), .Z(n523) );
  NAND2_X1 U479 ( .A1(n420), .A2(n523), .ZN(n422) );
  INV_X1 U480 ( .A(KEYINPUT64), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n577) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n426) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n433) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(KEYINPUT92), .Z(n431) );
  INV_X1 U486 ( .A(n427), .ZN(n428) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U489 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U492 ( .A(n437), .B(n436), .ZN(n470) );
  NAND2_X1 U493 ( .A1(n577), .A2(n470), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n438), .B(KEYINPUT55), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n439), .B(KEYINPUT121), .ZN(n564) );
  XOR2_X1 U496 ( .A(G190GAT), .B(G99GAT), .Z(n441) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G113GAT), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U499 ( .A(KEYINPUT84), .B(G71GAT), .Z(n443) );
  XNOR2_X1 U500 ( .A(G176GAT), .B(G183GAT), .ZN(n442) );
  XNOR2_X1 U501 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U502 ( .A(n445), .B(n444), .Z(n455) );
  XOR2_X1 U503 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n447) );
  XNOR2_X1 U504 ( .A(KEYINPUT89), .B(KEYINPUT86), .ZN(n446) );
  XNOR2_X1 U505 ( .A(n447), .B(n446), .ZN(n453) );
  XOR2_X1 U506 ( .A(n449), .B(n448), .Z(n451) );
  NAND2_X1 U507 ( .A1(G227GAT), .A2(G233GAT), .ZN(n450) );
  XNOR2_X1 U508 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U511 ( .A(n457), .B(n456), .Z(n469) );
  NAND2_X1 U512 ( .A1(n469), .A2(n560), .ZN(n458) );
  NOR2_X1 U513 ( .A1(n564), .A2(n458), .ZN(n462) );
  XNOR2_X1 U514 ( .A(KEYINPUT58), .B(KEYINPUT124), .ZN(n460) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n459) );
  XNOR2_X1 U516 ( .A(KEYINPUT27), .B(n497), .ZN(n472) );
  INV_X1 U517 ( .A(n472), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n523), .A2(n463), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(n464), .Z(n546) );
  XNOR2_X1 U520 ( .A(KEYINPUT28), .B(n470), .ZN(n530) );
  INV_X1 U521 ( .A(n530), .ZN(n465) );
  NOR2_X1 U522 ( .A1(n546), .A2(n465), .ZN(n533) );
  INV_X1 U523 ( .A(n469), .ZN(n565) );
  NAND2_X1 U524 ( .A1(n533), .A2(n565), .ZN(n477) );
  NAND2_X1 U525 ( .A1(n497), .A2(n469), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n466), .A2(n470), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n467), .B(KEYINPUT99), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT25), .ZN(n474) );
  NOR2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT26), .ZN(n578) );
  NAND2_X1 U531 ( .A1(n472), .A2(n578), .ZN(n473) );
  NAND2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n523), .A2(n475), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n491) );
  NAND2_X1 U535 ( .A1(n491), .A2(n488), .ZN(n478) );
  XOR2_X1 U536 ( .A(KEYINPUT103), .B(n478), .Z(n479) );
  NOR2_X1 U537 ( .A1(n591), .A2(n479), .ZN(n482) );
  INV_X1 U538 ( .A(KEYINPUT37), .ZN(n480) );
  NOR2_X1 U539 ( .A1(n509), .A2(n370), .ZN(n493) );
  AND2_X1 U540 ( .A1(n521), .A2(n493), .ZN(n484) );
  INV_X1 U541 ( .A(KEYINPUT38), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(n507) );
  NOR2_X1 U543 ( .A1(n507), .A2(n565), .ZN(n487) );
  NOR2_X1 U544 ( .A1(n560), .A2(n488), .ZN(n490) );
  XNOR2_X1 U545 ( .A(KEYINPUT82), .B(KEYINPUT16), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n490), .B(n489), .ZN(n492) );
  AND2_X1 U547 ( .A1(n492), .A2(n491), .ZN(n510) );
  NAND2_X1 U548 ( .A1(n493), .A2(n510), .ZN(n494) );
  XNOR2_X1 U549 ( .A(KEYINPUT100), .B(n494), .ZN(n502) );
  NOR2_X1 U550 ( .A1(n523), .A2(n502), .ZN(n495) );
  XOR2_X1 U551 ( .A(G1GAT), .B(n495), .Z(n496) );
  XNOR2_X1 U552 ( .A(KEYINPUT34), .B(n496), .ZN(G1324GAT) );
  XNOR2_X1 U553 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n499) );
  INV_X1 U554 ( .A(n497), .ZN(n525) );
  NOR2_X1 U555 ( .A1(n525), .A2(n502), .ZN(n498) );
  XNOR2_X1 U556 ( .A(n499), .B(n498), .ZN(G1325GAT) );
  NOR2_X1 U557 ( .A1(n502), .A2(n565), .ZN(n501) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(G1326GAT) );
  NOR2_X1 U560 ( .A1(n530), .A2(n502), .ZN(n503) );
  XOR2_X1 U561 ( .A(G22GAT), .B(n503), .Z(G1327GAT) );
  NOR2_X1 U562 ( .A1(n523), .A2(n507), .ZN(n504) );
  XNOR2_X1 U563 ( .A(n504), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n525), .A2(n507), .ZN(n506) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  NOR2_X1 U567 ( .A1(n530), .A2(n507), .ZN(n508) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n508), .Z(G1331GAT) );
  XNOR2_X1 U569 ( .A(n553), .B(KEYINPUT105), .ZN(n570) );
  AND2_X1 U570 ( .A1(n570), .A2(n509), .ZN(n522) );
  NAND2_X1 U571 ( .A1(n522), .A2(n510), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n523), .A2(n517), .ZN(n511) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n511), .Z(n512) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n512), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n525), .A2(n517), .ZN(n514) );
  XNOR2_X1 U576 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  NOR2_X1 U579 ( .A1(n565), .A2(n517), .ZN(n516) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n516), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n530), .A2(n517), .ZN(n519) );
  XNOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n523), .A2(n529), .ZN(n524) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n524), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n525), .A2(n529), .ZN(n526) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n526), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n565), .A2(n529), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n531), .Z(n532) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U596 ( .A1(n547), .A2(n533), .ZN(n534) );
  NOR2_X1 U597 ( .A1(n565), .A2(n534), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n581), .A2(n543), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT112), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n538) );
  NAND2_X1 U602 ( .A1(n543), .A2(n570), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U604 ( .A(G120GAT), .B(n539), .Z(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n541) );
  NAND2_X1 U606 ( .A1(n543), .A2(n586), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n542), .Z(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U610 ( .A1(n543), .A2(n560), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n550) );
  NAND2_X1 U613 ( .A1(n547), .A2(n578), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n546), .A2(n548), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n561), .A2(n581), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  INV_X1 U618 ( .A(n561), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n555) );
  XNOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(n556), .B(KEYINPUT52), .Z(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(KEYINPUT117), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n586), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n573), .A2(n581), .ZN(n566) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n568) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(n569), .Z(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n586), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT60), .ZN(n576) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(n576), .Z(n583) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n580) );
  INV_X1 U644 ( .A(KEYINPUT125), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n590) );
  INV_X1 U646 ( .A(n590), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U650 ( .A1(n587), .A2(n370), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

