//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n196), .C1(new_n197), .C2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n199), .B(G134), .C1(KEYINPUT64), .C2(KEYINPUT11), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n197), .A2(G137), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n201));
  INV_X1    g015(.A(G131), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n200), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(new_n189), .B(new_n192), .C1(KEYINPUT1), .C2(new_n187), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n197), .A2(G137), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n199), .A2(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n194), .A2(new_n203), .A3(new_n204), .A4(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT68), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n189), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n210));
  XNOR2_X1  g024(.A(G143), .B(G146), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G131), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(KEYINPUT67), .A3(new_n203), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(KEYINPUT67), .B1(new_n216), .B2(new_n203), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n214), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n209), .A2(new_n220), .A3(KEYINPUT30), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n213), .B1(new_n203), .B2(new_n216), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n208), .B1(new_n223), .B2(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n203), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n225), .A2(KEYINPUT65), .A3(new_n214), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G119), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT66), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(G116), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n232), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT2), .A2(G113), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT2), .A2(G113), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G116), .B(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n221), .A2(new_n227), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT69), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n209), .A2(new_n220), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(G237), .A2(G953), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G210), .ZN(new_n252));
  INV_X1    g066(.A(G101), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n254), .B(new_n255), .Z(new_n256));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n221), .A2(new_n227), .A3(new_n257), .A4(new_n245), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n247), .A2(new_n250), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT31), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n224), .A2(new_n226), .ZN(new_n261));
  INV_X1    g075(.A(new_n245), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n249), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n208), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT28), .B1(new_n266), .B2(new_n220), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n256), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n249), .B1(new_n246), .B2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n256), .A4(new_n258), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n260), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(G472), .A2(G902), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT32), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(KEYINPUT32), .A3(new_n276), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT70), .B(G902), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n248), .B(new_n245), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n267), .B1(new_n281), .B2(KEYINPUT28), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT29), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n270), .A2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n283), .B1(new_n269), .B2(new_n270), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n256), .B1(new_n272), .B2(new_n258), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G472), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n278), .A2(new_n279), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G469), .ZN(new_n291));
  INV_X1    g105(.A(new_n280), .ZN(new_n292));
  INV_X1    g106(.A(G107), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(G104), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n295));
  INV_X1    g109(.A(G104), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n295), .B1(new_n296), .B2(G107), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n293), .A2(KEYINPUT3), .A3(G104), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n296), .A2(G107), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n253), .B1(new_n300), .B2(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n296), .A2(G107), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n293), .A2(G104), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n299), .A2(new_n253), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(new_n204), .A3(new_n194), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT10), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n218), .A2(new_n219), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n299), .A2(new_n253), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n299), .A2(new_n253), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(KEYINPUT4), .A3(new_n311), .ZN(new_n312));
  OR3_X1    g126(.A1(new_n299), .A2(KEYINPUT4), .A3(new_n253), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n214), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n309), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n194), .A2(new_n204), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(new_n306), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n225), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT12), .ZN(new_n320));
  XNOR2_X1  g134(.A(G110), .B(G140), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G227), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n309), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT12), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(new_n318), .ZN(new_n327));
  AND4_X1   g141(.A1(new_n315), .A2(new_n320), .A3(new_n324), .A4(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT10), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n307), .B(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n314), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n324), .B1(new_n332), .B2(new_n315), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n291), .B(new_n292), .C1(new_n328), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(G469), .A2(G902), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n332), .A2(new_n315), .A3(new_n324), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n315), .A2(new_n320), .A3(new_n327), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n336), .B1(new_n338), .B2(new_n324), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n334), .B(new_n335), .C1(new_n339), .C2(new_n291), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  OAI21_X1  g155(.A(G221), .B1(new_n341), .B2(G902), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT90), .ZN(new_n344));
  AND2_X1   g158(.A1(KEYINPUT74), .A2(G125), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT74), .A2(G125), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT16), .ZN(new_n348));
  INV_X1    g162(.A(G140), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(G125), .A2(G140), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(new_n347), .B2(G140), .ZN(new_n352));
  OAI211_X1 g166(.A(G146), .B(new_n350), .C1(new_n352), .C2(new_n348), .ZN(new_n353));
  XNOR2_X1  g167(.A(G125), .B(G140), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT19), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OR2_X1    g170(.A1(KEYINPUT74), .A2(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT74), .A2(G125), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(G140), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(new_n351), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n356), .B1(new_n361), .B2(new_n355), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n353), .B1(new_n362), .B2(G146), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT86), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n251), .A2(G143), .A3(G214), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G143), .B1(new_n251), .B2(G214), .ZN(new_n367));
  OAI21_X1  g181(.A(G131), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n367), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n202), .A3(new_n365), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n353), .B(new_n372), .C1(new_n362), .C2(G146), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G113), .B(G122), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n375), .B(new_n296), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT84), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n369), .A3(new_n365), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT85), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n352), .A2(G146), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n354), .A2(new_n188), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n202), .B1(new_n369), .B2(new_n365), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n382), .A2(new_n383), .B1(new_n384), .B2(KEYINPUT18), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n374), .A2(new_n377), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n381), .A2(new_n385), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n348), .B1(new_n359), .B2(new_n360), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n357), .A2(new_n358), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n392), .A2(KEYINPUT16), .A3(G140), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n188), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n390), .B1(new_n394), .B2(new_n353), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n353), .A3(new_n390), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT88), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n371), .B2(KEYINPUT17), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT17), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT88), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n384), .A2(KEYINPUT17), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n389), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n387), .B(new_n388), .C1(new_n405), .C2(new_n377), .ZN(new_n406));
  NOR2_X1   g220(.A1(G475), .A2(G902), .ZN(new_n407));
  XOR2_X1   g221(.A(new_n407), .B(KEYINPUT89), .Z(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n344), .B1(new_n406), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n387), .B(new_n407), .C1(new_n405), .C2(new_n377), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT20), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n394), .A2(new_n353), .A3(new_n390), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n395), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n386), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n389), .A2(new_n376), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n416), .A2(new_n376), .B1(new_n417), .B2(new_n374), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n418), .A2(KEYINPUT90), .A3(new_n388), .A4(new_n408), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n410), .A2(new_n412), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n377), .A2(KEYINPUT91), .ZN(new_n421));
  AOI21_X1  g235(.A(G902), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n405), .A2(KEYINPUT91), .A3(new_n377), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G475), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G217), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n341), .A2(new_n427), .A3(G953), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n228), .B2(G122), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G107), .ZN(new_n430));
  XNOR2_X1  g244(.A(G116), .B(G122), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n431), .ZN(new_n433));
  XNOR2_X1  g247(.A(G128), .B(G143), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n197), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n434), .A2(new_n197), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n432), .B(new_n433), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n434), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(G128), .A3(new_n191), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT93), .A4(G134), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n431), .B(new_n293), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n435), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n197), .B1(new_n440), .B2(new_n434), .ZN(new_n446));
  AOI21_X1  g260(.A(KEYINPUT93), .B1(new_n446), .B2(new_n442), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n428), .B(new_n438), .C1(new_n445), .C2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n441), .A2(G134), .A3(new_n442), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(new_n443), .A3(new_n444), .A4(new_n435), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n428), .B1(new_n453), .B2(new_n438), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n292), .B1(new_n449), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(G478), .ZN(new_n456));
  NOR2_X1   g270(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(KEYINPUT94), .A2(KEYINPUT15), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n455), .A2(KEYINPUT95), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n438), .B1(new_n445), .B2(new_n447), .ZN(new_n463));
  INV_X1    g277(.A(new_n428), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n280), .B1(new_n465), .B2(new_n448), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n455), .A2(KEYINPUT95), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(G234), .A2(G237), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n471), .A2(G952), .A3(new_n322), .ZN(new_n472));
  XNOR2_X1  g286(.A(KEYINPUT21), .B(G898), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(KEYINPUT96), .Z(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n280), .A2(G953), .A3(new_n471), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g293(.A1(new_n343), .A2(new_n426), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n230), .A2(G128), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n187), .A2(G119), .ZN(new_n482));
  OR3_X1    g296(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT71), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT71), .B1(new_n481), .B2(new_n482), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT24), .B(G110), .Z(new_n486));
  OAI21_X1  g300(.A(new_n481), .B1(KEYINPUT72), .B2(KEYINPUT23), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT23), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT72), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n230), .B2(G128), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n485), .A2(new_n486), .B1(G110), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n353), .A3(new_n383), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n394), .A2(new_n353), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n486), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n492), .A2(KEYINPUT73), .A3(G110), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n492), .A2(G110), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT22), .B(G137), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n322), .A2(G221), .A3(G234), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n503), .B(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n501), .A3(new_n505), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n427), .B1(new_n292), .B2(G234), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n510), .A2(G902), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(new_n292), .A3(new_n508), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT25), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n507), .A2(KEYINPUT25), .A3(new_n292), .A4(new_n508), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n512), .B1(new_n517), .B2(new_n510), .ZN(new_n518));
  OAI21_X1  g332(.A(G214), .B1(G237), .B2(G902), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n316), .A2(new_n392), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n213), .A2(new_n347), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G224), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G953), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n523), .B(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n232), .A2(KEYINPUT5), .A3(new_n236), .ZN(new_n527));
  INV_X1    g341(.A(G113), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT5), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n229), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n530), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n533), .A2(new_n244), .A3(new_n306), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n312), .A2(new_n245), .A3(new_n313), .ZN(new_n536));
  XNOR2_X1  g350(.A(G110), .B(G122), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n537), .B(KEYINPUT77), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT78), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n535), .B2(new_n536), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n538), .B1(new_n541), .B2(KEYINPUT6), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT6), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n543), .B(new_n540), .C1(new_n535), .C2(new_n536), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n526), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT79), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n547), .B(new_n526), .C1(new_n542), .C2(new_n544), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n538), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n537), .B(KEYINPUT8), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT80), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n233), .A2(new_n234), .A3(KEYINPUT5), .ZN(new_n554));
  AOI22_X1  g368(.A1(new_n530), .A2(new_n554), .B1(new_n240), .B2(new_n243), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n306), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n554), .ZN(new_n557));
  OAI21_X1  g371(.A(G113), .B1(new_n233), .B2(KEYINPUT5), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n553), .B(new_n244), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n552), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n244), .B1(new_n557), .B2(new_n558), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(KEYINPUT80), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n563), .A2(KEYINPUT81), .A3(new_n306), .A4(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n531), .A2(new_n532), .B1(new_n240), .B2(new_n243), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n306), .B1(new_n566), .B2(new_n534), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n551), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT82), .B1(new_n524), .B2(G953), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n523), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n571), .B2(new_n525), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n525), .A2(new_n571), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n523), .A2(new_n569), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT83), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n550), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n568), .A2(KEYINPUT83), .A3(new_n575), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n549), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G210), .B1(G237), .B2(G902), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n549), .A2(new_n580), .A3(new_n582), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n520), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n290), .A2(new_n480), .A3(new_n518), .A4(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  NAND2_X1  g402(.A1(new_n275), .A2(new_n292), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n589), .A2(G472), .B1(new_n275), .B2(new_n276), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n340), .A2(new_n518), .A3(new_n342), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT97), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n584), .A2(new_n597), .A3(new_n585), .ZN(new_n598));
  AND3_X1   g412(.A1(new_n549), .A2(new_n580), .A3(new_n582), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT98), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n598), .A2(new_n519), .A3(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n425), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n418), .A2(new_n388), .A3(new_n408), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n603), .A2(new_n344), .B1(KEYINPUT20), .B2(new_n411), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n604), .B2(new_n419), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n449), .A2(new_n454), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(KEYINPUT99), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT99), .B(KEYINPUT33), .Z(new_n610));
  AOI21_X1  g424(.A(new_n609), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n280), .A2(new_n456), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n466), .B2(G478), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n455), .A2(KEYINPUT100), .A3(new_n456), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n605), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n601), .A2(KEYINPUT101), .A3(new_n478), .A4(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n598), .A2(new_n519), .A3(new_n478), .A4(new_n600), .ZN(new_n620));
  INV_X1    g434(.A(new_n617), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n596), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT34), .B(G104), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G6));
  NAND3_X1  g439(.A1(new_n418), .A2(new_n388), .A3(new_n407), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n626), .B1(new_n412), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT102), .B1(new_n411), .B2(KEYINPUT20), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OR3_X1    g444(.A1(new_n630), .A2(new_n602), .A3(new_n470), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n620), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(new_n596), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  AND2_X1   g449(.A1(new_n517), .A2(new_n510), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT103), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n502), .B(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n639), .A2(new_n511), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n480), .A2(new_n586), .A3(new_n590), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G110), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n643), .B(new_n645), .ZN(G12));
  NAND2_X1  g460(.A1(new_n598), .A2(new_n600), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n520), .A3(new_n343), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n275), .A2(KEYINPUT32), .A3(new_n276), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n649), .A2(new_n277), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n641), .B1(new_n650), .B2(new_n289), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n472), .B1(new_n476), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n631), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  AOI21_X1  g471(.A(new_n582), .B1(new_n549), .B2(new_n580), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n599), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT38), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n654), .B(KEYINPUT39), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n343), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(G472), .ZN(new_n665));
  INV_X1    g479(.A(new_n281), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n259), .B1(new_n666), .B2(new_n256), .ZN(new_n667));
  INV_X1    g481(.A(G902), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n650), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n605), .A2(new_n520), .A3(new_n470), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n641), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n660), .A2(new_n664), .A3(new_n670), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  NAND2_X1  g488(.A1(new_n614), .A2(new_n615), .ZN(new_n675));
  INV_X1    g489(.A(new_n611), .ZN(new_n676));
  INV_X1    g490(.A(new_n612), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n654), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n426), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n652), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  INV_X1    g497(.A(new_n518), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n650), .B2(new_n289), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n328), .A2(new_n333), .ZN(new_n686));
  OAI21_X1  g500(.A(G469), .B1(new_n686), .B2(new_n280), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n687), .A2(new_n342), .A3(new_n334), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT106), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n687), .A2(new_n690), .A3(new_n342), .A4(new_n334), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n618), .B2(new_n622), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT41), .B(G113), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NOR2_X1   g510(.A1(new_n632), .A2(new_n693), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n228), .ZN(G18));
  NOR2_X1   g512(.A1(new_n426), .A2(new_n479), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n290), .A2(new_n699), .A3(new_n642), .ZN(new_n700));
  INV_X1    g514(.A(new_n688), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n598), .A2(new_n519), .A3(new_n600), .A4(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT108), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n708), .B(new_n700), .C1(new_n704), .C2(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT109), .B(G119), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G21));
  AND2_X1   g526(.A1(new_n598), .A2(new_n600), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n477), .B1(new_n689), .B2(new_n691), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(new_n671), .A3(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n260), .B(new_n274), .C1(new_n256), .C2(new_n282), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n276), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n665), .B1(new_n275), .B2(new_n292), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n717), .B1(new_n718), .B2(KEYINPUT110), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n720), .B(new_n665), .C1(new_n275), .C2(new_n292), .ZN(new_n721));
  OR3_X1    g535(.A1(new_n719), .A2(new_n684), .A3(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n715), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(G122), .Z(G24));
  NOR4_X1   g538(.A1(new_n719), .A2(new_n721), .A3(new_n680), .A4(new_n641), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n704), .B2(new_n705), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND3_X1  g541(.A1(new_n584), .A2(new_n585), .A3(new_n519), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n334), .A2(new_n335), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n336), .B(KEYINPUT112), .ZN(new_n732));
  INV_X1    g546(.A(new_n324), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT111), .B1(new_n337), .B2(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n337), .A2(KEYINPUT111), .A3(new_n733), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n731), .B1(new_n736), .B2(new_n291), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(new_n342), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n584), .A2(KEYINPUT113), .A3(new_n585), .A4(new_n519), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n730), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n290), .A2(new_n518), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT42), .B1(new_n742), .B2(new_n681), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR4_X1   g558(.A1(new_n740), .A2(new_n741), .A3(new_n744), .A4(new_n680), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n202), .ZN(G33));
  AOI21_X1  g561(.A(KEYINPUT113), .B1(new_n659), .B2(new_n519), .ZN(new_n748));
  INV_X1    g562(.A(new_n739), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n685), .A3(new_n655), .A4(new_n738), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  NOR2_X1   g566(.A1(new_n426), .A2(new_n616), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT43), .ZN(new_n754));
  INV_X1    g568(.A(new_n590), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n642), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT44), .Z(new_n757));
  INV_X1    g571(.A(new_n750), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n334), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n291), .B1(new_n339), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n736), .B2(new_n761), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n763), .A2(new_n335), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n764), .B2(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n765), .B1(KEYINPUT46), .B2(new_n764), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n342), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n661), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G137), .ZN(G39));
  XNOR2_X1  g584(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n767), .B(new_n771), .Z(new_n772));
  NOR3_X1   g586(.A1(new_n290), .A2(new_n518), .A3(new_n680), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n750), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G140), .ZN(G42));
  NAND3_X1  g589(.A1(new_n518), .A2(new_n519), .A3(new_n342), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT115), .Z(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n753), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT116), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n687), .A2(new_n334), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT49), .ZN(new_n781));
  OR4_X1    g595(.A1(new_n670), .A2(new_n779), .A3(new_n660), .A4(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n648), .B(new_n651), .C1(new_n655), .C2(new_n681), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n636), .A2(new_n640), .A3(new_n654), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n737), .A2(new_n785), .A3(new_n342), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n737), .A2(new_n785), .A3(KEYINPUT118), .A4(new_n342), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n713), .A3(new_n670), .A4(new_n671), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n726), .A2(new_n784), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n726), .A2(new_n784), .A3(KEYINPUT52), .A4(new_n791), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n730), .A2(new_n738), .A3(new_n739), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n725), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n470), .A2(KEYINPUT117), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n800), .B(new_n462), .C1(new_n468), .C2(new_n469), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n425), .A2(new_n679), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n343), .A2(new_n802), .A3(new_n630), .A4(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n750), .A2(new_n651), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n751), .A2(new_n798), .A3(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n420), .A2(new_n799), .A3(new_n425), .A4(new_n801), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n807), .B1(new_n605), .B2(new_n616), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n586), .A3(new_n478), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n587), .B(new_n643), .C1(new_n596), .C2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n797), .A2(new_n685), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n744), .B1(new_n812), .B2(new_n680), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n742), .A2(KEYINPUT42), .A3(new_n681), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n632), .A2(new_n693), .B1(new_n715), .B2(new_n722), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(new_n694), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n710), .A2(new_n811), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n783), .B1(new_n796), .B2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT119), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n710), .A2(new_n817), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n794), .A2(new_n795), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n590), .A2(KEYINPUT97), .A3(new_n591), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT97), .B1(new_n590), .B2(new_n591), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n809), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n587), .A2(new_n643), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n751), .A3(new_n798), .A4(new_n805), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n746), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n821), .A2(new_n822), .A3(new_n829), .A4(KEYINPUT53), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n819), .A2(new_n820), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(KEYINPUT119), .B(new_n783), .C1(new_n796), .C2(new_n818), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT54), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n819), .A2(new_n830), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n833), .B1(KEYINPUT54), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  INV_X1    g650(.A(new_n722), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n472), .A3(new_n754), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n772), .A2(KEYINPUT120), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n780), .A2(new_n342), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n772), .B2(KEYINPUT120), .ZN(new_n841));
  AOI211_X1 g655(.A(new_n758), .B(new_n838), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n838), .A2(new_n519), .A3(new_n660), .A4(new_n688), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT50), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n750), .A2(new_n472), .A3(new_n701), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n754), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n719), .A2(new_n641), .A3(new_n721), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n845), .A2(new_n684), .A3(new_n670), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n426), .A2(new_n678), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n848), .A2(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n836), .B1(new_n842), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n772), .A2(new_n840), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n838), .A2(new_n758), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n836), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n844), .A3(new_n852), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n847), .A2(new_n741), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT48), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n850), .A2(new_n617), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(G952), .A3(new_n322), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n704), .A2(new_n705), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n838), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n835), .A2(new_n854), .A3(new_n858), .A4(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n782), .B1(new_n866), .B2(new_n867), .ZN(G75));
  NAND4_X1  g682(.A1(new_n831), .A2(new_n280), .A3(new_n583), .A4(new_n832), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT56), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n542), .A2(new_n544), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT121), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n870), .A3(new_n873), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g691(.A(new_n526), .B(KEYINPUT55), .Z(new_n878));
  AND2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n322), .A2(G952), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(G51));
  XOR2_X1   g696(.A(new_n335), .B(KEYINPUT57), .Z(new_n883));
  NAND3_X1  g697(.A1(new_n831), .A2(KEYINPUT54), .A3(new_n832), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(new_n833), .ZN(new_n886));
  INV_X1    g700(.A(new_n686), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(KEYINPUT122), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n831), .A2(new_n832), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n890), .A2(new_n292), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n763), .B(KEYINPUT123), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n888), .A2(KEYINPUT122), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n881), .B1(new_n889), .B2(new_n893), .ZN(G54));
  NAND3_X1  g708(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n895));
  INV_X1    g709(.A(new_n418), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n896), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n881), .ZN(G60));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  NOR2_X1   g716(.A1(new_n676), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n890), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n904), .B1(new_n906), .B2(new_n884), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n900), .B1(new_n907), .B2(new_n881), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n903), .B1(new_n885), .B2(new_n833), .ZN(new_n909));
  INV_X1    g723(.A(new_n881), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(KEYINPUT124), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n676), .B1(new_n835), .B2(new_n902), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n908), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(KEYINPUT125), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n908), .A2(new_n911), .A3(new_n912), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  NAND4_X1  g733(.A1(new_n831), .A2(new_n639), .A3(new_n832), .A4(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n831), .A2(new_n832), .A3(new_n919), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n910), .B(new_n920), .C1(new_n921), .C2(new_n509), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g737(.A(G953), .B1(new_n475), .B2(new_n524), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n821), .A2(new_n827), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n926), .B2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n874), .B1(G898), .B2(new_n322), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(G69));
  NAND2_X1  g743(.A1(new_n221), .A2(new_n227), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n362), .Z(new_n931));
  NAND2_X1  g745(.A1(new_n726), .A2(new_n784), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n673), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT62), .Z(new_n935));
  NAND4_X1  g749(.A1(new_n750), .A2(new_n685), .A3(new_n662), .A4(new_n808), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n769), .A2(new_n935), .A3(new_n774), .A4(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n937), .B2(G953), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n931), .B1(G900), .B2(G953), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n774), .A2(new_n751), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n685), .A2(new_n713), .A3(new_n671), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n768), .B1(new_n759), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n940), .A2(new_n815), .A3(new_n933), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n943), .B2(G953), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n938), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n945), .B(new_n948), .Z(G72));
  NAND2_X1  g763(.A1(G472), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT63), .Z(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n943), .B2(new_n925), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n270), .A3(new_n258), .A4(new_n272), .ZN(new_n953));
  INV_X1    g767(.A(new_n259), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n954), .A2(new_n287), .A3(KEYINPUT127), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n287), .A2(KEYINPUT127), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n834), .A2(new_n951), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n910), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n937), .A2(new_n926), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n951), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n270), .B1(new_n272), .B2(new_n258), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(G57));
endmodule


