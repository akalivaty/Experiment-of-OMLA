//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1311, new_n1312, new_n1313, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396, new_n1397, new_n1398, new_n1399, new_n1400;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  AND2_X1   g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  INV_X1    g0011(.A(new_n201), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G50), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT64), .Z(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G97), .ZN(new_n219));
  INV_X1    g0019(.A(G257), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n221), .A2(new_n222), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n209), .B1(new_n211), .B2(new_n215), .C1(new_n228), .C2(KEYINPUT1), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT67), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G226), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n234), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G58), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT13), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(KEYINPUT71), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(G232), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  AND2_X1   g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NOR2_X1   g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(G226), .B2(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(G33), .A2(G97), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n252), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G41), .ZN(new_n260));
  INV_X1    g0060(.A(G45), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(new_n252), .A3(G274), .ZN(new_n263));
  INV_X1    g0063(.A(G238), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n252), .A2(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n263), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n250), .B1(new_n259), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n259), .A2(new_n268), .A3(new_n250), .ZN(new_n271));
  OAI21_X1  g0071(.A(G179), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(KEYINPUT73), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(KEYINPUT72), .B2(KEYINPUT14), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT13), .B1(new_n259), .B2(new_n268), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n259), .A2(new_n268), .A3(KEYINPUT13), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(KEYINPUT72), .A2(KEYINPUT14), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT73), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(G179), .C1(new_n270), .C2(new_n271), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n275), .B(new_n280), .C1(new_n277), .C2(new_n278), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n273), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT74), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  INV_X1    g0089(.A(G68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT70), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n291), .A2(new_n265), .A3(G13), .A4(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT12), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n292), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G1), .A2(G13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G20), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G1), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n296), .A2(G68), .A3(new_n300), .A4(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(G33), .A3(G77), .ZN(new_n305));
  INV_X1    g0105(.A(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n305), .B1(new_n301), .B2(G68), .C1(new_n307), .C2(new_n202), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT11), .ZN(new_n309));
  AND3_X1   g0109(.A1(new_n308), .A2(new_n309), .A3(new_n299), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n309), .B1(new_n308), .B2(new_n299), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n287), .B1(new_n295), .B2(new_n312), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n310), .A2(new_n311), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n314), .A2(KEYINPUT74), .A3(new_n294), .A4(new_n304), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n286), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n259), .A2(new_n268), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n248), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n320), .B2(new_n276), .ZN(new_n321));
  INV_X1    g0121(.A(G190), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n249), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n269), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n314), .A2(new_n294), .A3(new_n304), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n321), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(G20), .A2(G77), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT15), .B(G87), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n301), .A2(G33), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n328), .B1(new_n329), .B2(new_n330), .C1(new_n307), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n299), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n296), .A2(G77), .A3(new_n300), .A4(new_n303), .ZN(new_n334));
  AND2_X1   g0134(.A1(new_n289), .A2(new_n292), .ZN(new_n335));
  INV_X1    g0135(.A(G77), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n255), .A2(new_n256), .ZN(new_n339));
  INV_X1    g0139(.A(G107), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n252), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n264), .A2(G1698), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G232), .B2(G1698), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n306), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n252), .A2(G244), .A3(new_n266), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n263), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n274), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n349), .A2(new_n354), .A3(new_n263), .A4(new_n351), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n338), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(G200), .B1(new_n350), .B2(new_n352), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n332), .A2(new_n299), .B1(new_n336), .B2(new_n335), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n349), .A2(G190), .A3(new_n263), .A4(new_n351), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n357), .A2(new_n358), .A3(new_n359), .A4(new_n334), .ZN(new_n360));
  AND4_X1   g0160(.A1(new_n317), .A2(new_n327), .A3(new_n356), .A4(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(G1698), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n347), .A2(G222), .A3(new_n362), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(KEYINPUT68), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n345), .B2(new_n346), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(G223), .B1(new_n339), .B2(G77), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n252), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G226), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n263), .B1(new_n370), .B2(new_n267), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n274), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n335), .A2(new_n299), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n302), .A2(new_n202), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(new_n202), .B2(new_n335), .ZN(new_n375));
  INV_X1    g0175(.A(new_n307), .ZN(new_n376));
  AOI22_X1  g0176(.A1(G150), .A2(new_n376), .B1(new_n203), .B2(G20), .ZN(new_n377));
  NOR2_X1   g0177(.A1(KEYINPUT8), .A2(G58), .ZN(new_n378));
  INV_X1    g0178(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT69), .B(G58), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT8), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n377), .B1(new_n382), .B2(new_n330), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n299), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n375), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n371), .ZN(new_n386));
  INV_X1    g0186(.A(new_n368), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(new_n364), .B2(new_n365), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n354), .B(new_n386), .C1(new_n388), .C2(new_n252), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n372), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT9), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n375), .A2(new_n384), .A3(KEYINPUT9), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT10), .ZN(new_n396));
  OAI211_X1 g0196(.A(G190), .B(new_n386), .C1(new_n388), .C2(new_n252), .ZN(new_n397));
  OAI21_X1  g0197(.A(G200), .B1(new_n369), .B2(new_n371), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n395), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(new_n393), .A3(new_n397), .A4(new_n394), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT10), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n391), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n382), .A2(new_n302), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n373), .A2(new_n403), .B1(new_n382), .B2(new_n335), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(G159), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n307), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(G58), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(KEYINPUT69), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT69), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(G58), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n201), .B1(new_n413), .B2(G68), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n408), .B1(new_n414), .B2(new_n301), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n345), .A2(new_n301), .A3(new_n346), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n301), .A4(new_n346), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n290), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n300), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n415), .B2(new_n420), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n405), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n263), .B1(new_n253), .B2(new_n267), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  OR2_X1    g0227(.A1(G223), .A2(G1698), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n370), .A2(G1698), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n428), .B(new_n429), .C1(new_n255), .C2(new_n256), .ZN(new_n430));
  NAND2_X1  g0230(.A1(G33), .A2(G87), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n252), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(new_n433), .A3(G179), .ZN(new_n434));
  OAI21_X1  g0234(.A(G169), .B1(new_n426), .B2(new_n432), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT18), .B1(new_n425), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT7), .B1(new_n339), .B2(new_n301), .ZN(new_n439));
  INV_X1    g0239(.A(new_n419), .ZN(new_n440));
  OAI21_X1  g0240(.A(G68), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n212), .B1(new_n380), .B2(new_n290), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n407), .B1(new_n442), .B2(G20), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n441), .A2(new_n443), .A3(KEYINPUT16), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n424), .A2(new_n444), .A3(new_n299), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n445), .A2(new_n404), .B1(new_n435), .B2(new_n434), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n318), .B1(new_n427), .B2(new_n433), .ZN(new_n449));
  AND2_X1   g0249(.A1(KEYINPUT75), .A2(G190), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT75), .A2(G190), .ZN(new_n451));
  OR2_X1    g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NOR3_X1   g0253(.A1(new_n426), .A2(new_n432), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n455), .A2(new_n445), .A3(new_n404), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT17), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n455), .A2(new_n445), .A3(KEYINPUT17), .A4(new_n404), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n438), .A2(new_n448), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n361), .A2(new_n402), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n335), .A2(G97), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n306), .A2(G1), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n296), .A2(new_n300), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n464), .B1(G97), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n376), .A2(G77), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n340), .A2(KEYINPUT6), .A3(G97), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT6), .ZN(new_n472));
  XNOR2_X1  g0272(.A(G97), .B(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n469), .B1(new_n474), .B2(new_n301), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n340), .B1(new_n418), .B2(new_n419), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n299), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT76), .ZN(new_n478));
  OAI21_X1  g0278(.A(G107), .B1(new_n439), .B2(new_n440), .ZN(new_n479));
  AND2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  NOR2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n472), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n470), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(G20), .B1(G77), .B2(new_n376), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT76), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n299), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n468), .B1(new_n478), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n261), .A2(G1), .ZN(new_n489));
  AND2_X1   g0289(.A1(KEYINPUT5), .A2(G41), .ZN(new_n490));
  NOR2_X1   g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G257), .A3(new_n252), .ZN(new_n493));
  INV_X1    g0293(.A(G274), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n210), .B2(new_n251), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT5), .B(G41), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n489), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G244), .B(new_n362), .C1(new_n255), .C2(new_n256), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(G1698), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n502), .B(G244), .C1(new_n256), .C2(new_n255), .ZN(new_n503));
  OAI211_X1 g0303(.A(G250), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n252), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G190), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT77), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n508), .B2(new_n318), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n512));
  INV_X1    g0312(.A(G244), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n345), .B2(new_n346), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT4), .B1(new_n514), .B2(new_n362), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n507), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n498), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(KEYINPUT77), .A3(G200), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n488), .A2(new_n509), .A3(new_n511), .A4(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n468), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n486), .B1(new_n485), .B2(new_n299), .ZN(new_n522));
  AOI211_X1 g0322(.A(KEYINPUT76), .B(new_n300), .C1(new_n479), .C2(new_n484), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n516), .A2(new_n354), .A3(new_n517), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(G169), .B2(new_n508), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n520), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT19), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n301), .B1(new_n258), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n481), .A2(new_n217), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n301), .B(G68), .C1(new_n255), .C2(new_n256), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n530), .B1(new_n330), .B2(new_n219), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n299), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n335), .A2(new_n329), .ZN(new_n538));
  INV_X1    g0338(.A(new_n329), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n296), .A2(new_n300), .A3(new_n539), .A4(new_n466), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n264), .A2(new_n362), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n513), .A2(G1698), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(new_n255), .C2(new_n256), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G116), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n252), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n218), .B1(new_n265), .B2(G45), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n252), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n252), .A2(G274), .ZN(new_n549));
  INV_X1    g0349(.A(new_n489), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n274), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n495), .A2(new_n489), .B1(new_n252), .B2(new_n547), .ZN(new_n553));
  NOR2_X1   g0353(.A1(G238), .A2(G1698), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n513), .B2(G1698), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n555), .A2(new_n347), .B1(G33), .B2(G116), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n354), .B(new_n553), .C1(new_n556), .C2(new_n252), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n541), .A2(new_n552), .A3(new_n557), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n536), .A2(new_n299), .B1(new_n335), .B2(new_n329), .ZN(new_n559));
  OAI21_X1  g0359(.A(G200), .B1(new_n546), .B2(new_n551), .ZN(new_n560));
  OAI211_X1 g0360(.A(G190), .B(new_n553), .C1(new_n556), .C2(new_n252), .ZN(new_n561));
  AOI211_X1 g0361(.A(new_n465), .B(new_n299), .C1(new_n289), .C2(new_n292), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(G87), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n559), .A2(new_n560), .A3(new_n561), .A4(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n492), .A2(G264), .A3(new_n252), .ZN(new_n566));
  INV_X1    g0366(.A(G294), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n306), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G250), .A2(G1698), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n569), .B1(new_n220), .B2(G1698), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n568), .B1(new_n570), .B2(new_n347), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n497), .B(new_n566), .C1(new_n571), .C2(new_n252), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n220), .A2(G1698), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G250), .B2(G1698), .ZN(new_n575));
  OAI22_X1  g0375(.A1(new_n575), .A2(new_n339), .B1(new_n306), .B2(new_n567), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n507), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT82), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n578), .A3(new_n497), .A4(new_n566), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(G169), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT83), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n572), .B2(new_n354), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n496), .A2(new_n489), .B1(new_n210), .B2(new_n251), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n576), .A2(new_n507), .B1(new_n583), .B2(G264), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT83), .A3(G179), .A4(new_n497), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n580), .A2(new_n582), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(G116), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n330), .A2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT23), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n301), .B2(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n340), .A2(KEYINPUT23), .A3(G20), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT22), .ZN(new_n593));
  AOI21_X1  g0393(.A(G20), .B1(new_n345), .B2(new_n346), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(G87), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n301), .B(G87), .C1(new_n255), .C2(new_n256), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(KEYINPUT22), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n592), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT24), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT24), .B(new_n592), .C1(new_n595), .C2(new_n597), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n600), .A2(new_n299), .A3(new_n601), .ZN(new_n602));
  XOR2_X1   g0402(.A(KEYINPUT81), .B(KEYINPUT25), .Z(new_n603));
  NAND3_X1  g0403(.A1(new_n335), .A2(new_n340), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(KEYINPUT81), .B(KEYINPUT25), .C1(new_n296), .C2(G107), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n605), .C1(new_n467), .C2(new_n340), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n586), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT84), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n300), .B1(new_n598), .B2(new_n599), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n606), .B1(new_n612), .B2(new_n601), .ZN(new_n613));
  AOI21_X1  g0413(.A(G190), .B1(new_n573), .B2(new_n579), .ZN(new_n614));
  AOI21_X1  g0414(.A(G200), .B1(new_n584), .B2(new_n497), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n586), .A2(KEYINPUT84), .A3(new_n608), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n611), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n297), .A2(new_n298), .B1(G20), .B2(new_n587), .ZN(new_n619));
  AOI21_X1  g0419(.A(G20), .B1(G33), .B2(G283), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n306), .A2(G97), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT80), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT80), .B1(new_n620), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n619), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT20), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(KEYINPUT20), .B(new_n619), .C1(new_n622), .C2(new_n623), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n296), .A2(G116), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n629), .B1(new_n562), .B2(G116), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n492), .A2(G270), .A3(new_n252), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n632), .A2(KEYINPUT78), .A3(new_n497), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT78), .B1(new_n632), .B2(new_n497), .ZN(new_n634));
  OAI211_X1 g0434(.A(G257), .B(new_n362), .C1(new_n255), .C2(new_n256), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n345), .A2(G303), .A3(new_n346), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT79), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n367), .A2(new_n638), .A3(G264), .ZN(new_n639));
  OAI211_X1 g0439(.A(G264), .B(G1698), .C1(new_n255), .C2(new_n256), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT79), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n637), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n633), .A2(new_n634), .B1(new_n642), .B2(new_n252), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n631), .A2(new_n643), .A3(KEYINPUT21), .A4(G169), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n632), .A2(new_n497), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT78), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n632), .A2(new_n497), .A3(KEYINPUT78), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n635), .A2(new_n636), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n638), .B1(new_n367), .B2(G264), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n640), .A2(KEYINPUT79), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n647), .A2(new_n648), .B1(new_n652), .B2(new_n507), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(G179), .A3(new_n631), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n644), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n631), .A2(new_n643), .A3(G169), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT21), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n647), .A2(new_n648), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n507), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(new_n452), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n628), .A2(new_n630), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n661), .B(new_n662), .C1(new_n318), .C2(new_n653), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n655), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n618), .A2(new_n664), .ZN(new_n665));
  AND4_X1   g0465(.A1(new_n463), .A2(new_n529), .A3(new_n565), .A4(new_n665), .ZN(G372));
  XNOR2_X1  g0466(.A(new_n446), .B(KEYINPUT18), .ZN(new_n667));
  INV_X1    g0467(.A(new_n356), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n327), .A2(new_n668), .B1(new_n286), .B2(new_n316), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n458), .A2(new_n459), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n667), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n399), .A2(new_n401), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n391), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n558), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n524), .A2(new_n565), .A3(new_n527), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n478), .A2(new_n487), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n526), .B1(new_n679), .B2(new_n521), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(KEYINPUT26), .A3(new_n565), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n675), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n585), .A2(new_n582), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n613), .B1(new_n683), .B2(new_n580), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n644), .A2(new_n654), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n274), .B1(new_n659), .B2(new_n660), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT21), .B1(new_n686), .B2(new_n631), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n520), .A2(new_n528), .A3(new_n565), .A4(new_n616), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n682), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n674), .B1(new_n462), .B2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n692), .B(KEYINPUT85), .Z(G369));
  NAND2_X1  g0493(.A1(new_n655), .A2(new_n658), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n265), .A2(new_n301), .A3(G13), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(KEYINPUT27), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT86), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G213), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n695), .B2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G343), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n694), .A2(new_n631), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n703), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n662), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n664), .B2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT87), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT87), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n611), .A2(new_n616), .A3(new_n617), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n613), .B2(new_n705), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n684), .A2(new_n703), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n710), .A2(G330), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n694), .A2(new_n705), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n716), .A2(new_n618), .B1(new_n609), .B2(new_n703), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(G399));
  NOR2_X1   g0519(.A1(new_n532), .A2(G116), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT88), .ZN(new_n721));
  INV_X1    g0521(.A(new_n207), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(new_n265), .ZN(new_n724));
  INV_X1    g0524(.A(new_n213), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n721), .A2(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n726), .B(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n659), .A2(new_n660), .A3(G179), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n546), .A2(new_n551), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n508), .A2(new_n731), .A3(new_n584), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n729), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT90), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n731), .A2(G179), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n643), .A2(new_n518), .A3(new_n572), .A4(new_n735), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n734), .B1(new_n733), .B2(new_n736), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n508), .A2(new_n731), .A3(new_n584), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(KEYINPUT30), .A3(G179), .A4(new_n653), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n737), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT31), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n705), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT91), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT91), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n733), .A2(new_n736), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n740), .B1(new_n748), .B2(new_n734), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n747), .B(new_n744), .C1(new_n749), .C2(new_n737), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n740), .A2(new_n733), .A3(new_n736), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n703), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n743), .ZN(new_n753));
  AND4_X1   g0553(.A1(new_n520), .A2(new_n528), .A3(new_n565), .A4(new_n705), .ZN(new_n754));
  AND4_X1   g0554(.A1(new_n658), .A2(new_n663), .A3(new_n654), .A4(new_n644), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n711), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n746), .A2(new_n750), .A3(new_n753), .A4(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(G330), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT29), .ZN(new_n759));
  AOI21_X1  g0559(.A(KEYINPUT84), .B1(new_n586), .B2(new_n608), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n586), .A2(KEYINPUT84), .A3(new_n608), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n694), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n682), .B1(new_n762), .B2(new_n689), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n759), .B1(new_n763), .B2(new_n705), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n690), .A2(new_n705), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(KEYINPUT29), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n758), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n728), .B1(new_n767), .B2(G1), .ZN(G364));
  INV_X1    g0568(.A(G330), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n708), .B2(new_n709), .ZN(new_n770));
  INV_X1    g0570(.A(G13), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n265), .B1(new_n772), .B2(G45), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n723), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G330), .B2(new_n710), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n775), .B(KEYINPUT93), .Z(new_n779));
  NAND2_X1  g0579(.A1(new_n347), .A2(new_n207), .ZN(new_n780));
  INV_X1    g0580(.A(G355), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n780), .A2(new_n781), .B1(G116), .B2(new_n207), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n722), .A2(new_n347), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n214), .B2(new_n261), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n243), .A2(new_n261), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(G13), .A2(G33), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n298), .B1(G20), .B2(new_n274), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n779), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n301), .A2(new_n354), .A3(G200), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n452), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n322), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n301), .ZN(new_n799));
  OAI22_X1  g0599(.A1(new_n797), .A2(new_n380), .B1(new_n219), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n301), .A2(new_n354), .A3(new_n318), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n452), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n800), .B1(G50), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n301), .A2(G179), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n805), .A2(new_n322), .A3(new_n318), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(new_n406), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n805), .A2(G190), .A3(G200), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n809), .A2(new_n217), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n801), .A2(new_n322), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n347), .B1(new_n811), .B2(new_n290), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n805), .A2(new_n322), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n810), .B(new_n812), .C1(G107), .C2(new_n814), .ZN(new_n815));
  AND3_X1   g0615(.A1(new_n795), .A2(KEYINPUT94), .A3(new_n322), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT94), .B1(new_n795), .B2(new_n322), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G77), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n804), .A2(new_n808), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G322), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n797), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n806), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n347), .B(new_n823), .C1(G329), .C2(new_n824), .ZN(new_n825));
  XOR2_X1   g0625(.A(KEYINPUT33), .B(G317), .Z(new_n826));
  OAI22_X1  g0626(.A1(new_n811), .A2(new_n826), .B1(new_n799), .B2(new_n567), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(G326), .B2(new_n803), .ZN(new_n828));
  INV_X1    g0628(.A(new_n809), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n829), .A2(G303), .B1(new_n814), .B2(G283), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n825), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n818), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n821), .B1(new_n831), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n794), .B1(new_n834), .B2(new_n791), .ZN(new_n835));
  INV_X1    g0635(.A(new_n790), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n835), .B1(new_n710), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT95), .Z(new_n838));
  NAND2_X1  g0638(.A1(new_n777), .A2(KEYINPUT92), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n778), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  INV_X1    g0641(.A(new_n779), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n791), .A2(new_n788), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(new_n336), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n811), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n803), .A2(G137), .B1(new_n845), .B2(G150), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n797), .C1(new_n818), .C2(new_n406), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT98), .Z(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  OR2_X1    g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n813), .A2(new_n290), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n339), .B(new_n852), .C1(G132), .C2(new_n824), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n202), .B2(new_n809), .C1(new_n380), .C2(new_n799), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n849), .B2(new_n850), .ZN(new_n855));
  INV_X1    g0655(.A(G283), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n818), .A2(new_n587), .B1(new_n856), .B2(new_n811), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n857), .A2(KEYINPUT96), .B1(G303), .B2(new_n803), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(KEYINPUT96), .B2(new_n857), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT97), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n217), .A2(new_n813), .B1(new_n809), .B2(new_n340), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n339), .B1(new_n806), .B2(new_n832), .C1(new_n799), .C2(new_n219), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n861), .B(new_n862), .C1(G294), .C2(new_n796), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n851), .A2(new_n855), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n791), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n844), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT99), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(KEYINPUT99), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n703), .A2(new_n338), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n356), .A3(new_n360), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n356), .A2(new_n869), .A3(new_n360), .A4(KEYINPUT100), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(new_n356), .C2(new_n705), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n867), .B(new_n868), .C1(new_n789), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n873), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n705), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n689), .A2(new_n688), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT26), .B1(new_n680), .B2(new_n565), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n558), .A2(new_n564), .ZN(new_n881));
  NOR4_X1   g0681(.A1(new_n488), .A2(new_n881), .A3(new_n526), .A4(new_n677), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n558), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n878), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT101), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n690), .A2(KEYINPUT101), .A3(new_n878), .ZN(new_n887));
  INV_X1    g0687(.A(new_n874), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n886), .A2(new_n887), .B1(new_n765), .B2(new_n888), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n758), .A2(new_n889), .B1(new_n723), .B2(new_n774), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n758), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n875), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT102), .Z(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(G384));
  AOI211_X1 g0694(.A(new_n587), .B(new_n211), .C1(new_n483), .C2(KEYINPUT35), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(KEYINPUT35), .B2(new_n483), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT36), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n336), .B(new_n213), .C1(new_n413), .C2(G68), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n290), .A2(G50), .ZN(new_n899));
  OAI211_X1 g0699(.A(G1), .B(new_n771), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT103), .Z(new_n902));
  INV_X1    g0702(.A(KEYINPUT106), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n445), .A2(new_n404), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n436), .ZN(new_n906));
  INV_X1    g0706(.A(new_n701), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n906), .A2(new_n908), .A3(new_n456), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n906), .A2(new_n908), .A3(new_n911), .A4(new_n456), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n908), .B1(new_n667), .B2(new_n670), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n904), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT104), .B1(new_n415), .B2(new_n420), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT104), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n441), .A2(new_n443), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n916), .A2(new_n918), .A3(new_n423), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n405), .B1(new_n919), .B2(new_n422), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n456), .B1(new_n920), .B2(new_n437), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n701), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT37), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n912), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n460), .A2(new_n922), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n924), .A2(new_n925), .A3(KEYINPUT38), .ZN(new_n926));
  XNOR2_X1  g0726(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n915), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  AND4_X1   g0729(.A1(new_n911), .A2(new_n906), .A3(new_n908), .A4(new_n456), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n444), .A2(new_n299), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n441), .A2(new_n443), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT16), .B1(new_n932), .B2(KEYINPUT104), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n931), .B1(new_n933), .B2(new_n918), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n907), .B1(new_n934), .B2(new_n405), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n436), .B1(new_n934), .B2(new_n405), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n456), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n930), .B1(KEYINPUT37), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n935), .B1(new_n667), .B2(new_n670), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n904), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n929), .B1(new_n940), .B2(new_n926), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n903), .B1(new_n928), .B2(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n924), .A2(KEYINPUT38), .A3(new_n925), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n924), .B2(new_n925), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT39), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n915), .A2(new_n926), .A3(new_n927), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n317), .A2(new_n703), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n667), .A2(new_n907), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n356), .A2(new_n703), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n886), .B2(new_n887), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n316), .B(new_n703), .C1(new_n286), .C2(new_n326), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n313), .A2(new_n315), .A3(new_n703), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n956), .B(new_n326), .C1(new_n286), .C2(new_n316), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n940), .A2(new_n926), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n951), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n950), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n463), .B1(new_n766), .B2(new_n764), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n674), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n962), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n752), .A2(KEYINPUT107), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT107), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n751), .A2(new_n967), .A3(new_n703), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n966), .A2(new_n743), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n751), .A2(new_n744), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n756), .A3(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n956), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n317), .A2(new_n327), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n888), .B1(new_n973), .B2(new_n954), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n460), .A2(new_n905), .A3(new_n907), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n910), .A2(new_n912), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT38), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n943), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(KEYINPUT40), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n874), .B1(new_n955), .B2(new_n957), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n665), .A2(new_n754), .B1(new_n744), .B2(new_n751), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n981), .B1(new_n982), .B2(new_n969), .ZN(new_n983));
  AOI21_X1  g0783(.A(KEYINPUT40), .B1(new_n940), .B2(new_n926), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n980), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n462), .B1(new_n969), .B2(new_n982), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n769), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n965), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n265), .B2(new_n772), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n965), .A2(new_n989), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n902), .B1(new_n991), .B2(new_n992), .ZN(G367));
  NAND2_X1  g0793(.A1(new_n559), .A2(new_n563), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n703), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n565), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n558), .B2(new_n995), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT109), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n529), .B1(new_n488), .B2(new_n705), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n680), .A2(new_n703), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n999), .B1(new_n715), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT108), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n770), .A2(KEYINPUT109), .A3(new_n714), .A4(new_n1005), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1004), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n998), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT108), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n998), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n716), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1005), .A2(new_n711), .A3(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n761), .A2(new_n760), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n528), .B1(new_n1000), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1017), .A2(KEYINPUT42), .B1(new_n1019), .B2(new_n705), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(KEYINPUT42), .B2(new_n1017), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1009), .A2(new_n1014), .A3(new_n1023), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n723), .B(KEYINPUT41), .Z(new_n1027));
  INV_X1    g0827(.A(KEYINPUT45), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n1002), .B2(new_n717), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n718), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT44), .B1(new_n1002), .B2(new_n717), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1002), .A2(KEYINPUT44), .A3(new_n717), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n715), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1016), .A2(new_n711), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n714), .B2(new_n1016), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n770), .B(new_n1038), .ZN(new_n1039));
  OAI211_X1 g0839(.A(new_n715), .B(new_n1031), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .A4(new_n767), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1027), .B1(new_n1041), .B2(new_n767), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT110), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n773), .B1(new_n1042), .B2(KEYINPUT110), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1025), .B(new_n1026), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n234), .A2(new_n784), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n793), .B1(new_n722), .B2(new_n539), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n842), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n811), .A2(new_n567), .B1(new_n799), .B2(new_n340), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n802), .A2(new_n832), .B1(new_n219), .B2(new_n813), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n819), .C2(G283), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n829), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1052));
  INV_X1    g0852(.A(G303), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n797), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(KEYINPUT46), .B1(new_n829), .B2(G116), .ZN(new_n1055));
  INV_X1    g0855(.A(G317), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n339), .B1(new_n806), .B2(new_n1056), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1051), .A2(new_n1052), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n818), .A2(new_n202), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n813), .A2(new_n336), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n799), .A2(new_n290), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(new_n413), .C2(new_n829), .ZN(new_n1063));
  INV_X1    g0863(.A(G137), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n347), .B1(new_n806), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G159), .B2(new_n845), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G143), .A2(new_n803), .B1(new_n796), .B2(G150), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1059), .B1(new_n1060), .B2(new_n1068), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT47), .Z(new_n1070));
  OAI221_X1 g0870(.A(new_n1048), .B1(new_n836), .B2(new_n997), .C1(new_n1070), .C2(new_n865), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1045), .A2(new_n1071), .ZN(G387));
  NAND3_X1  g0872(.A1(new_n712), .A2(new_n713), .A3(new_n790), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n783), .B1(new_n239), .B2(new_n261), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n721), .B2(new_n780), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n261), .B1(new_n290), .B2(new_n336), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n331), .A2(G50), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n721), .B(new_n1078), .C1(KEYINPUT50), .C2(new_n1077), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1075), .A2(new_n1079), .B1(new_n340), .B2(new_n722), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n779), .B1(new_n1080), .B2(new_n793), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n796), .A2(G317), .B1(new_n845), .B2(G311), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n1053), .B2(new_n818), .C1(new_n822), .C2(new_n802), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT48), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n799), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(G283), .B1(new_n829), .B2(G294), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT49), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n813), .A2(new_n587), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n347), .B(new_n1093), .C1(G326), .C2(new_n824), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n809), .A2(new_n336), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n797), .A2(new_n202), .B1(new_n406), .B2(new_n802), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n539), .C2(new_n1087), .ZN(new_n1098));
  INV_X1    g0898(.A(G150), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n347), .B1(new_n806), .B2(new_n1099), .C1(new_n219), .C2(new_n813), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n378), .B1(new_n413), .B2(KEYINPUT8), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n1101), .B2(new_n845), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1098), .B(new_n1102), .C1(new_n290), .C2(new_n818), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1081), .B1(new_n1104), .B2(new_n791), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1039), .A2(new_n774), .B1(new_n1073), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1039), .A2(new_n767), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n723), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1039), .A2(new_n767), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(G393));
  INV_X1    g0910(.A(KEYINPUT111), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1036), .A2(new_n1040), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT111), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1107), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT113), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1112), .A2(new_n1117), .A3(new_n1107), .A4(new_n1113), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1041), .A2(new_n723), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1114), .A2(new_n774), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n792), .B1(new_n219), .B2(new_n207), .C1(new_n246), .C2(new_n784), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n779), .A2(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G317), .A2(new_n803), .B1(new_n796), .B2(G311), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n811), .A2(new_n1053), .B1(new_n856), .B2(new_n809), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n339), .B1(new_n806), .B2(new_n822), .C1(new_n340), .C2(new_n813), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(G116), .C2(new_n1087), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n567), .B2(new_n818), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n811), .A2(new_n202), .B1(new_n290), .B2(new_n809), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n347), .B1(new_n806), .B2(new_n847), .C1(new_n217), .C2(new_n813), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(G77), .C2(new_n1087), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n331), .B2(new_n818), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G150), .A2(new_n803), .B1(new_n796), .B2(G159), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT51), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n1126), .A2(new_n1130), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g0937(.A(new_n1137), .B(KEYINPUT112), .Z(new_n1138));
  OAI221_X1 g0938(.A(new_n1124), .B1(new_n1005), .B2(new_n836), .C1(new_n865), .C2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1121), .A2(new_n1122), .A3(new_n1139), .ZN(G390));
  NAND3_X1  g0940(.A1(new_n757), .A2(G330), .A3(new_n874), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n958), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n971), .A2(G330), .A3(new_n974), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n884), .A2(new_n885), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT101), .B1(new_n690), .B2(new_n878), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n1146), .B1(new_n356), .B2(new_n703), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1018), .A2(new_n616), .A3(new_n755), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n520), .A2(new_n528), .A3(new_n565), .A4(new_n705), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n970), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n751), .A2(new_n967), .A3(new_n703), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n967), .B1(new_n751), .B2(new_n703), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1152), .A2(new_n1153), .A3(KEYINPUT31), .ZN(new_n1154));
  OAI211_X1 g0954(.A(G330), .B(new_n874), .C1(new_n1151), .C2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n958), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT114), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(KEYINPUT114), .A3(new_n958), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n952), .B1(new_n763), .B2(new_n878), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n757), .A2(G330), .A3(new_n974), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1148), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n463), .A2(G330), .A3(new_n971), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n963), .A2(new_n674), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n949), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n953), .B2(new_n958), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1169), .A2(new_n942), .A3(new_n947), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1160), .A2(new_n958), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n915), .A2(new_n926), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1168), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1170), .A2(new_n1161), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1143), .B1(new_n1170), .B2(new_n1175), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1167), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1165), .B1(new_n1148), .B2(new_n1162), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n958), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n949), .B1(new_n1147), .B2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1161), .B(new_n1175), .C1(new_n948), .C2(new_n1181), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n945), .A2(KEYINPUT106), .A3(new_n946), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT106), .B1(new_n945), .B2(new_n946), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1174), .B1(new_n1185), .B2(new_n1169), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1179), .B(new_n1182), .C1(new_n1143), .C2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1178), .A2(new_n1187), .A3(new_n723), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1182), .B(new_n774), .C1(new_n1186), .C2(new_n1143), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT116), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n843), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n779), .B1(new_n1101), .B2(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n811), .A2(new_n340), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n852), .B(new_n1193), .C1(G283), .C2(new_n803), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n347), .B(new_n810), .C1(G294), .C2(new_n824), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1194), .B(new_n1195), .C1(new_n219), .C2(new_n818), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n796), .A2(G116), .B1(new_n1087), .B2(G77), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT115), .Z(new_n1198));
  AOI22_X1  g0998(.A1(new_n803), .A2(G128), .B1(G159), .B2(new_n1087), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n796), .A2(G132), .B1(new_n845), .B2(G137), .ZN(new_n1200));
  INV_X1    g1000(.A(G125), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n347), .B1(new_n806), .B2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G50), .B2(new_n814), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1199), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n809), .A2(new_n1099), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT53), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(KEYINPUT54), .B(G143), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1206), .B1(new_n818), .B2(new_n1207), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n1196), .A2(new_n1198), .B1(new_n1204), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1192), .B1(new_n1209), .B2(new_n791), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n948), .B2(new_n789), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1189), .A2(new_n1190), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1190), .B1(new_n1189), .B2(new_n1211), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1188), .B1(new_n1212), .B2(new_n1213), .ZN(G378));
  OAI21_X1  g1014(.A(new_n775), .B1(G50), .B2(new_n1191), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n673), .A2(new_n390), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n701), .B1(new_n375), .B2(new_n384), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n402), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g1020(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1221), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n402), .A2(new_n1219), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n1217), .B(new_n391), .C1(new_n399), .C2(new_n401), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1223), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1222), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1228), .A2(new_n789), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n797), .A2(new_n340), .B1(new_n587), .B2(new_n802), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(G97), .B2(new_n845), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n260), .B(new_n339), .C1(new_n806), .C2(new_n856), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n813), .A2(new_n380), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(new_n1062), .A3(new_n1096), .A4(new_n1233), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1231), .B(new_n1234), .C1(new_n329), .C2(new_n818), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT58), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(G50), .B1(new_n306), .B2(new_n260), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1238), .B1(new_n347), .B2(G41), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G128), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n797), .A2(new_n1241), .B1(new_n1201), .B2(new_n802), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G132), .B2(new_n845), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1207), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1087), .A2(G150), .B1(new_n829), .B2(new_n1244), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1243), .B(new_n1245), .C1(new_n1064), .C2(new_n818), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(new_n1246), .B(KEYINPUT117), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n814), .A2(G159), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G33), .B(G41), .C1(new_n824), .C2(G124), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n1248), .A2(KEYINPUT59), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1240), .B1(new_n1236), .B2(new_n1235), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1215), .B(new_n1229), .C1(new_n1254), .C2(new_n791), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT118), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1228), .B1(new_n986), .B2(G330), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n769), .B(new_n1227), .C1(new_n980), .C2(new_n985), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1256), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n950), .A2(new_n961), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1172), .A2(new_n971), .A3(new_n974), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n1262), .A2(KEYINPUT40), .B1(new_n984), .B2(new_n983), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1227), .B1(new_n1263), .B2(new_n769), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n986), .A2(G330), .A3(new_n1228), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1266), .A2(new_n962), .A3(new_n1256), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1261), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1255), .B1(new_n1268), .B2(new_n774), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1165), .B1(new_n1270), .B2(new_n1179), .ZN(new_n1271));
  AND4_X1   g1071(.A1(new_n950), .A2(new_n1264), .A3(new_n961), .A4(new_n1265), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1264), .A2(new_n1265), .B1(new_n950), .B2(new_n961), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT57), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n723), .B1(new_n1271), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1187), .A2(new_n1166), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT57), .B1(new_n1276), .B2(new_n1268), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1269), .B1(new_n1275), .B2(new_n1277), .ZN(G375));
  NAND2_X1  g1078(.A1(new_n1163), .A2(new_n774), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n842), .B1(new_n290), .B2(new_n843), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n797), .A2(new_n1064), .B1(new_n202), .B2(new_n799), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G159), .B2(new_n829), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n819), .A2(G150), .ZN(new_n1283));
  OAI221_X1 g1083(.A(new_n347), .B1(new_n806), .B2(new_n1241), .C1(new_n380), .C2(new_n813), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n803), .A2(G132), .B1(new_n845), .B2(new_n1244), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1282), .A2(new_n1283), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n797), .A2(new_n856), .B1(new_n219), .B2(new_n809), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G294), .B2(new_n803), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n347), .B(new_n1061), .C1(G303), .C2(new_n824), .ZN(new_n1290));
  AOI22_X1  g1090(.A1(new_n845), .A2(G116), .B1(new_n1087), .B2(new_n539), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n818), .A2(new_n340), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1287), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n1294), .A2(KEYINPUT119), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(KEYINPUT119), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n791), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1280), .B1(new_n1295), .B2(new_n1297), .C1(new_n1180), .C2(new_n789), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1279), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1027), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1148), .A2(new_n1162), .A3(new_n1165), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1167), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(G381));
  OR3_X1    g1104(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1305));
  NOR4_X1   g1105(.A1(G387), .A2(new_n1305), .A3(G390), .A4(G381), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1189), .A2(new_n1211), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1188), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  OR2_X1    g1109(.A1(new_n1309), .A2(G375), .ZN(G407));
  NOR2_X1   g1110(.A1(new_n699), .A2(G343), .ZN(new_n1311));
  XOR2_X1   g1111(.A(new_n1311), .B(KEYINPUT120), .Z(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G407), .B(G213), .C1(G375), .C2(new_n1313), .ZN(G409));
  AND3_X1   g1114(.A1(new_n1121), .A2(new_n1122), .A3(new_n1139), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(G387), .A2(new_n1315), .ZN(new_n1316));
  XNOR2_X1  g1116(.A(new_n840), .B(G393), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(G390), .A2(new_n1045), .A3(new_n1071), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1320));
  OR2_X1    g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT61), .ZN(new_n1322));
  OAI211_X1 g1122(.A(G378), .B(new_n1269), .C1(new_n1275), .C2(new_n1277), .ZN(new_n1323));
  AND3_X1   g1123(.A1(new_n1276), .A2(new_n1301), .A3(new_n1268), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n774), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1215), .B1(new_n1254), .B2(new_n791), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n789), .B2(new_n1228), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(new_n1308), .B1(new_n1324), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1323), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(KEYINPUT121), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1311), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT121), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1323), .A2(new_n1329), .A3(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1148), .A2(new_n1162), .A3(KEYINPUT60), .A4(new_n1165), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n723), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1167), .A2(KEYINPUT60), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1336), .B1(new_n1337), .B2(new_n1302), .ZN(new_n1338));
  OAI21_X1  g1138(.A(G384), .B1(new_n1338), .B2(new_n1299), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1302), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1340), .B1(KEYINPUT60), .B2(new_n1167), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n893), .B(new_n1300), .C1(new_n1341), .C2(new_n1336), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1331), .A2(new_n1332), .A3(new_n1334), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT125), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1312), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1330), .B2(new_n1346), .ZN(new_n1347));
  AOI211_X1 g1147(.A(KEYINPUT125), .B(new_n1312), .C1(new_n1323), .C2(new_n1329), .ZN(new_n1348));
  OR2_X1    g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT122), .ZN(new_n1350));
  INV_X1    g1150(.A(G2897), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1332), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1352), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1343), .A2(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1354), .A2(KEYINPUT123), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT123), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1343), .A2(new_n1356), .A3(new_n1353), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1355), .A2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1343), .ZN(new_n1359));
  NOR2_X1   g1159(.A1(new_n1346), .A2(new_n1351), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1358), .A2(new_n1361), .ZN(new_n1362));
  OAI221_X1 g1162(.A(new_n1322), .B1(new_n1344), .B2(KEYINPUT62), .C1(new_n1349), .C2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT62), .ZN(new_n1364));
  AOI21_X1  g1164(.A(new_n1364), .B1(new_n1349), .B2(new_n1343), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1321), .B1(new_n1363), .B2(new_n1365), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1331), .A2(new_n1332), .A3(new_n1334), .ZN(new_n1367));
  INV_X1    g1167(.A(KEYINPUT124), .ZN(new_n1368));
  AOI22_X1  g1168(.A1(new_n1355), .A2(new_n1357), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1367), .A2(new_n1368), .A3(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1368), .B1(new_n1367), .B2(new_n1369), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1370), .A2(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT63), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1344), .A2(new_n1373), .ZN(new_n1374));
  NOR3_X1   g1174(.A1(new_n1319), .A2(new_n1320), .A3(KEYINPUT61), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1359), .A2(new_n1373), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1376), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1377));
  NAND3_X1  g1177(.A1(new_n1374), .A2(new_n1375), .A3(new_n1377), .ZN(new_n1378));
  NOR3_X1   g1178(.A1(new_n1372), .A2(KEYINPUT126), .A3(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT126), .ZN(new_n1380));
  AND3_X1   g1180(.A1(new_n1374), .A2(new_n1377), .A3(new_n1375), .ZN(new_n1381));
  AND3_X1   g1181(.A1(new_n1323), .A2(new_n1329), .A3(new_n1333), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1333), .B1(new_n1323), .B2(new_n1329), .ZN(new_n1383));
  NOR3_X1   g1183(.A1(new_n1382), .A2(new_n1383), .A3(new_n1311), .ZN(new_n1384));
  OAI21_X1  g1184(.A(KEYINPUT124), .B1(new_n1384), .B2(new_n1362), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1367), .A2(new_n1368), .A3(new_n1369), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1380), .B1(new_n1381), .B2(new_n1387), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1366), .B1(new_n1379), .B2(new_n1388), .ZN(G405));
  OR2_X1    g1189(.A1(new_n1321), .A2(new_n1359), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1321), .A2(new_n1359), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1392));
  AND2_X1   g1192(.A1(G375), .A2(new_n1308), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1393), .A2(new_n1394), .ZN(new_n1395));
  INV_X1    g1195(.A(KEYINPUT127), .ZN(new_n1396));
  AOI21_X1  g1196(.A(new_n1395), .B1(new_n1396), .B2(new_n1393), .ZN(new_n1397));
  INV_X1    g1197(.A(new_n1397), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1392), .A2(new_n1398), .ZN(new_n1399));
  NAND3_X1  g1199(.A1(new_n1390), .A2(new_n1397), .A3(new_n1391), .ZN(new_n1400));
  NAND2_X1  g1200(.A1(new_n1399), .A2(new_n1400), .ZN(G402));
endmodule


