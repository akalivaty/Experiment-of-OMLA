//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1266, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G58), .A2(G232), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n210), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(G20), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n213), .B1(KEYINPUT1), .B2(new_n222), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n222), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n232), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G50), .B(G68), .Z(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(G1), .A2(G13), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT8), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n252), .A2(new_n254), .B1(G20), .B2(new_n204), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n208), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT67), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n257), .B1(G20), .B2(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G150), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n248), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT68), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n246), .A3(new_n245), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n207), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  OAI22_X1  g0066(.A1(new_n264), .A2(new_n266), .B1(G50), .B2(new_n263), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT69), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G222), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(G223), .A3(G1698), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n272), .B(new_n273), .C1(new_n214), .C2(new_n270), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n246), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n223), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n279), .A2(G274), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G41), .A2(G45), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G1), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n207), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n207), .A2(new_n288), .B1(new_n223), .B2(new_n278), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n280), .A2(new_n285), .B1(new_n289), .B2(G226), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n276), .A2(new_n277), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n276), .A2(new_n290), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n269), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n269), .A2(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n262), .A2(new_n298), .A3(new_n268), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n292), .A2(G200), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n276), .A2(G190), .A3(new_n290), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n296), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n262), .A2(new_n298), .A3(new_n268), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n298), .B1(new_n262), .B2(new_n268), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n304), .B(new_n296), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n295), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n263), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n214), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT70), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n259), .A2(new_n252), .ZN(new_n314));
  INV_X1    g0114(.A(new_n254), .ZN(new_n315));
  XNOR2_X1  g0115(.A(KEYINPUT15), .B(G87), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n315), .A2(new_n316), .B1(new_n214), .B2(new_n208), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n247), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n265), .A2(G77), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n264), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(KEYINPUT71), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n264), .A2(new_n322), .A3(new_n319), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n313), .B(new_n318), .C1(new_n321), .C2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT72), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n270), .A2(G232), .A3(new_n271), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n270), .A2(G238), .A3(G1698), .ZN(new_n328));
  INV_X1    g0128(.A(G107), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n270), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n275), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n280), .A2(new_n285), .B1(new_n289), .B2(G244), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G200), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n331), .A2(G190), .A3(new_n332), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n324), .A2(new_n325), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n326), .A2(new_n334), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n333), .A2(new_n293), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n324), .C1(G179), .C2(new_n333), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n310), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT77), .ZN(new_n343));
  XNOR2_X1  g0143(.A(new_n342), .B(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT3), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G33), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n345), .A2(new_n347), .A3(G226), .A4(G1698), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n345), .A2(new_n347), .A3(G223), .A4(new_n271), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n344), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n275), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n280), .A2(new_n285), .B1(new_n289), .B2(G232), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(KEYINPUT78), .A3(G179), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT78), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n351), .A2(new_n352), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n355), .B1(new_n356), .B2(new_n277), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n293), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n252), .A2(new_n265), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n360), .A2(new_n264), .B1(new_n263), .B2(new_n252), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n361), .B(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n270), .B2(G20), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n346), .A2(G33), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT7), .B(new_n208), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n203), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT74), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(KEYINPUT74), .A2(G58), .A3(G68), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n225), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G20), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n259), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT75), .B1(new_n369), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n248), .B1(new_n378), .B2(KEYINPUT16), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT16), .ZN(new_n380));
  OAI211_X1 g0180(.A(KEYINPUT75), .B(new_n380), .C1(new_n369), .C2(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n363), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT18), .B1(new_n359), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(new_n381), .A3(new_n247), .ZN(new_n385));
  INV_X1    g0185(.A(new_n363), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n356), .A2(new_n355), .A3(new_n277), .ZN(new_n389));
  INV_X1    g0189(.A(new_n358), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT78), .B1(new_n353), .B2(G179), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G200), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n353), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(G190), .B2(new_n353), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n385), .A2(new_n386), .A3(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT17), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n382), .A2(KEYINPUT17), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n395), .A2(new_n404), .A3(KEYINPUT79), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n383), .A2(new_n393), .A3(new_n401), .A4(new_n402), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT79), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n270), .A2(G232), .A3(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n345), .A2(new_n347), .A3(G226), .A4(new_n271), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n275), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n280), .A2(new_n285), .B1(new_n289), .B2(G238), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n414), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n413), .A2(new_n415), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G190), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n259), .A2(G50), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n254), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n248), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT11), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT12), .B1(new_n263), .B2(G68), .ZN(new_n427));
  OR3_X1    g0227(.A1(new_n263), .A2(KEYINPUT12), .A3(G68), .ZN(new_n428));
  INV_X1    g0228(.A(new_n264), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n203), .B1(new_n207), .B2(G20), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n427), .A2(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n425), .A2(KEYINPUT11), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n418), .A2(new_n422), .A3(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n420), .A2(G179), .A3(new_n421), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT14), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(G169), .C1(new_n416), .C2(new_n417), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT73), .ZN(new_n442));
  INV_X1    g0242(.A(new_n432), .ZN(new_n443));
  INV_X1    g0243(.A(new_n433), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n432), .A2(KEYINPUT73), .A3(new_n433), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n435), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n341), .A2(new_n405), .A3(new_n408), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n345), .A2(new_n347), .A3(G244), .A4(new_n271), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT4), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(G283), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n253), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G250), .A2(G1698), .ZN(new_n456));
  NAND2_X1  g0256(.A1(KEYINPUT4), .A2(G244), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G1698), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n270), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n275), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n287), .A2(G1), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G257), .A3(new_n279), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT5), .B(G41), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n467), .A2(new_n279), .A3(G274), .A4(new_n462), .ZN(new_n468));
  AND2_X1   g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n461), .A2(G190), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n396), .B1(new_n461), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(KEYINPUT81), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT80), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n270), .A2(new_n364), .A3(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n345), .A2(new_n347), .ZN(new_n475));
  AOI21_X1  g0275(.A(KEYINPUT7), .B1(new_n475), .B2(new_n208), .ZN(new_n476));
  OAI21_X1  g0276(.A(G107), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT6), .ZN(new_n478));
  AND2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n329), .A2(KEYINPUT6), .A3(G97), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n483), .A2(G20), .B1(G77), .B2(new_n259), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n248), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n263), .A2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n207), .A2(G33), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n263), .A2(new_n487), .A3(new_n246), .A4(new_n245), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n486), .B1(new_n489), .B2(G97), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n473), .B1(new_n485), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n483), .A2(G20), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n259), .A2(G77), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n329), .B1(new_n365), .B2(new_n368), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n247), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(KEYINPUT80), .A3(new_n490), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT81), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n461), .A2(new_n469), .A3(new_n499), .A4(G190), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n472), .A2(new_n492), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n461), .A2(new_n469), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G169), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n461), .A2(G179), .A3(new_n469), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n497), .A2(new_n490), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT82), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n508), .A2(G116), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(KEYINPUT82), .ZN(new_n511));
  OAI21_X1  g0311(.A(G33), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n345), .A2(new_n347), .A3(G244), .A4(G1698), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n345), .A2(new_n347), .A3(G238), .A4(new_n271), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n275), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n279), .A2(G274), .A3(new_n462), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n207), .A2(G45), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n279), .A2(G250), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n516), .A2(new_n277), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(G169), .B1(new_n516), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n208), .ZN(new_n526));
  INV_X1    g0326(.A(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n480), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT83), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n528), .A3(KEYINPUT83), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT19), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n533), .B1(new_n315), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n270), .A2(new_n208), .A3(G68), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n532), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n247), .ZN(new_n538));
  INV_X1    g0338(.A(new_n316), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n263), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n489), .A2(new_n539), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G190), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n516), .A2(new_n521), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n520), .B1(new_n275), .B2(new_n515), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(G200), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n488), .A2(new_n527), .ZN(new_n548));
  AOI211_X1 g0348(.A(new_n540), .B(new_n548), .C1(new_n537), .C2(new_n247), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n524), .A2(new_n543), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n501), .A2(new_n507), .A3(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n345), .A2(new_n347), .A3(G257), .A4(G1698), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n345), .A2(new_n347), .A3(G250), .A4(new_n271), .ZN(new_n553));
  NAND2_X1  g0353(.A1(G33), .A2(G294), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n275), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n275), .B1(new_n462), .B2(new_n467), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G264), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n558), .A3(new_n468), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n396), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n555), .A2(new_n275), .B1(new_n557), .B2(G264), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n544), .A3(new_n468), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n345), .A2(new_n347), .A3(new_n208), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n270), .A2(new_n566), .A3(new_n208), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT24), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n510), .A2(KEYINPUT82), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n508), .A2(G116), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n253), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n208), .B2(G107), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n329), .A2(KEYINPUT23), .A3(G20), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n572), .A2(new_n208), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n569), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n569), .B1(new_n568), .B2(new_n576), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n247), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT25), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n263), .B2(G107), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n263), .A2(new_n581), .A3(G107), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n583), .A2(new_n584), .B1(new_n329), .B2(new_n488), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n563), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n559), .A2(new_n293), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n561), .A2(new_n277), .A3(new_n468), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n580), .B2(new_n586), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G20), .B1(G33), .B2(G283), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n253), .A2(G97), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n594), .A2(new_n595), .B1(new_n245), .B2(new_n246), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n570), .A2(new_n571), .A3(G20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT20), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n597), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n570), .A2(new_n571), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n488), .A2(new_n510), .B1(new_n263), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n293), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n270), .A2(G264), .A3(G1698), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n270), .A2(G257), .A3(new_n271), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n475), .A2(G303), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n275), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n465), .A2(G270), .A3(new_n279), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n468), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT84), .B1(new_n612), .B2(new_n468), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n606), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n601), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT20), .B1(new_n596), .B2(new_n597), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n605), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n611), .B(G190), .C1(new_n613), .C2(new_n614), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n612), .A2(new_n468), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT84), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n612), .A2(KEYINPUT84), .A3(new_n468), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n275), .B2(new_n610), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n622), .B(new_n623), .C1(new_n628), .C2(new_n396), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n626), .A2(new_n627), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(G179), .A3(new_n611), .A4(new_n621), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n606), .A2(new_n615), .A3(KEYINPUT21), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n618), .A2(new_n629), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n450), .A2(new_n551), .A3(new_n593), .A4(new_n634), .ZN(G372));
  INV_X1    g0435(.A(new_n295), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n440), .A2(new_n438), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n420), .A2(new_n421), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n439), .B1(new_n638), .B2(G169), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n447), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n435), .B2(new_n339), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n404), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n395), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n304), .B1(new_n306), .B2(new_n307), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(KEYINPUT10), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n308), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n636), .B1(new_n643), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n546), .A2(new_n277), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n516), .A2(new_n521), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n293), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n543), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n632), .A2(new_n631), .ZN(new_n653));
  AOI21_X1  g0453(.A(KEYINPUT21), .B1(new_n606), .B2(new_n615), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n568), .A2(new_n576), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(KEYINPUT24), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n248), .B1(new_n657), .B2(new_n577), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n590), .B(new_n589), .C1(new_n658), .C2(new_n585), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n588), .B1(new_n655), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n652), .B1(new_n660), .B2(new_n551), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n492), .A2(new_n498), .B1(new_n503), .B2(new_n504), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT26), .B1(new_n662), .B2(new_n550), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n547), .A2(new_n549), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n651), .A3(new_n505), .A4(new_n506), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n647), .B1(new_n449), .B2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(G13), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n672), .A2(G1), .A3(G20), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT85), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n674), .B2(KEYINPUT27), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT27), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n673), .A2(KEYINPUT85), .A3(new_n677), .ZN(new_n678));
  OAI221_X1 g0478(.A(G213), .B1(KEYINPUT27), .B2(new_n674), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n622), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n633), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n618), .A2(new_n631), .A3(new_n632), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n682), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G330), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT86), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n681), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n658), .B2(new_n585), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n593), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n592), .A2(new_n690), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n659), .A2(new_n587), .A3(new_n681), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n684), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n698), .B1(new_n592), .B2(new_n681), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n211), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n528), .A2(G116), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G1), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n226), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n666), .A2(new_n651), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n507), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT90), .B1(new_n709), .B2(KEYINPUT26), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n662), .A2(new_n550), .A3(KEYINPUT26), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT90), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n667), .A2(new_n712), .A3(new_n665), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n690), .B1(new_n714), .B2(new_n661), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n587), .B1(new_n684), .B2(new_n592), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n501), .A2(new_n550), .A3(new_n507), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n651), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n663), .B1(KEYINPUT26), .B2(new_n709), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n681), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT89), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(KEYINPUT89), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n717), .A2(new_n724), .B1(new_n716), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G330), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n551), .A2(new_n634), .A3(new_n696), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT88), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n659), .A2(new_n587), .A3(new_n681), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n633), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT88), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(new_n733), .A3(new_n551), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n502), .A2(new_n277), .A3(new_n559), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n546), .A2(KEYINPUT87), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n736), .A2(new_n615), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n546), .A2(new_n561), .A3(new_n461), .A4(new_n469), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n611), .B(G179), .C1(new_n613), .C2(new_n614), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(KEYINPUT30), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n744), .B1(new_n740), .B2(new_n741), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n739), .A2(new_n743), .A3(new_n745), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n746), .A2(KEYINPUT31), .A3(new_n690), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n746), .B2(new_n690), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n728), .B1(new_n735), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n727), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n707), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n686), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(new_n728), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT91), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n672), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n207), .B1(new_n757), .B2(G45), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n702), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n689), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n753), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n760), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n211), .A2(G355), .A3(new_n270), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n701), .A2(new_n270), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(G45), .B2(new_n226), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n240), .A2(new_n287), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n767), .B1(G116), .B2(new_n211), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n223), .B1(new_n208), .B2(G169), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT92), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n764), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n766), .B1(new_n771), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n208), .A2(new_n277), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n544), .A2(new_n396), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n544), .A2(G179), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n208), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n785), .B1(G294), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT94), .Z(new_n790));
  NOR2_X1   g0590(.A1(new_n208), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n779), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n396), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n792), .A2(new_n793), .B1(new_n795), .B2(new_n454), .ZN(new_n796));
  XOR2_X1   g0596(.A(KEYINPUT33), .B(G317), .Z(new_n797));
  NAND2_X1  g0597(.A1(new_n778), .A2(new_n794), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n791), .A2(new_n782), .ZN(new_n799));
  INV_X1    g0599(.A(G329), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n797), .A2(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n778), .A2(G190), .A3(new_n396), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n475), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n796), .A2(new_n801), .A3(new_n804), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n787), .A2(new_n534), .B1(new_n798), .B2(new_n203), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT93), .ZN(new_n807));
  INV_X1    g0607(.A(new_n792), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G87), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n202), .B2(new_n802), .ZN(new_n810));
  INV_X1    g0610(.A(G159), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT32), .B1(new_n799), .B2(new_n811), .ZN(new_n812));
  OAI211_X1 g0612(.A(new_n812), .B(new_n270), .C1(new_n329), .C2(new_n795), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n780), .A2(new_n201), .B1(new_n783), .B2(new_n214), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n799), .A2(KEYINPUT32), .A3(new_n811), .ZN(new_n815));
  NOR4_X1   g0615(.A1(new_n810), .A2(new_n813), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n790), .A2(new_n805), .B1(new_n807), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n775), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n777), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT95), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n756), .A2(new_n761), .B1(new_n765), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n818), .A2(new_n763), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n795), .A2(new_n527), .B1(new_n799), .B2(new_n784), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT96), .Z(new_n825));
  OAI22_X1  g0625(.A1(new_n780), .A2(new_n793), .B1(new_n792), .B2(new_n329), .ZN(new_n826));
  INV_X1    g0626(.A(new_n603), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n827), .A2(new_n783), .B1(new_n798), .B2(new_n454), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n475), .B1(new_n802), .B2(new_n829), .C1(new_n534), .C2(new_n787), .ZN(new_n830));
  NOR4_X1   g0630(.A1(new_n825), .A2(new_n826), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G137), .ZN(new_n832));
  INV_X1    g0632(.A(G150), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n780), .A2(new_n832), .B1(new_n798), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT97), .Z(new_n835));
  INV_X1    g0635(.A(new_n802), .ZN(new_n836));
  INV_X1    g0636(.A(new_n783), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n836), .A2(G143), .B1(new_n837), .B2(G159), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT34), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n270), .B1(new_n792), .B2(new_n201), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n795), .A2(new_n203), .B1(new_n799), .B2(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(G58), .C2(new_n788), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n831), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n760), .B1(G77), .B2(new_n823), .C1(new_n845), .C2(new_n818), .ZN(new_n846));
  OR2_X1    g0646(.A1(new_n846), .A2(KEYINPUT98), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(KEYINPUT98), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n339), .A2(new_n690), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n690), .A2(new_n324), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n337), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n850), .B1(new_n339), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n847), .B(new_n848), .C1(new_n763), .C2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n340), .A2(new_n690), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n661), .B2(new_n668), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT99), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n690), .B1(new_n661), .B2(new_n668), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n859), .B2(new_n853), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(new_n339), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(new_n849), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n722), .A2(KEYINPUT99), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n857), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n766), .B1(new_n864), .B2(new_n750), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n855), .B1(new_n720), .B2(new_n721), .ZN(new_n866));
  INV_X1    g0666(.A(new_n863), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT99), .B1(new_n722), .B2(new_n862), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n750), .B(new_n866), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n854), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT100), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT100), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n873), .B(new_n854), .C1(new_n865), .C2(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(G384));
  AOI211_X1 g0675(.A(new_n510), .B(new_n224), .C1(new_n483), .C2(KEYINPUT35), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(KEYINPUT35), .B2(new_n483), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT36), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n214), .A2(new_n201), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n879), .A2(new_n374), .B1(G50), .B2(new_n203), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(G1), .A3(new_n672), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT101), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n361), .B1(new_n379), .B2(new_n381), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n399), .B1(new_n679), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n359), .A2(new_n885), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT37), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n387), .A2(new_n392), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n387), .A2(new_n680), .ZN(new_n890));
  XNOR2_X1  g0690(.A(KEYINPUT102), .B(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n399), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n885), .A2(new_n679), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n394), .B2(new_n403), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n896));
  INV_X1    g0696(.A(new_n891), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n399), .B1(new_n359), .B2(new_n382), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n382), .A2(new_n679), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n892), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n406), .A2(new_n899), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT38), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n884), .B1(new_n896), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n893), .A2(new_n895), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT38), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n441), .A2(new_n447), .A3(new_n681), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n904), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n395), .A2(new_n680), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n907), .A2(new_n908), .ZN(new_n914));
  INV_X1    g0714(.A(new_n435), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n447), .A2(new_n690), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n640), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n447), .B(new_n690), .C1(new_n441), .C2(new_n435), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n866), .B2(new_n849), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n913), .B1(new_n914), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT103), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n912), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g0724(.A(KEYINPUT103), .B(new_n913), .C1(new_n914), .C2(new_n921), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n726), .A2(new_n449), .ZN(new_n927));
  INV_X1    g0727(.A(new_n647), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n926), .B(new_n929), .ZN(new_n930));
  NOR4_X1   g0730(.A1(new_n719), .A2(new_n731), .A3(new_n633), .A4(KEYINPUT88), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n733), .B1(new_n732), .B2(new_n551), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n749), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n862), .B1(new_n917), .B2(new_n918), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n933), .B(new_n934), .C1(new_n896), .C2(new_n903), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT40), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n919), .A2(new_n853), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n735), .B2(new_n749), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n914), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n449), .B1(new_n735), .B2(new_n749), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n728), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n942), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n930), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n207), .B2(new_n757), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n930), .A2(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n883), .B1(new_n946), .B2(new_n947), .ZN(G367));
  INV_X1    g0748(.A(new_n768), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n232), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n776), .B1(new_n211), .B2(new_n316), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n760), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n780), .ZN(new_n953));
  INV_X1    g0753(.A(new_n799), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n953), .A2(G143), .B1(new_n954), .B2(G137), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n201), .B2(new_n783), .C1(new_n833), .C2(new_n802), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n787), .A2(new_n203), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n270), .B1(new_n798), .B2(new_n811), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n792), .A2(new_n202), .B1(new_n795), .B2(new_n214), .ZN(new_n959));
  NOR4_X1   g0759(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n270), .B1(new_n836), .B2(G303), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT110), .B(G317), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n961), .B1(new_n534), .B2(new_n795), .C1(new_n799), .C2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n827), .A2(new_n792), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n964), .A2(KEYINPUT46), .B1(new_n329), .B2(new_n787), .ZN(new_n965));
  NAND2_X1  g0765(.A1(KEYINPUT46), .A2(G116), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n829), .A2(new_n798), .B1(new_n792), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT109), .B(G311), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n780), .A2(new_n968), .B1(new_n783), .B2(new_n454), .ZN(new_n969));
  NOR4_X1   g0769(.A1(new_n963), .A2(new_n965), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n960), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT47), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n818), .B1(new_n971), .B2(KEYINPUT47), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n952), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n681), .A2(new_n549), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n652), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(KEYINPUT104), .C1(new_n708), .C2(new_n975), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(KEYINPUT104), .B2(new_n976), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n764), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n974), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n695), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT44), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n492), .A2(new_n498), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n505), .A3(new_n690), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT105), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n984), .A2(new_n690), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n989), .A2(new_n501), .A3(new_n507), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n987), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  OR3_X1    g0791(.A1(new_n699), .A2(new_n983), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n983), .B1(new_n699), .B2(new_n991), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n992), .A2(KEYINPUT108), .A3(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n699), .A2(new_n991), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT45), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT45), .B1(new_n699), .B2(new_n991), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n998), .A2(new_n999), .B1(KEYINPUT108), .B2(new_n993), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n982), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n998), .A2(new_n999), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n993), .A2(KEYINPUT108), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n1002), .A2(new_n695), .A3(new_n994), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n655), .A2(new_n690), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n697), .B1(new_n694), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n689), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n751), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n751), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n702), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n759), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n991), .A2(new_n698), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT42), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n991), .A2(new_n592), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n690), .B1(new_n1016), .B2(new_n507), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n689), .A2(new_n694), .A3(new_n991), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT106), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n979), .A2(KEYINPUT43), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1021), .A2(KEYINPUT106), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1024), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1020), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1021), .B(KEYINPUT106), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n1023), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1031), .A2(new_n1019), .A3(new_n1018), .A4(new_n1026), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n981), .B1(new_n1013), .B2(new_n1033), .ZN(G387));
  INV_X1    g0834(.A(G77), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n287), .B1(new_n203), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n704), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(KEYINPUT111), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n252), .A2(KEYINPUT50), .A3(new_n201), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT50), .B1(new_n252), .B2(new_n201), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1038), .B1(KEYINPUT111), .B2(new_n1037), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1041), .B(new_n768), .C1(new_n236), .C2(new_n287), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1037), .A2(new_n211), .A3(new_n270), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(G107), .C2(new_n211), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n766), .B1(new_n1044), .B2(new_n776), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n475), .B1(new_n799), .B2(new_n781), .C1(new_n827), .C2(new_n795), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n802), .A2(new_n962), .B1(new_n783), .B2(new_n793), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n780), .A2(new_n803), .B1(new_n798), .B2(new_n968), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT113), .Z(new_n1050));
  AND2_X1   g0850(.A1(new_n1050), .A2(KEYINPUT48), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1050), .A2(KEYINPUT48), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n787), .A2(new_n454), .B1(new_n792), .B2(new_n829), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT112), .ZN(new_n1054));
  NOR3_X1   g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1046), .B1(new_n1055), .B2(KEYINPUT49), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(KEYINPUT49), .B2(new_n1055), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n792), .A2(new_n214), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n270), .B1(new_n795), .B2(new_n534), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(G68), .C2(new_n837), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n953), .A2(G159), .B1(new_n954), .B2(G150), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n798), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n836), .A2(G50), .B1(new_n1062), .B2(new_n252), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n788), .A2(new_n539), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1045), .B1(new_n694), .B2(new_n980), .C1(new_n1066), .C2(new_n818), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT114), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n759), .B2(new_n1008), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n751), .A2(new_n1008), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1009), .A2(new_n702), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(G393));
  NAND3_X1  g0872(.A1(new_n1001), .A2(new_n759), .A3(new_n1004), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n776), .B1(new_n534), .B2(new_n211), .C1(new_n949), .C2(new_n243), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n766), .B1(new_n1074), .B2(KEYINPUT115), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(KEYINPUT115), .B2(new_n1074), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n836), .A2(G311), .B1(new_n953), .B2(G317), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n454), .A2(new_n792), .B1(new_n783), .B2(new_n829), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n798), .A2(new_n793), .B1(new_n799), .B2(new_n803), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n475), .B1(new_n795), .B2(new_n329), .C1(new_n787), .C2(new_n827), .ZN(new_n1081));
  OR4_X1    g0881(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n787), .A2(new_n1035), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n795), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n475), .B(new_n1083), .C1(G87), .C2(new_n1084), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n802), .A2(new_n811), .B1(new_n780), .B2(new_n833), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT51), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n252), .A2(new_n837), .B1(new_n808), .B2(G68), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(G50), .A2(new_n1062), .B1(new_n954), .B2(G143), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1082), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1076), .B1(new_n775), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n991), .B2(new_n980), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n702), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1073), .B(new_n1093), .C1(new_n1094), .C2(new_n1095), .ZN(G390));
  NAND3_X1  g0896(.A1(new_n933), .A2(G330), .A3(new_n934), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT117), .A4(G330), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n933), .A2(G330), .A3(new_n853), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1099), .A2(new_n1100), .B1(new_n920), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n857), .A2(new_n850), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT118), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1101), .A2(new_n1104), .A3(new_n920), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n850), .B1(new_n715), .B2(new_n861), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1097), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1101), .B2(new_n920), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1102), .A2(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n450), .A2(new_n750), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1110), .B(new_n647), .C1(new_n726), .C2(new_n449), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n919), .B1(new_n857), .B2(new_n850), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n904), .A2(new_n909), .B1(new_n1114), .B2(new_n910), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n910), .B(KEYINPUT116), .Z(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n896), .B2(new_n903), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n713), .A2(new_n711), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n712), .B1(new_n667), .B2(new_n665), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n681), .B(new_n861), .C1(new_n1120), .C2(new_n720), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n920), .B1(new_n1121), .B2(new_n849), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1099), .B(new_n1100), .C1(new_n1115), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1114), .A2(new_n910), .ZN(new_n1125));
  AND3_X1   g0925(.A1(new_n907), .A2(KEYINPUT39), .A3(new_n908), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n901), .A2(new_n902), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n906), .ZN(new_n1128));
  AOI21_X1  g0928(.A(KEYINPUT39), .B1(new_n1128), .B2(new_n908), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1125), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  OR2_X1    g0930(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1097), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1124), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n703), .B1(new_n1113), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1133), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1101), .A2(new_n920), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT117), .B1(new_n750), .B2(new_n934), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1100), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1103), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1136), .A2(KEYINPUT118), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(new_n1097), .A3(new_n1106), .A4(new_n1105), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1111), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1135), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1134), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n762), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n760), .B1(new_n823), .B2(new_n252), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n792), .A2(new_n833), .ZN(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G137), .A2(new_n1062), .B1(new_n954), .B2(G125), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n201), .C2(new_n795), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT54), .B(G143), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G128), .A2(new_n953), .B1(new_n837), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n475), .B1(new_n836), .B2(G132), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1156), .B(new_n1157), .C1(new_n811), .C2(new_n787), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n836), .A2(G116), .B1(new_n954), .B2(G294), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n534), .B2(new_n783), .C1(new_n329), .C2(new_n798), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G283), .A2(new_n953), .B1(new_n1084), .B2(G68), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1083), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1161), .A2(new_n1162), .A3(new_n475), .A4(new_n809), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1153), .A2(new_n1158), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1148), .B1(new_n1164), .B2(new_n775), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1147), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n1133), .B2(new_n758), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1146), .A2(new_n1168), .ZN(G378));
  AND2_X1   g0969(.A1(new_n914), .A2(new_n921), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT103), .B1(new_n1170), .B2(new_n913), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n922), .A2(new_n923), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n912), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n679), .B1(new_n262), .B2(new_n268), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n646), .B2(new_n295), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n636), .B(new_n1176), .C1(new_n645), .C2(new_n308), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1175), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n310), .A2(new_n1176), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n646), .A2(new_n295), .A3(new_n1177), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n1174), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n941), .B2(G330), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n728), .B(new_n1184), .C1(new_n936), .C2(new_n940), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1173), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n941), .A2(G330), .A3(new_n1185), .ZN(new_n1189));
  AOI21_X1  g0989(.A(KEYINPUT40), .B1(new_n907), .B2(new_n908), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(KEYINPUT40), .A2(new_n935), .B1(new_n1190), .B2(new_n938), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1184), .B1(new_n1191), .B2(new_n728), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n926), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1188), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1103), .B1(new_n1196), .B2(new_n1136), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1195), .A2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1112), .B1(new_n1198), .B2(new_n1133), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1194), .A2(new_n1199), .A3(KEYINPUT57), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n702), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1194), .B2(new_n1199), .ZN(new_n1202));
  OR2_X1    g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n760), .B1(new_n823), .B2(G50), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n953), .A2(G125), .ZN(new_n1205));
  INV_X1    g1005(.A(G128), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n802), .C1(new_n792), .C2(new_n1154), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n842), .A2(new_n798), .B1(new_n783), .B2(new_n832), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT120), .Z(new_n1209));
  AOI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(G150), .C2(new_n788), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(KEYINPUT59), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n253), .A2(new_n286), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT121), .B(G124), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n954), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n811), .B2(new_n795), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n783), .A2(new_n316), .B1(new_n799), .B2(new_n454), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n475), .A2(new_n286), .ZN(new_n1220));
  NOR4_X1   g1020(.A1(new_n1219), .A2(new_n957), .A3(new_n1058), .A4(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n795), .A2(new_n202), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G107), .B2(new_n836), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G116), .A2(new_n953), .B1(new_n1062), .B2(G97), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1221), .A2(new_n1223), .A3(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT58), .ZN(new_n1226));
  OR2_X1    g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1220), .A2(new_n201), .A3(new_n1214), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n775), .B1(new_n1218), .B2(new_n1230), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT122), .Z(new_n1232));
  AOI211_X1 g1032(.A(new_n1204), .B(new_n1232), .C1(new_n762), .C2(new_n1184), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1194), .B2(new_n759), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1203), .A2(new_n1234), .ZN(G375));
  OAI21_X1  g1035(.A(new_n759), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n760), .B1(new_n823), .B2(G68), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n780), .A2(new_n842), .B1(new_n799), .B2(new_n1206), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(new_n475), .A3(new_n1222), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(G150), .A2(new_n837), .B1(new_n1062), .B2(new_n1155), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n836), .A2(G137), .B1(new_n808), .B2(G159), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n788), .A2(G50), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1239), .A2(new_n1240), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1064), .B1(new_n329), .B2(new_n783), .C1(new_n827), .C2(new_n798), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n802), .A2(new_n454), .B1(new_n780), .B2(new_n829), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n792), .A2(new_n534), .B1(new_n799), .B2(new_n793), .ZN(new_n1246));
  OR3_X1    g1046(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n475), .B1(new_n795), .B2(new_n1035), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT124), .Z(new_n1249));
  OAI21_X1  g1049(.A(new_n1243), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1237), .B1(new_n1250), .B2(new_n775), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n919), .B2(new_n763), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1236), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1141), .A2(new_n1143), .A3(new_n1111), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(new_n1012), .B(KEYINPUT123), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1113), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(G381));
  OR3_X1    g1058(.A1(G390), .A2(G396), .A3(G393), .ZN(new_n1259));
  NOR4_X1   g1059(.A1(new_n1259), .A2(G384), .A3(G387), .A4(G381), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1167), .B1(new_n1134), .B2(new_n1145), .ZN(new_n1261));
  INV_X1    g1061(.A(G375), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .ZN(G407));
  INV_X1    g1063(.A(G213), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1264), .A2(G343), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1262), .A2(new_n1261), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(G407), .A2(G213), .A3(new_n1266), .ZN(G409));
  NAND2_X1  g1067(.A1(new_n1265), .A2(G2897), .ZN(new_n1268));
  INV_X1    g1068(.A(G384), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1141), .A2(new_n1111), .A3(new_n1143), .A4(KEYINPUT60), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1270), .A2(new_n702), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT60), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1255), .B1(new_n1144), .B2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1269), .B1(new_n1274), .B2(new_n1254), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1253), .B(G384), .C1(new_n1271), .C2(new_n1273), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1268), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1272), .B1(new_n1109), .B2(new_n1112), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1270), .A2(new_n702), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1254), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(G384), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1274), .A2(new_n1269), .A3(new_n1254), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1268), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1234), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1194), .A2(new_n1199), .A3(new_n1256), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1234), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1261), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1265), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1277), .A2(new_n1286), .A3(KEYINPUT125), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1289), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1299), .B1(new_n1296), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(G390), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1302), .ZN(new_n1303));
  XNOR2_X1  g1103(.A(G393), .B(new_n821), .ZN(new_n1304));
  OAI211_X1 g1104(.A(G390), .B(new_n981), .C1(new_n1013), .C2(new_n1033), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1304), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1306), .A2(new_n1307), .A3(KEYINPUT61), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1265), .B1(new_n1290), .B2(new_n1293), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1300), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1309), .A2(KEYINPUT63), .A3(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1298), .A2(new_n1301), .A3(new_n1308), .A4(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT62), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1309), .A2(new_n1313), .A3(new_n1310), .ZN(new_n1314));
  XOR2_X1   g1114(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1309), .B2(new_n1287), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1313), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1314), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1312), .B1(new_n1318), .B2(new_n1319), .ZN(G405));
  NAND2_X1  g1120(.A1(G375), .A2(new_n1261), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1290), .A3(new_n1310), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G378), .B1(new_n1203), .B2(new_n1234), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1290), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1300), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1322), .A2(new_n1319), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1319), .B1(new_n1322), .B2(new_n1325), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(G402));
endmodule


