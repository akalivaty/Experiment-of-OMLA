

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n608), .A2(n607), .ZN(n611) );
  XNOR2_X1 U553 ( .A(KEYINPUT96), .B(KEYINPUT30), .ZN(n653) );
  XNOR2_X1 U554 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U555 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n659) );
  XNOR2_X1 U556 ( .A(n660), .B(n659), .ZN(n661) );
  AND2_X1 U557 ( .A1(n663), .A2(n669), .ZN(n664) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n533) );
  AND2_X1 U559 ( .A1(n540), .A2(G2104), .ZN(n873) );
  NAND2_X1 U560 ( .A1(n874), .A2(G138), .ZN(n536) );
  NOR2_X1 U561 ( .A1(n588), .A2(G651), .ZN(n786) );
  OR2_X1 U562 ( .A1(n538), .A2(n539), .ZN(n544) );
  AND2_X1 U563 ( .A1(n546), .A2(n545), .ZN(G164) );
  INV_X1 U564 ( .A(G651), .ZN(n525) );
  NOR2_X1 U565 ( .A1(G543), .A2(n525), .ZN(n520) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n520), .Z(n785) );
  NAND2_X1 U567 ( .A1(G63), .A2(n785), .ZN(n522) );
  XOR2_X1 U568 ( .A(KEYINPUT0), .B(G543), .Z(n588) );
  NAND2_X1 U569 ( .A1(G51), .A2(n786), .ZN(n521) );
  NAND2_X1 U570 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U571 ( .A(KEYINPUT6), .B(n523), .ZN(n530) );
  NOR2_X1 U572 ( .A1(G543), .A2(G651), .ZN(n781) );
  NAND2_X1 U573 ( .A1(n781), .A2(G89), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n524), .B(KEYINPUT4), .ZN(n527) );
  NOR2_X1 U575 ( .A1(n588), .A2(n525), .ZN(n779) );
  NAND2_X1 U576 ( .A1(G76), .A2(n779), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U578 ( .A(n528), .B(KEYINPUT5), .Z(n529) );
  NOR2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT74), .B(n531), .Z(n532) );
  XNOR2_X1 U581 ( .A(KEYINPUT7), .B(n532), .ZN(G168) );
  INV_X1 U582 ( .A(KEYINPUT85), .ZN(n538) );
  INV_X1 U583 ( .A(G2105), .ZN(n540) );
  NAND2_X1 U584 ( .A1(G102), .A2(n873), .ZN(n537) );
  XNOR2_X1 U585 ( .A(KEYINPUT64), .B(n533), .ZN(n535) );
  INV_X1 U586 ( .A(KEYINPUT17), .ZN(n534) );
  XNOR2_X2 U587 ( .A(n535), .B(n534), .ZN(n874) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n539) );
  NAND2_X1 U589 ( .A1(n538), .A2(n539), .ZN(n546) );
  AND2_X1 U590 ( .A1(G2104), .A2(G2105), .ZN(n880) );
  NAND2_X1 U591 ( .A1(G114), .A2(n880), .ZN(n542) );
  NOR2_X1 U592 ( .A1(G2104), .A2(n540), .ZN(n878) );
  NAND2_X1 U593 ( .A1(G126), .A2(n878), .ZN(n541) );
  AND2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n543) );
  AND2_X1 U595 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U596 ( .A1(G137), .A2(n874), .ZN(n549) );
  NAND2_X1 U597 ( .A1(G101), .A2(n873), .ZN(n547) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n547), .Z(n548) );
  NAND2_X1 U599 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U600 ( .A1(G113), .A2(n880), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G125), .A2(n878), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X2 U603 ( .A1(n553), .A2(n552), .ZN(G160) );
  NAND2_X1 U604 ( .A1(G86), .A2(n781), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G61), .A2(n785), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n558) );
  NAND2_X1 U607 ( .A1(n779), .A2(G73), .ZN(n556) );
  XOR2_X1 U608 ( .A(KEYINPUT2), .B(n556), .Z(n557) );
  NOR2_X1 U609 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U610 ( .A1(n786), .A2(G48), .ZN(n559) );
  NAND2_X1 U611 ( .A1(n560), .A2(n559), .ZN(G305) );
  XNOR2_X1 U612 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n564) );
  NAND2_X1 U613 ( .A1(G90), .A2(n781), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G77), .A2(n779), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U616 ( .A(n564), .B(n563), .ZN(n570) );
  NAND2_X1 U617 ( .A1(G52), .A2(n786), .ZN(n565) );
  XNOR2_X1 U618 ( .A(n565), .B(KEYINPUT66), .ZN(n568) );
  NAND2_X1 U619 ( .A1(n785), .A2(G64), .ZN(n566) );
  XOR2_X1 U620 ( .A(KEYINPUT65), .B(n566), .Z(n567) );
  NAND2_X1 U621 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X1 U622 ( .A1(n570), .A2(n569), .ZN(G171) );
  NAND2_X1 U623 ( .A1(G91), .A2(n781), .ZN(n572) );
  NAND2_X1 U624 ( .A1(G78), .A2(n779), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U626 ( .A1(n785), .A2(G65), .ZN(n573) );
  XOR2_X1 U627 ( .A(KEYINPUT68), .B(n573), .Z(n574) );
  NOR2_X1 U628 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U629 ( .A1(n786), .A2(G53), .ZN(n576) );
  NAND2_X1 U630 ( .A1(n577), .A2(n576), .ZN(G299) );
  XNOR2_X1 U631 ( .A(KEYINPUT75), .B(KEYINPUT8), .ZN(n578) );
  XNOR2_X1 U632 ( .A(n578), .B(G168), .ZN(G286) );
  NAND2_X1 U633 ( .A1(G88), .A2(n781), .ZN(n580) );
  NAND2_X1 U634 ( .A1(G75), .A2(n779), .ZN(n579) );
  NAND2_X1 U635 ( .A1(n580), .A2(n579), .ZN(n584) );
  NAND2_X1 U636 ( .A1(G62), .A2(n785), .ZN(n582) );
  NAND2_X1 U637 ( .A1(G50), .A2(n786), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U639 ( .A1(n584), .A2(n583), .ZN(G166) );
  INV_X1 U640 ( .A(G166), .ZN(G303) );
  NAND2_X1 U641 ( .A1(G49), .A2(n786), .ZN(n586) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n585) );
  NAND2_X1 U643 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U644 ( .A1(n785), .A2(n587), .ZN(n590) );
  NAND2_X1 U645 ( .A1(n588), .A2(G87), .ZN(n589) );
  NAND2_X1 U646 ( .A1(n590), .A2(n589), .ZN(G288) );
  NAND2_X1 U647 ( .A1(G85), .A2(n781), .ZN(n592) );
  NAND2_X1 U648 ( .A1(G72), .A2(n779), .ZN(n591) );
  NAND2_X1 U649 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U650 ( .A1(G60), .A2(n785), .ZN(n594) );
  NAND2_X1 U651 ( .A1(G47), .A2(n786), .ZN(n593) );
  NAND2_X1 U652 ( .A1(n594), .A2(n593), .ZN(n595) );
  OR2_X1 U653 ( .A1(n596), .A2(n595), .ZN(G290) );
  NOR2_X1 U654 ( .A1(G164), .A2(G1384), .ZN(n701) );
  NAND2_X1 U655 ( .A1(G40), .A2(G160), .ZN(n597) );
  XNOR2_X1 U656 ( .A(n597), .B(KEYINPUT86), .ZN(n702) );
  INV_X1 U657 ( .A(n702), .ZN(n598) );
  NAND2_X1 U658 ( .A1(n701), .A2(n598), .ZN(n649) );
  NAND2_X1 U659 ( .A1(G8), .A2(n649), .ZN(n698) );
  NOR2_X1 U660 ( .A1(G1981), .A2(G305), .ZN(n599) );
  XOR2_X1 U661 ( .A(n599), .B(KEYINPUT24), .Z(n600) );
  NOR2_X1 U662 ( .A1(n698), .A2(n600), .ZN(n692) );
  XNOR2_X1 U663 ( .A(G1981), .B(G305), .ZN(n957) );
  NOR2_X1 U664 ( .A1(G1966), .A2(n698), .ZN(n651) );
  INV_X1 U665 ( .A(n651), .ZN(n663) );
  XNOR2_X1 U666 ( .A(G2078), .B(KEYINPUT92), .ZN(n601) );
  XNOR2_X1 U667 ( .A(n601), .B(KEYINPUT25), .ZN(n995) );
  INV_X1 U668 ( .A(n649), .ZN(n634) );
  NOR2_X1 U669 ( .A1(n995), .A2(n649), .ZN(n603) );
  AND2_X1 U670 ( .A1(n649), .A2(G1961), .ZN(n602) );
  NOR2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n656) );
  NAND2_X1 U672 ( .A1(G171), .A2(n656), .ZN(n648) );
  INV_X1 U673 ( .A(G299), .ZN(n794) );
  XOR2_X1 U674 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n605) );
  NAND2_X1 U675 ( .A1(G2072), .A2(n634), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n605), .B(n604), .ZN(n608) );
  NAND2_X1 U677 ( .A1(G1956), .A2(n649), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT94), .B(n606), .Z(n607) );
  NOR2_X1 U679 ( .A1(n794), .A2(n611), .ZN(n610) );
  XNOR2_X1 U680 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n609) );
  XNOR2_X1 U681 ( .A(n610), .B(n609), .ZN(n645) );
  NAND2_X1 U682 ( .A1(n794), .A2(n611), .ZN(n643) );
  NAND2_X1 U683 ( .A1(n781), .A2(G81), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(KEYINPUT12), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G68), .A2(n779), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U687 ( .A(KEYINPUT13), .B(n615), .Z(n619) );
  NAND2_X1 U688 ( .A1(G56), .A2(n785), .ZN(n616) );
  XNOR2_X1 U689 ( .A(n616), .B(KEYINPUT14), .ZN(n617) );
  XNOR2_X1 U690 ( .A(n617), .B(KEYINPUT71), .ZN(n618) );
  NOR2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n786), .A2(G43), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n950) );
  INV_X1 U694 ( .A(G1996), .ZN(n994) );
  NOR2_X1 U695 ( .A1(n649), .A2(n994), .ZN(n622) );
  XOR2_X1 U696 ( .A(n622), .B(KEYINPUT26), .Z(n624) );
  NAND2_X1 U697 ( .A1(n649), .A2(G1341), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U699 ( .A1(n950), .A2(n625), .ZN(n638) );
  NAND2_X1 U700 ( .A1(n785), .A2(G66), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G92), .A2(n781), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G79), .A2(n779), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U704 ( .A1(G54), .A2(n786), .ZN(n628) );
  XNOR2_X1 U705 ( .A(KEYINPUT73), .B(n628), .ZN(n629) );
  NOR2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U708 ( .A(KEYINPUT15), .B(n633), .Z(n951) );
  NAND2_X1 U709 ( .A1(G1348), .A2(n649), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G2067), .A2(n634), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n639) );
  NOR2_X1 U712 ( .A1(n951), .A2(n639), .ZN(n637) );
  OR2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n951), .A2(n639), .ZN(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U718 ( .A(KEYINPUT29), .B(n646), .Z(n647) );
  NAND2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n662) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n649), .ZN(n665) );
  INV_X1 U721 ( .A(n665), .ZN(n650) );
  NAND2_X1 U722 ( .A1(G8), .A2(n650), .ZN(n652) );
  OR2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n655), .A2(G168), .ZN(n658) );
  NOR2_X1 U725 ( .A1(G171), .A2(n656), .ZN(n657) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n669) );
  XNOR2_X1 U728 ( .A(KEYINPUT98), .B(n664), .ZN(n668) );
  NAND2_X1 U729 ( .A1(G8), .A2(n665), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT91), .B(n666), .Z(n667) );
  NAND2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n678) );
  NAND2_X1 U732 ( .A1(n669), .A2(G286), .ZN(n674) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n698), .ZN(n671) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n649), .ZN(n670) );
  NOR2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U736 ( .A1(n672), .A2(G303), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U738 ( .A1(n675), .A2(G8), .ZN(n676) );
  XNOR2_X1 U739 ( .A(n676), .B(KEYINPUT32), .ZN(n677) );
  NAND2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n693) );
  INV_X1 U741 ( .A(n693), .ZN(n680) );
  OR2_X1 U742 ( .A1(G1976), .A2(G288), .ZN(n684) );
  INV_X1 U743 ( .A(G1971), .ZN(n979) );
  NAND2_X1 U744 ( .A1(G166), .A2(n979), .ZN(n679) );
  NAND2_X1 U745 ( .A1(n684), .A2(n679), .ZN(n943) );
  NOR2_X1 U746 ( .A1(n680), .A2(n943), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n698), .A2(n681), .ZN(n682) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n944) );
  NAND2_X1 U749 ( .A1(n682), .A2(n944), .ZN(n683) );
  INV_X1 U750 ( .A(KEYINPUT33), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n683), .A2(n686), .ZN(n689) );
  OR2_X1 U752 ( .A1(n698), .A2(n684), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n687), .B(KEYINPUT99), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U756 ( .A1(n957), .A2(n690), .ZN(n691) );
  NOR2_X1 U757 ( .A1(n692), .A2(n691), .ZN(n700) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n694) );
  NAND2_X1 U759 ( .A1(G8), .A2(n694), .ZN(n695) );
  NAND2_X1 U760 ( .A1(n693), .A2(n695), .ZN(n696) );
  XNOR2_X1 U761 ( .A(KEYINPUT100), .B(n696), .ZN(n697) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n733) );
  NOR2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n746) );
  NAND2_X1 U765 ( .A1(G104), .A2(n873), .ZN(n704) );
  NAND2_X1 U766 ( .A1(G140), .A2(n874), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n706) );
  XOR2_X1 U768 ( .A(KEYINPUT34), .B(KEYINPUT87), .Z(n705) );
  XNOR2_X1 U769 ( .A(n706), .B(n705), .ZN(n711) );
  NAND2_X1 U770 ( .A1(G116), .A2(n880), .ZN(n708) );
  NAND2_X1 U771 ( .A1(G128), .A2(n878), .ZN(n707) );
  NAND2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U773 ( .A(KEYINPUT35), .B(n709), .Z(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U775 ( .A(n712), .B(KEYINPUT36), .ZN(n713) );
  XNOR2_X1 U776 ( .A(n713), .B(KEYINPUT88), .ZN(n893) );
  XNOR2_X1 U777 ( .A(KEYINPUT37), .B(G2067), .ZN(n744) );
  NOR2_X1 U778 ( .A1(n893), .A2(n744), .ZN(n915) );
  NAND2_X1 U779 ( .A1(n746), .A2(n915), .ZN(n742) );
  NAND2_X1 U780 ( .A1(n880), .A2(G107), .ZN(n714) );
  XOR2_X1 U781 ( .A(KEYINPUT89), .B(n714), .Z(n716) );
  NAND2_X1 U782 ( .A1(n878), .A2(G119), .ZN(n715) );
  NAND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U784 ( .A(KEYINPUT90), .B(n717), .Z(n721) );
  NAND2_X1 U785 ( .A1(n874), .A2(G131), .ZN(n719) );
  NAND2_X1 U786 ( .A1(G95), .A2(n873), .ZN(n718) );
  AND2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n859) );
  AND2_X1 U789 ( .A1(n859), .A2(G1991), .ZN(n730) );
  NAND2_X1 U790 ( .A1(n878), .A2(G129), .ZN(n723) );
  NAND2_X1 U791 ( .A1(G141), .A2(n874), .ZN(n722) );
  NAND2_X1 U792 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U793 ( .A1(n873), .A2(G105), .ZN(n724) );
  XOR2_X1 U794 ( .A(KEYINPUT38), .B(n724), .Z(n725) );
  NOR2_X1 U795 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n880), .A2(G117), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n888) );
  AND2_X1 U798 ( .A1(n888), .A2(G1996), .ZN(n729) );
  NOR2_X1 U799 ( .A1(n730), .A2(n729), .ZN(n920) );
  INV_X1 U800 ( .A(n920), .ZN(n731) );
  NAND2_X1 U801 ( .A1(n731), .A2(n746), .ZN(n736) );
  AND2_X1 U802 ( .A1(n742), .A2(n736), .ZN(n732) );
  AND2_X1 U803 ( .A1(n733), .A2(n732), .ZN(n735) );
  XNOR2_X1 U804 ( .A(G1986), .B(G290), .ZN(n941) );
  NAND2_X1 U805 ( .A1(n941), .A2(n746), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n749) );
  NOR2_X1 U807 ( .A1(G1996), .A2(n888), .ZN(n926) );
  INV_X1 U808 ( .A(n736), .ZN(n739) );
  NOR2_X1 U809 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U810 ( .A1(G1991), .A2(n859), .ZN(n922) );
  NOR2_X1 U811 ( .A1(n737), .A2(n922), .ZN(n738) );
  NOR2_X1 U812 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U813 ( .A1(n926), .A2(n740), .ZN(n741) );
  XNOR2_X1 U814 ( .A(KEYINPUT39), .B(n741), .ZN(n743) );
  NAND2_X1 U815 ( .A1(n743), .A2(n742), .ZN(n745) );
  NAND2_X1 U816 ( .A1(n893), .A2(n744), .ZN(n914) );
  NAND2_X1 U817 ( .A1(n745), .A2(n914), .ZN(n747) );
  NAND2_X1 U818 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U819 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U820 ( .A(n750), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U821 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U822 ( .A(G57), .ZN(G237) );
  XOR2_X1 U823 ( .A(KEYINPUT10), .B(KEYINPUT69), .Z(n752) );
  NAND2_X1 U824 ( .A1(G7), .A2(G661), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n752), .B(n751), .ZN(G223) );
  XOR2_X1 U826 ( .A(G223), .B(KEYINPUT70), .Z(n816) );
  NAND2_X1 U827 ( .A1(n816), .A2(G567), .ZN(n753) );
  XOR2_X1 U828 ( .A(KEYINPUT11), .B(n753), .Z(G234) );
  INV_X1 U829 ( .A(G860), .ZN(n761) );
  OR2_X1 U830 ( .A1(n950), .A2(n761), .ZN(G153) );
  INV_X1 U831 ( .A(G171), .ZN(G301) );
  NAND2_X1 U832 ( .A1(G868), .A2(G301), .ZN(n754) );
  XNOR2_X1 U833 ( .A(n754), .B(KEYINPUT72), .ZN(n756) );
  INV_X1 U834 ( .A(n951), .ZN(n777) );
  OR2_X1 U835 ( .A1(G868), .A2(n777), .ZN(n755) );
  NAND2_X1 U836 ( .A1(n756), .A2(n755), .ZN(G284) );
  XOR2_X1 U837 ( .A(G868), .B(KEYINPUT76), .Z(n757) );
  NOR2_X1 U838 ( .A1(G286), .A2(n757), .ZN(n759) );
  NOR2_X1 U839 ( .A1(G868), .A2(G299), .ZN(n758) );
  NOR2_X1 U840 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U841 ( .A(KEYINPUT77), .B(n760), .Z(G297) );
  NAND2_X1 U842 ( .A1(n761), .A2(G559), .ZN(n762) );
  NAND2_X1 U843 ( .A1(n762), .A2(n777), .ZN(n763) );
  XNOR2_X1 U844 ( .A(n763), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U845 ( .A1(G868), .A2(n950), .ZN(n766) );
  NAND2_X1 U846 ( .A1(G868), .A2(n777), .ZN(n764) );
  NOR2_X1 U847 ( .A1(G559), .A2(n764), .ZN(n765) );
  NOR2_X1 U848 ( .A1(n766), .A2(n765), .ZN(G282) );
  NAND2_X1 U849 ( .A1(n878), .A2(G123), .ZN(n767) );
  XNOR2_X1 U850 ( .A(n767), .B(KEYINPUT18), .ZN(n769) );
  NAND2_X1 U851 ( .A1(G135), .A2(n874), .ZN(n768) );
  NAND2_X1 U852 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U853 ( .A(KEYINPUT78), .B(n770), .ZN(n774) );
  NAND2_X1 U854 ( .A1(G99), .A2(n873), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G111), .A2(n880), .ZN(n771) );
  NAND2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U857 ( .A1(n774), .A2(n773), .ZN(n918) );
  XNOR2_X1 U858 ( .A(n918), .B(G2096), .ZN(n776) );
  INV_X1 U859 ( .A(G2100), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(G156) );
  NAND2_X1 U861 ( .A1(G559), .A2(n777), .ZN(n778) );
  XNOR2_X1 U862 ( .A(n778), .B(n950), .ZN(n797) );
  NOR2_X1 U863 ( .A1(n797), .A2(G860), .ZN(n791) );
  NAND2_X1 U864 ( .A1(n779), .A2(G80), .ZN(n780) );
  XOR2_X1 U865 ( .A(KEYINPUT79), .B(n780), .Z(n783) );
  NAND2_X1 U866 ( .A1(n781), .A2(G93), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U868 ( .A(KEYINPUT80), .B(n784), .ZN(n790) );
  NAND2_X1 U869 ( .A1(G67), .A2(n785), .ZN(n788) );
  NAND2_X1 U870 ( .A1(G55), .A2(n786), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U872 ( .A1(n790), .A2(n789), .ZN(n822) );
  XNOR2_X1 U873 ( .A(n791), .B(n822), .ZN(G145) );
  XNOR2_X1 U874 ( .A(KEYINPUT19), .B(G305), .ZN(n792) );
  XNOR2_X1 U875 ( .A(n792), .B(G288), .ZN(n793) );
  XNOR2_X1 U876 ( .A(G166), .B(n793), .ZN(n796) );
  XNOR2_X1 U877 ( .A(G290), .B(n794), .ZN(n795) );
  XNOR2_X1 U878 ( .A(n796), .B(n795), .ZN(n823) );
  XNOR2_X1 U879 ( .A(n823), .B(n797), .ZN(n798) );
  NAND2_X1 U880 ( .A1(n798), .A2(G868), .ZN(n799) );
  XNOR2_X1 U881 ( .A(KEYINPUT81), .B(n799), .ZN(n800) );
  XNOR2_X1 U882 ( .A(n822), .B(n800), .ZN(G295) );
  NAND2_X1 U883 ( .A1(G2078), .A2(G2084), .ZN(n801) );
  XOR2_X1 U884 ( .A(KEYINPUT20), .B(n801), .Z(n802) );
  NAND2_X1 U885 ( .A1(G2090), .A2(n802), .ZN(n803) );
  XNOR2_X1 U886 ( .A(KEYINPUT21), .B(n803), .ZN(n804) );
  NAND2_X1 U887 ( .A1(n804), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U888 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U889 ( .A1(G483), .A2(G661), .ZN(n814) );
  XOR2_X1 U890 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n806) );
  NAND2_X1 U891 ( .A1(G132), .A2(G82), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n806), .B(n805), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n807), .A2(G96), .ZN(n808) );
  NOR2_X1 U894 ( .A1(n808), .A2(G218), .ZN(n809) );
  XNOR2_X1 U895 ( .A(n809), .B(KEYINPUT83), .ZN(n820) );
  NAND2_X1 U896 ( .A1(n820), .A2(G2106), .ZN(n813) );
  NAND2_X1 U897 ( .A1(G120), .A2(G108), .ZN(n810) );
  NOR2_X1 U898 ( .A1(G237), .A2(n810), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G69), .A2(n811), .ZN(n821) );
  NAND2_X1 U900 ( .A1(n821), .A2(G567), .ZN(n812) );
  NAND2_X1 U901 ( .A1(n813), .A2(n812), .ZN(n913) );
  NOR2_X1 U902 ( .A1(n814), .A2(n913), .ZN(n815) );
  XNOR2_X1 U903 ( .A(n815), .B(KEYINPUT84), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G36), .A2(n819), .ZN(G176) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U906 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U907 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U908 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(G188) );
  XNOR2_X1 U910 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U912 ( .A(G132), .ZN(G219) );
  INV_X1 U913 ( .A(G120), .ZN(G236) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  INV_X1 U915 ( .A(G82), .ZN(G220) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  XOR2_X1 U918 ( .A(n822), .B(KEYINPUT112), .Z(n825) );
  XNOR2_X1 U919 ( .A(G171), .B(n823), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n826), .B(n950), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n827), .B(n951), .ZN(n828) );
  XOR2_X1 U923 ( .A(G286), .B(n828), .Z(n829) );
  NOR2_X1 U924 ( .A1(G37), .A2(n829), .ZN(n830) );
  XOR2_X1 U925 ( .A(KEYINPUT113), .B(n830), .Z(G397) );
  XOR2_X1 U926 ( .A(G2474), .B(G1961), .Z(n832) );
  XNOR2_X1 U927 ( .A(G1996), .B(G1991), .ZN(n831) );
  XNOR2_X1 U928 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U929 ( .A(n833), .B(KEYINPUT103), .Z(n835) );
  XNOR2_X1 U930 ( .A(G1971), .B(G1976), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U932 ( .A(G1981), .B(G1956), .Z(n837) );
  XNOR2_X1 U933 ( .A(G1986), .B(G1966), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U935 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U936 ( .A(KEYINPUT104), .B(KEYINPUT41), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n843) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2090), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(G227) );
  NAND2_X1 U947 ( .A1(G124), .A2(n878), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n850), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U949 ( .A1(n880), .A2(G112), .ZN(n852) );
  NAND2_X1 U950 ( .A1(G136), .A2(n874), .ZN(n851) );
  NAND2_X1 U951 ( .A1(n852), .A2(n851), .ZN(n855) );
  NAND2_X1 U952 ( .A1(G100), .A2(n873), .ZN(n853) );
  XNOR2_X1 U953 ( .A(KEYINPUT105), .B(n853), .ZN(n854) );
  NOR2_X1 U954 ( .A1(n855), .A2(n854), .ZN(n856) );
  NAND2_X1 U955 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(KEYINPUT106), .B(n858), .Z(G162) );
  XOR2_X1 U957 ( .A(G160), .B(n859), .Z(n868) );
  NAND2_X1 U958 ( .A1(G103), .A2(n873), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G139), .A2(n874), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n878), .A2(G127), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT110), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G115), .A2(n880), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT47), .B(n865), .Z(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(n928) );
  XNOR2_X1 U967 ( .A(n868), .B(n928), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n870) );
  XNOR2_X1 U969 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U971 ( .A(n872), .B(n871), .Z(n890) );
  NAND2_X1 U972 ( .A1(G106), .A2(n873), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U975 ( .A(n877), .B(KEYINPUT45), .ZN(n885) );
  NAND2_X1 U976 ( .A1(n878), .A2(G130), .ZN(n879) );
  XOR2_X1 U977 ( .A(KEYINPUT107), .B(n879), .Z(n882) );
  NAND2_X1 U978 ( .A1(n880), .A2(G118), .ZN(n881) );
  NAND2_X1 U979 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U980 ( .A(KEYINPUT108), .B(n883), .Z(n884) );
  NAND2_X1 U981 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U982 ( .A(n886), .B(G164), .ZN(n887) );
  XOR2_X1 U983 ( .A(n888), .B(n887), .Z(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U985 ( .A(n918), .B(n891), .Z(n892) );
  XNOR2_X1 U986 ( .A(G162), .B(n892), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U988 ( .A1(G37), .A2(n895), .ZN(G395) );
  XOR2_X1 U989 ( .A(G2454), .B(G2435), .Z(n897) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2427), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n904) );
  XOR2_X1 U992 ( .A(KEYINPUT101), .B(G2446), .Z(n899) );
  XNOR2_X1 U993 ( .A(G2443), .B(G2430), .ZN(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n900), .B(G2451), .Z(n902) );
  XNOR2_X1 U996 ( .A(G1341), .B(G1348), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U998 ( .A(n904), .B(n903), .ZN(n905) );
  NAND2_X1 U999 ( .A1(n905), .A2(G14), .ZN(n906) );
  XOR2_X1 U1000 ( .A(KEYINPUT102), .B(n906), .Z(G401) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n907), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G397), .A2(n908), .ZN(n912) );
  NOR2_X1 U1004 ( .A1(n913), .A2(G401), .ZN(n909) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(n909), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(n910), .ZN(n911) );
  NAND2_X1 U1007 ( .A1(n912), .A2(n911), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(n913), .ZN(G319) );
  INV_X1 U1010 ( .A(G69), .ZN(G235) );
  INV_X1 U1011 ( .A(n914), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n924) );
  XOR2_X1 U1013 ( .A(G2084), .B(G160), .Z(n917) );
  NOR2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1015 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1017 ( .A1(n924), .A2(n923), .ZN(n935) );
  XOR2_X1 U1018 ( .A(G2090), .B(G162), .Z(n925) );
  NOR2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1020 ( .A(KEYINPUT51), .B(n927), .Z(n933) );
  XOR2_X1 U1021 ( .A(G2072), .B(n928), .Z(n930) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1024 ( .A(KEYINPUT50), .B(n931), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1026 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1027 ( .A(KEYINPUT52), .B(n936), .ZN(n938) );
  INV_X1 U1028 ( .A(KEYINPUT55), .ZN(n937) );
  NAND2_X1 U1029 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1030 ( .A1(n939), .A2(G29), .ZN(n1022) );
  XNOR2_X1 U1031 ( .A(G16), .B(KEYINPUT56), .ZN(n965) );
  XNOR2_X1 U1032 ( .A(G1961), .B(G301), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n963) );
  NOR2_X1 U1034 ( .A1(G166), .A2(n979), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n945) );
  NAND2_X1 U1036 ( .A1(n945), .A2(n944), .ZN(n948) );
  XOR2_X1 U1037 ( .A(G1956), .B(G299), .Z(n946) );
  XNOR2_X1 U1038 ( .A(KEYINPUT121), .B(n946), .ZN(n947) );
  NOR2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(KEYINPUT122), .B(n949), .ZN(n955) );
  XNOR2_X1 U1041 ( .A(n950), .B(G1341), .ZN(n953) );
  XNOR2_X1 U1042 ( .A(n951), .B(G1348), .ZN(n952) );
  NOR2_X1 U1043 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1044 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1045 ( .A(G1966), .B(KEYINPUT120), .Z(n956) );
  XNOR2_X1 U1046 ( .A(G168), .B(n956), .ZN(n958) );
  NOR2_X1 U1047 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1048 ( .A(KEYINPUT57), .B(n959), .ZN(n960) );
  NOR2_X1 U1049 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1050 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(n993) );
  INV_X1 U1052 ( .A(G16), .ZN(n991) );
  XNOR2_X1 U1053 ( .A(KEYINPUT59), .B(G1348), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(n966), .B(G4), .ZN(n971) );
  XOR2_X1 U1055 ( .A(G1341), .B(KEYINPUT123), .Z(n967) );
  XNOR2_X1 U1056 ( .A(G19), .B(n967), .ZN(n969) );
  XNOR2_X1 U1057 ( .A(G20), .B(G1956), .ZN(n968) );
  NOR2_X1 U1058 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1059 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1060 ( .A(KEYINPUT124), .B(G1981), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G6), .B(n972), .ZN(n973) );
  NOR2_X1 U1062 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1063 ( .A(KEYINPUT60), .B(n975), .Z(n977) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G21), .ZN(n976) );
  NOR2_X1 U1065 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1066 ( .A(KEYINPUT125), .B(n978), .Z(n986) );
  XOR2_X1 U1067 ( .A(G1986), .B(G24), .Z(n981) );
  XNOR2_X1 U1068 ( .A(n979), .B(G22), .ZN(n980) );
  NAND2_X1 U1069 ( .A1(n981), .A2(n980), .ZN(n983) );
  XNOR2_X1 U1070 ( .A(G23), .B(G1976), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NAND2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1074 ( .A(G5), .B(G1961), .ZN(n987) );
  NOR2_X1 U1075 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(KEYINPUT61), .B(n989), .ZN(n990) );
  NAND2_X1 U1077 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(n993), .A2(n992), .ZN(n1020) );
  XNOR2_X1 U1079 ( .A(G32), .B(n994), .ZN(n999) );
  XOR2_X1 U1080 ( .A(n995), .B(G27), .Z(n997) );
  XNOR2_X1 U1081 ( .A(G33), .B(G2072), .ZN(n996) );
  NOR2_X1 U1082 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1083 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XOR2_X1 U1084 ( .A(KEYINPUT117), .B(G2067), .Z(n1000) );
  XNOR2_X1 U1085 ( .A(G26), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1086 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1087 ( .A(KEYINPUT118), .B(n1003), .ZN(n1007) );
  XOR2_X1 U1088 ( .A(G25), .B(G1991), .Z(n1004) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(G28), .ZN(n1005) );
  XOR2_X1 U1090 ( .A(KEYINPUT116), .B(n1005), .Z(n1006) );
  NAND2_X1 U1091 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(n1008), .B(KEYINPUT53), .ZN(n1011) );
  XOR2_X1 U1093 ( .A(G2084), .B(G34), .Z(n1009) );
  XNOR2_X1 U1094 ( .A(KEYINPUT54), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1096 ( .A(G35), .B(G2090), .ZN(n1012) );
  NOR2_X1 U1097 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1098 ( .A(KEYINPUT55), .B(n1014), .ZN(n1016) );
  INV_X1 U1099 ( .A(G29), .ZN(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1101 ( .A1(n1017), .A2(G11), .ZN(n1018) );
  XOR2_X1 U1102 ( .A(KEYINPUT119), .B(n1018), .Z(n1019) );
  NOR2_X1 U1103 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1104 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  XOR2_X1 U1106 ( .A(KEYINPUT126), .B(G311), .Z(G150) );
endmodule

