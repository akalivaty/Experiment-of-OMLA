//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n620, new_n621, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147, new_n1149;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n464), .B2(G125), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI211_X1 g042(.A(KEYINPUT67), .B(G125), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n461), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n464), .A2(new_n472), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n471), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  AOI21_X1  g056(.A(new_n472), .B1(new_n462), .B2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n466), .A2(new_n467), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(G136), .B2(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n466), .B2(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n464), .A2(new_n494), .A3(new_n491), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n472), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n482), .A2(G126), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT68), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(new_n508), .A3(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n503), .A2(G651), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n513), .B1(new_n504), .B2(new_n506), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(new_n508), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G50), .A2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  XOR2_X1   g096(.A(KEYINPUT70), .B(G88), .Z(new_n522));
  OAI21_X1  g097(.A(new_n517), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n520), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(new_n513), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n512), .B2(new_n515), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n510), .B1(new_n514), .B2(new_n508), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT68), .B(KEYINPUT6), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT69), .B1(new_n532), .B2(new_n513), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n531), .A2(KEYINPUT71), .A3(new_n533), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n530), .A2(G51), .A3(new_n534), .A4(G543), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n531), .A2(G89), .A3(new_n520), .A4(new_n533), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(KEYINPUT7), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n538), .A2(new_n539), .B1(new_n520), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n535), .A2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  INV_X1    g119(.A(G543), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n531), .A2(new_n533), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n529), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n547), .A2(new_n534), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G52), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n521), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n521), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n550), .A2(G90), .B1(G651), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(new_n548), .A2(G43), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n521), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n550), .A2(G81), .B1(G651), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT72), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n557), .A2(new_n564), .A3(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  AOI22_X1  g147(.A1(new_n520), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n513), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n574), .B1(new_n550), .B2(G91), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n548), .A2(G53), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n547), .A2(new_n534), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI211_X1 g155(.A(KEYINPUT73), .B(KEYINPUT9), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n576), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G299));
  AND3_X1   g158(.A1(new_n549), .A2(KEYINPUT74), .A3(new_n554), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT74), .B1(new_n549), .B2(new_n554), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n584), .A2(new_n585), .ZN(G301));
  NAND2_X1  g161(.A1(new_n548), .A2(G49), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT75), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n516), .A2(new_n520), .ZN(new_n589));
  INV_X1    g164(.A(G87), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n550), .A2(KEYINPUT75), .A3(G87), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n587), .A2(new_n593), .A3(new_n594), .ZN(G288));
  NAND3_X1  g170(.A1(new_n516), .A2(G48), .A3(G543), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT76), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n520), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n513), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n550), .B2(G86), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(G305));
  NAND2_X1  g176(.A1(new_n548), .A2(G47), .ZN(new_n602));
  NAND2_X1  g177(.A1(G72), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n521), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n550), .A2(G85), .B1(G651), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n602), .A2(new_n606), .ZN(G290));
  NAND2_X1  g182(.A1(new_n550), .A2(G92), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n520), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n610), .A2(new_n513), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n548), .A2(G54), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n614), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g190(.A(new_n614), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(new_n582), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(new_n582), .B2(G868), .ZN(G280));
  AND2_X1   g194(.A1(new_n612), .A2(new_n613), .ZN(new_n620));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(G860), .ZN(G148));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n566), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n614), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n488), .A2(G135), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT77), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n482), .A2(G123), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n472), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT78), .Z(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n464), .A2(new_n474), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT13), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2100), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2443), .B(G2446), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT80), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n651), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT81), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT84), .B(KEYINPUT17), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n663), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n661), .ZN(new_n668));
  INV_X1    g243(.A(new_n663), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n669), .A2(KEYINPUT83), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(KEYINPUT83), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(new_n662), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n668), .A2(new_n663), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT87), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n689), .B1(new_n684), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(new_n691), .B2(new_n684), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n693), .A2(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n693), .A2(KEYINPUT20), .ZN(new_n695));
  OAI221_X1 g270(.A(new_n690), .B1(new_n689), .B2(new_n685), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1981), .B(G1986), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(G229));
  NAND2_X1  g278(.A1(new_n482), .A2(G119), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n472), .A2(G107), .ZN(new_n705));
  OAI21_X1  g280(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n706));
  INV_X1    g281(.A(G131), .ZN(new_n707));
  OAI221_X1 g282(.A(new_n704), .B1(new_n705), .B2(new_n706), .C1(new_n707), .C2(new_n476), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT88), .B(G29), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n709), .S(new_n711), .Z(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT90), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT35), .B(G1991), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n714), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G23), .ZN(new_n719));
  INV_X1    g294(.A(G288), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(new_n718), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT33), .B(G1976), .Z(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  OR2_X1    g299(.A1(G6), .A2(G16), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G305), .B2(new_n718), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT32), .B(G1981), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n718), .A2(G22), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT92), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G303), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(G1971), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n726), .B2(new_n728), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n723), .A2(new_n724), .A3(new_n729), .A4(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(KEYINPUT34), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(KEYINPUT34), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G24), .ZN(new_n739));
  INV_X1    g314(.A(G290), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n739), .B1(new_n740), .B2(G16), .ZN(new_n741));
  INV_X1    g316(.A(G1986), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n717), .A2(new_n737), .A3(new_n738), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n744), .B(new_n745), .Z(new_n746));
  NOR2_X1   g321(.A1(G171), .A2(new_n718), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G5), .B2(new_n718), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT97), .ZN(new_n751));
  INV_X1    g326(.A(G29), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G33), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT25), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G139), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n476), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n472), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n752), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G2072), .Z(new_n763));
  INV_X1    g338(.A(G2084), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT24), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G34), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G34), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n710), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n480), .B2(new_n752), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n752), .A2(G32), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT26), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G129), .B2(new_n482), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n488), .A2(G141), .B1(G105), .B2(new_n474), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n770), .B1(new_n776), .B2(new_n752), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT95), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT27), .B(G1996), .Z(new_n779));
  OAI221_X1 g354(.A(new_n763), .B1(new_n764), .B2(new_n769), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT96), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n634), .A2(new_n710), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n710), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n710), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(G28), .ZN(new_n788));
  OR2_X1    g363(.A1(new_n788), .A2(KEYINPUT30), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n788), .B2(KEYINPUT30), .ZN(new_n790));
  OR2_X1    g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  NAND2_X1  g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n789), .A2(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n786), .A2(new_n787), .A3(new_n793), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n778), .A2(new_n779), .B1(new_n764), .B2(new_n769), .ZN(new_n795));
  AND3_X1   g370(.A1(new_n782), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n718), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G168), .B2(new_n718), .ZN(new_n798));
  INV_X1    g373(.A(G1966), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n748), .A2(new_n749), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n781), .A2(new_n796), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n751), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT98), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n803), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n620), .A2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G4), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1348), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n710), .A2(G26), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT28), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n488), .A2(G140), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n482), .A2(G128), .ZN(new_n815));
  OR2_X1    g390(.A1(G104), .A2(G2105), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n816), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(new_n752), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT94), .ZN(new_n821));
  INV_X1    g396(.A(G2067), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n711), .A2(G35), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G162), .B2(new_n711), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT29), .B(G2090), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NOR4_X1   g402(.A1(new_n810), .A2(new_n811), .A3(new_n823), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n718), .A2(G20), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT23), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n582), .B2(new_n718), .ZN(new_n831));
  INV_X1    g406(.A(G1956), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n718), .A2(G19), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n567), .B2(new_n718), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(G1341), .Z(new_n836));
  NAND3_X1  g411(.A1(new_n828), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n805), .A2(new_n806), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n746), .A2(new_n838), .ZN(G150));
  INV_X1    g414(.A(G150), .ZN(G311));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n621), .ZN(new_n841));
  XNOR2_X1  g416(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n550), .A2(G93), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT100), .B(G55), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n844), .B1(new_n513), .B2(new_n845), .C1(new_n579), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n566), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n562), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n843), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(new_n852), .B2(new_n851), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n847), .A2(G860), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT101), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n634), .B(new_n480), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G162), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n761), .B(new_n775), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n708), .B(new_n638), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n818), .B(new_n501), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n488), .A2(G142), .B1(G130), .B2(new_n482), .ZN(new_n865));
  OAI21_X1  g440(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n867));
  INV_X1    g442(.A(G118), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n866), .A2(new_n867), .B1(new_n868), .B2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n869), .B1(new_n867), .B2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n864), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n863), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT103), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n875), .B(new_n876), .C1(new_n860), .C2(new_n873), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g453(.A(KEYINPUT42), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n850), .A2(new_n625), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n848), .B(new_n849), .C1(G559), .C2(new_n614), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n620), .A2(new_n582), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n614), .A2(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n880), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n880), .A2(new_n881), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n879), .B(new_n885), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n887), .A2(new_n888), .B1(new_n880), .B2(new_n881), .ZN(new_n892));
  INV_X1    g467(.A(new_n885), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT42), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(G290), .B(G166), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n891), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n891), .B2(new_n894), .ZN(new_n899));
  OAI21_X1  g474(.A(G868), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n847), .A2(new_n623), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n901), .B1(new_n900), .B2(new_n902), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(G295));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n902), .ZN(G331));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n584), .A2(new_n585), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(G168), .ZN(new_n909));
  NOR2_X1   g484(.A1(G171), .A2(G168), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n850), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(G301), .A2(G286), .ZN(new_n913));
  OAI211_X1 g488(.A(new_n848), .B(new_n849), .C1(new_n913), .C2(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n884), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n887), .A2(new_n888), .A3(new_n912), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT106), .B1(new_n919), .B2(new_n897), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  INV_X1    g496(.A(new_n897), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n917), .A2(new_n918), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n897), .B(KEYINPUT105), .ZN(new_n926));
  AOI21_X1  g501(.A(G37), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n925), .B1(new_n924), .B2(new_n927), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n907), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n924), .A2(new_n927), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(KEYINPUT44), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(G397));
  AOI21_X1  g510(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(KEYINPUT45), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(G40), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n470), .B2(G2105), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n740), .A2(new_n742), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n818), .B(new_n822), .ZN(new_n944));
  INV_X1    g519(.A(G1996), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n775), .B(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n708), .B(new_n715), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n943), .A2(new_n944), .A3(new_n946), .A4(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n740), .A2(new_n742), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n942), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(G286), .B2(G8), .ZN(new_n952));
  INV_X1    g527(.A(G8), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT114), .B(new_n953), .C1(new_n535), .C2(new_n542), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n956), .A2(G1384), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n958), .B1(new_n496), .B2(new_n500), .ZN(new_n959));
  OAI22_X1  g534(.A1(KEYINPUT109), .A2(new_n959), .B1(new_n936), .B2(KEYINPUT45), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n501), .A2(KEYINPUT109), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n940), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n799), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n501), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n936), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n764), .A3(new_n940), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n953), .B1(new_n963), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT115), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n955), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g547(.A(KEYINPUT115), .B(new_n953), .C1(new_n963), .C2(new_n969), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT51), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT116), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT116), .ZN(new_n976));
  OAI211_X1 g551(.A(new_n976), .B(KEYINPUT51), .C1(new_n972), .C2(new_n973), .ZN(new_n977));
  INV_X1    g552(.A(new_n955), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n978), .A2(KEYINPUT51), .A3(new_n970), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n975), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n955), .B1(new_n963), .B2(new_n969), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT117), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT62), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT117), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n981), .A2(new_n987), .A3(new_n983), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n941), .A2(new_n965), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n953), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT76), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n596), .B(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n600), .ZN(new_n995));
  OAI21_X1  g570(.A(G1981), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n597), .A2(new_n997), .A3(new_n600), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n992), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n998), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n991), .B1(G288), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1003), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1001), .A2(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1004), .A2(KEYINPUT52), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT107), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT107), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(new_n1010), .A3(KEYINPUT52), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n959), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n938), .A2(new_n785), .A3(new_n940), .A4(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1016));
  NAND3_X1  g591(.A1(new_n966), .A2(new_n940), .A3(new_n968), .ZN(new_n1017));
  AOI22_X1  g592(.A1(new_n1015), .A2(new_n1016), .B1(new_n1017), .B2(new_n749), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n785), .A2(KEYINPUT53), .ZN(new_n1019));
  OR3_X1    g594(.A1(new_n960), .A2(new_n962), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(G166), .B2(new_n953), .ZN(new_n1023));
  NAND3_X1  g598(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n1026));
  AOI21_X1  g601(.A(G2090), .B1(new_n1017), .B2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1027), .B1(new_n1026), .B2(new_n1017), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n937), .A2(new_n959), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n940), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n733), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1025), .B1(new_n1032), .B2(G8), .ZN(new_n1033));
  OR2_X1    g608(.A1(new_n1017), .A2(G2090), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n953), .B1(new_n1034), .B2(new_n1031), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(new_n1025), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  AND4_X1   g612(.A1(new_n908), .A2(new_n1013), .A3(new_n1021), .A4(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n989), .A2(KEYINPUT123), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n979), .B1(new_n974), .B2(KEYINPUT116), .ZN(new_n1040));
  AOI211_X1 g615(.A(KEYINPUT117), .B(new_n982), .C1(new_n1040), .C2(new_n977), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n987), .B1(new_n981), .B2(new_n983), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT62), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT123), .B1(new_n989), .B2(new_n1038), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n939), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n470), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(G2105), .B1(new_n470), .B2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT120), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1019), .ZN(new_n1054));
  OAI211_X1 g629(.A(KEYINPUT120), .B(new_n1047), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1053), .A2(new_n1029), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1018), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G171), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(KEYINPUT54), .C1(new_n908), .C2(new_n1021), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1037), .A2(new_n1007), .A3(new_n1012), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(G301), .A2(new_n1018), .A3(new_n1056), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n1061), .A2(KEYINPUT121), .B1(new_n1021), .B2(new_n908), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n1057), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT54), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1060), .A2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT61), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1017), .A2(new_n832), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1030), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1075));
  AOI211_X1 g650(.A(KEYINPUT57), .B(new_n576), .C1(new_n578), .C2(new_n581), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n582), .A2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1080), .A2(new_n1076), .A3(new_n1073), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1069), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1075), .A2(new_n1077), .A3(new_n1074), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1073), .B1(new_n1080), .B2(new_n1076), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT61), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT110), .B(KEYINPUT58), .Z(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(G1341), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1030), .A2(G1996), .B1(new_n990), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n563), .A2(new_n1088), .A3(KEYINPUT111), .A4(new_n565), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT59), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1082), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(KEYINPUT112), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT112), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1082), .A2(new_n1093), .A3(new_n1085), .A4(new_n1090), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1017), .A2(new_n809), .B1(new_n990), .B2(new_n822), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT60), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT113), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(new_n614), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1099), .A2(new_n1100), .B1(KEYINPUT60), .B2(new_n1095), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1092), .A2(new_n1094), .A3(new_n1101), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n614), .A2(new_n1095), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1083), .B1(new_n1078), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1065), .B(KEYINPUT122), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1068), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n970), .A2(G168), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1033), .A2(KEYINPUT63), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1013), .B1(new_n1036), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(G1976), .B(G288), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1111));
  INV_X1    g686(.A(new_n998), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n991), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  AND2_X1   g689(.A1(new_n970), .A2(G168), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1013), .B(new_n1115), .C1(new_n1025), .C2(new_n1035), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1114), .B1(KEYINPUT63), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1107), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n950), .B1(new_n1046), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n942), .A2(new_n945), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT46), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  XNOR2_X1  g697(.A(new_n1122), .B(KEYINPUT124), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n944), .A2(new_n776), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1120), .A2(new_n1121), .B1(new_n1124), .B2(new_n942), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT47), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n709), .A2(new_n716), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(new_n944), .A3(new_n946), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(G2067), .B2(new_n818), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n942), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n740), .A2(new_n742), .A3(new_n942), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1132), .B(KEYINPUT125), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT48), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n946), .A2(new_n944), .A3(new_n947), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n942), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1127), .B(new_n1131), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT126), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1119), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g717(.A(new_n658), .ZN(new_n1144));
  INV_X1    g718(.A(G319), .ZN(new_n1145));
  NOR3_X1   g719(.A1(new_n1144), .A2(new_n1145), .A3(G227), .ZN(new_n1146));
  NAND3_X1  g720(.A1(new_n877), .A2(new_n702), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g721(.A(new_n1147), .B1(new_n933), .B2(new_n928), .ZN(G308));
  NAND2_X1  g722(.A1(new_n933), .A2(new_n928), .ZN(new_n1149));
  NAND4_X1  g723(.A1(new_n1149), .A2(new_n702), .A3(new_n877), .A4(new_n1146), .ZN(G225));
endmodule


