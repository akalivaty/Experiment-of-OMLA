//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  XOR2_X1   g000(.A(G43gat), .B(G50gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n204), .A2(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  OR3_X1    g009(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(KEYINPUT89), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n212), .B1(KEYINPUT89), .B2(new_n211), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT88), .ZN(new_n214));
  AND3_X1   g013(.A1(new_n202), .A2(new_n214), .A3(new_n203), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(new_n202), .B2(new_n203), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n208), .B(new_n213), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n211), .A2(new_n209), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n204), .B1(new_n218), .B2(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT17), .ZN(new_n221));
  XNOR2_X1  g020(.A(G15gat), .B(G22gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(G1gat), .ZN(new_n224));
  INV_X1    g023(.A(G8gat), .ZN(new_n225));
  OAI221_X1 g024(.A(new_n224), .B1(KEYINPUT90), .B2(new_n225), .C1(G1gat), .C2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n220), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT18), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n232), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n228), .B(new_n220), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n231), .B(KEYINPUT13), .Z(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n236), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G141gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(G197gat), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT11), .B(G169gat), .Z(new_n243));
  XNOR2_X1  g042(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(new_n244), .B(KEYINPUT12), .Z(new_n245));
  NAND2_X1  g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n235), .A2(new_n236), .A3(new_n247), .A4(new_n239), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G228gat), .A2(G233gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n252));
  XOR2_X1   g051(.A(G197gat), .B(G204gat), .Z(new_n253));
  AOI21_X1  g052(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  OR2_X1    g058(.A1(new_n255), .A2(new_n256), .ZN(new_n260));
  AND2_X1   g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n252), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265));
  INV_X1    g064(.A(G155gat), .ZN(new_n266));
  INV_X1    g065(.A(G162gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(KEYINPUT2), .ZN(new_n269));
  INV_X1    g068(.A(G141gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(G148gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(G148gat), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n271), .B1(new_n272), .B2(KEYINPUT80), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT80), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n274), .A2(new_n270), .A3(G148gat), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n269), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G141gat), .B(G148gat), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n265), .B(new_n268), .C1(new_n277), .C2(KEYINPUT2), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n264), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n256), .B1(new_n255), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n281), .B2(new_n255), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n259), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n276), .A2(new_n252), .A3(new_n278), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n262), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT83), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n280), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n251), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n284), .B(KEYINPUT76), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n251), .B1(new_n294), .B2(new_n287), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n252), .B1(new_n285), .B2(KEYINPUT29), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n279), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n293), .A2(new_n298), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  XNOR2_X1  g101(.A(G78gat), .B(G106gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT31), .B(G50gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n293), .A2(new_n298), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n299), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT85), .ZN(new_n309));
  INV_X1    g108(.A(G22gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n305), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n293), .B(new_n298), .C1(new_n309), .C2(new_n310), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n302), .A2(new_n308), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  OR2_X1    g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(KEYINPUT66), .B2(KEYINPUT23), .ZN(new_n318));
  AND2_X1   g117(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT67), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n316), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  INV_X1    g123(.A(G183gat), .ZN(new_n325));
  INV_X1    g124(.A(G190gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(KEYINPUT68), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(KEYINPUT68), .B2(new_n327), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n330));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI221_X1 g132(.A(new_n320), .B1(new_n321), .B2(new_n323), .C1(new_n329), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT25), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n316), .A2(KEYINPUT26), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n317), .B(new_n336), .C1(new_n323), .C2(KEYINPUT26), .ZN(new_n337));
  NAND2_X1  g136(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n338));
  AOI21_X1  g137(.A(G190gat), .B1(new_n338), .B2(KEYINPUT27), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT28), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(KEYINPUT27), .B(G183gat), .Z(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  NOR3_X1   g143(.A1(new_n343), .A2(new_n344), .A3(G190gat), .ZN(new_n345));
  OAI221_X1 g144(.A(new_n337), .B1(new_n325), .B2(new_n326), .C1(new_n342), .C2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n332), .B1(KEYINPUT24), .B2(new_n327), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT65), .B(G169gat), .ZN(new_n349));
  INV_X1    g148(.A(G176gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(KEYINPUT23), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n347), .A2(new_n348), .A3(new_n320), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n346), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n315), .B1(new_n353), .B2(new_n262), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT78), .B1(new_n353), .B2(new_n315), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n356), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n294), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n315), .B1(new_n353), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n353), .B2(new_n315), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(new_n284), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n358), .A2(new_n294), .B1(new_n284), .B2(new_n362), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT30), .A3(new_n367), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AND3_X1   g171(.A1(new_n359), .A2(new_n363), .A3(new_n367), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n367), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT79), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n372), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G113gat), .B(G120gat), .Z(new_n380));
  INV_X1    g179(.A(KEYINPUT71), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n383));
  XNOR2_X1  g182(.A(G127gat), .B(G134gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT71), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n382), .A2(new_n383), .A3(new_n384), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(KEYINPUT70), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT70), .ZN(new_n389));
  INV_X1    g188(.A(G134gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(G127gat), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n388), .B(new_n391), .C1(KEYINPUT1), .C2(new_n385), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(new_n279), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n397), .A2(new_n393), .A3(new_n286), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(G225gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n393), .B(new_n279), .Z(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n400), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(KEYINPUT39), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(G1gat), .B(G29gat), .Z(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT82), .ZN(new_n407));
  XOR2_X1   g206(.A(G57gat), .B(G85gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n407), .B(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(KEYINPUT86), .A2(KEYINPUT39), .ZN(new_n413));
  NAND2_X1  g212(.A1(KEYINPUT86), .A2(KEYINPUT39), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n399), .A2(new_n401), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n405), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT40), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT5), .B1(new_n403), .B2(new_n400), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n399), .B2(new_n401), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n396), .A2(KEYINPUT5), .A3(new_n400), .A4(new_n398), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n411), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n416), .A2(new_n417), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n418), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n314), .B1(new_n379), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n368), .B1(new_n364), .B2(KEYINPUT37), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n370), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT38), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT87), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n420), .A2(new_n421), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT6), .B1(new_n431), .B2(new_n412), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n422), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n420), .A2(KEYINPUT6), .A3(new_n411), .A4(new_n421), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n376), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n426), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n358), .A2(new_n294), .B1(new_n284), .B2(new_n362), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT38), .B1(new_n437), .B2(KEYINPUT37), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n435), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n440), .B(KEYINPUT38), .C1(new_n426), .C2(new_n428), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n430), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n353), .A2(new_n393), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT73), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT73), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n353), .A2(new_n445), .A3(new_n393), .ZN(new_n446));
  INV_X1    g245(.A(new_n393), .ZN(new_n447));
  NAND4_X1  g246(.A1(new_n335), .A2(new_n447), .A3(new_n346), .A4(new_n352), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n448), .A2(KEYINPUT72), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(KEYINPUT72), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n444), .A2(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(G227gat), .ZN(new_n452));
  INV_X1    g251(.A(G233gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT64), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT32), .B1(new_n451), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n458), .B1(new_n451), .B2(new_n456), .ZN(new_n459));
  XOR2_X1   g258(.A(G15gat), .B(G43gat), .Z(new_n460));
  XNOR2_X1  g259(.A(G71gat), .B(G99gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n454), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n451), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n465), .A2(KEYINPUT34), .B1(new_n451), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n462), .ZN(new_n468));
  OAI221_X1 g267(.A(KEYINPUT32), .B1(new_n458), .B2(new_n468), .C1(new_n451), .C2(new_n456), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n463), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n467), .B1(new_n463), .B2(new_n469), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT36), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT36), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(new_n470), .B2(new_n471), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n425), .A2(new_n442), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n433), .A2(new_n434), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n372), .B(new_n477), .C1(new_n375), .C2(new_n378), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n314), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n369), .A2(new_n371), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n374), .B1(new_n373), .B2(KEYINPUT30), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n376), .A2(KEYINPUT79), .A3(new_n377), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n308), .A2(new_n302), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n312), .A2(new_n313), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n472), .A2(new_n477), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n314), .A2(new_n470), .A3(new_n471), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT35), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n490), .A2(new_n491), .A3(new_n477), .A4(new_n484), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n250), .B1(new_n480), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT7), .ZN(new_n496));
  NOR2_X1   g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT8), .ZN(new_n498));
  NAND2_X1  g297(.A1(G99gat), .A2(G106gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(KEYINPUT96), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(G99gat), .A3(G106gat), .ZN(new_n502));
  AOI211_X1 g301(.A(KEYINPUT97), .B(new_n497), .C1(new_n500), .C2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT97), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n499), .A2(KEYINPUT96), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n505), .A2(new_n502), .A3(KEYINPUT8), .ZN(new_n506));
  INV_X1    g305(.A(new_n497), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n496), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G99gat), .B(G106gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n510), .B(new_n496), .C1(new_n503), .C2(new_n508), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n512), .A2(KEYINPUT98), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n506), .A2(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT97), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n506), .A2(new_n504), .A3(new_n507), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n510), .B1(new_n519), .B2(new_n496), .ZN(new_n520));
  INV_X1    g319(.A(new_n513), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n221), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n512), .A2(KEYINPUT98), .A3(new_n513), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT98), .B1(new_n512), .B2(new_n513), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n220), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n529), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n523), .A2(new_n531), .A3(new_n526), .A4(new_n527), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n532), .A2(KEYINPUT99), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(KEYINPUT99), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT100), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n536), .B1(new_n533), .B2(new_n534), .ZN(new_n537));
  XNOR2_X1  g336(.A(G134gat), .B(G162gat), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n540), .ZN(new_n542));
  OAI221_X1 g341(.A(new_n530), .B1(new_n536), .B2(new_n542), .C1(new_n533), .C2(new_n534), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(G183gat), .B(G211gat), .Z(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G64gat), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(G57gat), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n548), .A2(KEYINPUT93), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(G57gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(KEYINPUT93), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(G71gat), .B(G78gat), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(G57gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G64gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n550), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n554), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n550), .A3(KEYINPUT91), .ZN(new_n562));
  AOI211_X1 g361(.A(KEYINPUT92), .B(new_n553), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n557), .A2(G64gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n560), .B1(new_n548), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n562), .A3(new_n555), .ZN(new_n567));
  INV_X1    g366(.A(new_n553), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n556), .B1(new_n563), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n572));
  OR3_X1    g371(.A1(new_n571), .A2(KEYINPUT95), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT95), .B1(new_n571), .B2(new_n572), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n578), .A3(new_n574), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n546), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n546), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n229), .B1(new_n584), .B2(new_n570), .ZN(new_n585));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(G231gat), .A2(G233gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n585), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n583), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n570), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n524), .B2(new_n525), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n570), .B1(new_n520), .B2(new_n521), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n555), .B1(new_n598), .B2(KEYINPUT91), .ZN(new_n599));
  INV_X1    g398(.A(new_n562), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n568), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT92), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n567), .A2(new_n564), .A3(new_n568), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n604), .A2(new_n512), .A3(new_n513), .A4(new_n556), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n597), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n593), .B1(new_n596), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n592), .B1(new_n597), .B2(new_n605), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G120gat), .B(G148gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT102), .ZN(new_n612));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n608), .A2(new_n609), .A3(new_n614), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n544), .A2(new_n591), .A3(new_n618), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(KEYINPUT103), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n494), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n477), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g426(.A(KEYINPUT16), .B(G8gat), .Z(new_n628));
  NAND3_X1  g427(.A1(new_n624), .A2(new_n379), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(G8gat), .B1(new_n623), .B2(new_n484), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  MUX2_X1   g430(.A(new_n629), .B(new_n631), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g431(.A(G15gat), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n473), .A2(new_n475), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n623), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n472), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n623), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n637), .A2(KEYINPUT104), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(KEYINPUT104), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(G1326gat));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n487), .ZN(new_n641));
  XOR2_X1   g440(.A(KEYINPUT43), .B(G22gat), .Z(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n618), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n591), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n544), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT105), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n494), .A2(new_n205), .A3(new_n625), .A4(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT45), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n425), .A2(new_n442), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n479), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n478), .A2(KEYINPUT106), .A3(new_n314), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n651), .A2(new_n653), .A3(new_n634), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n493), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n646), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n480), .A2(new_n493), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n544), .A2(new_n658), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n657), .A2(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n645), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(new_n250), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n664), .A2(new_n625), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n650), .B1(new_n665), .B2(new_n205), .ZN(G1328gat));
  NAND2_X1  g465(.A1(new_n494), .A2(new_n648), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(G36gat), .A3(new_n484), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n664), .A2(new_n379), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n670), .B1(new_n671), .B2(new_n206), .ZN(G1329gat));
  INV_X1    g471(.A(new_n634), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n661), .A2(G43gat), .A3(new_n673), .A4(new_n663), .ZN(new_n674));
  INV_X1    g473(.A(G43gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n675), .B1(new_n667), .B2(new_n636), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT48), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n682));
  INV_X1    g481(.A(new_n654), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT106), .B1(new_n478), .B2(new_n314), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(new_n476), .B1(new_n489), .B2(new_n492), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n658), .B1(new_n686), .B2(new_n544), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n659), .A2(new_n660), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n314), .A4(new_n663), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G50gat), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n667), .A2(G50gat), .A3(new_n487), .ZN(new_n691));
  AOI211_X1 g490(.A(new_n681), .B(new_n682), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  AND4_X1   g491(.A1(new_n679), .A2(new_n690), .A3(new_n680), .A4(new_n691), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(G1331gat));
  NOR2_X1   g493(.A1(new_n583), .A2(new_n590), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n589), .B1(new_n581), .B2(new_n582), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR4_X1   g496(.A1(new_n646), .A2(new_n249), .A3(new_n697), .A4(new_n618), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n656), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n477), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(new_n557), .ZN(G1332gat));
  AOI211_X1 g500(.A(new_n484), .B(new_n699), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n702));
  NOR2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1333gat));
  NOR3_X1   g503(.A1(new_n699), .A2(G71gat), .A3(new_n636), .ZN(new_n705));
  INV_X1    g504(.A(new_n699), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n673), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(G71gat), .B2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g508(.A1(new_n706), .A2(new_n314), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n591), .A2(new_n249), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n618), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n661), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n625), .ZN(new_n716));
  INV_X1    g515(.A(G85gat), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n656), .A2(new_n646), .A3(new_n712), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT51), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n656), .A2(KEYINPUT51), .A3(new_n646), .A4(new_n712), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n644), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n625), .A2(new_n717), .ZN(new_n724));
  OAI22_X1  g523(.A1(new_n716), .A2(new_n717), .B1(new_n723), .B2(new_n724), .ZN(G1336gat));
  INV_X1    g524(.A(KEYINPUT110), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n720), .A2(new_n726), .A3(new_n721), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n484), .A2(G92gat), .A3(new_n618), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT109), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n718), .A2(KEYINPUT110), .A3(new_n719), .ZN(new_n730));
  AND3_X1   g529(.A1(new_n727), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n687), .A2(new_n688), .A3(new_n379), .A4(new_n714), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n732), .A2(G92gat), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT52), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT52), .B1(new_n722), .B2(new_n729), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(KEYINPUT111), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n732), .A2(KEYINPUT111), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n734), .A2(new_n739), .ZN(G1337gat));
  AND2_X1   g539(.A1(new_n715), .A2(new_n673), .ZN(new_n741));
  INV_X1    g540(.A(G99gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n472), .A2(new_n742), .ZN(new_n743));
  OAI22_X1  g542(.A1(new_n741), .A2(new_n742), .B1(new_n723), .B2(new_n743), .ZN(G1338gat));
  NOR3_X1   g543(.A1(new_n487), .A2(G106gat), .A3(new_n618), .ZN(new_n745));
  XOR2_X1   g544(.A(new_n745), .B(KEYINPUT112), .Z(new_n746));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n730), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n687), .A2(new_n688), .A3(new_n314), .A4(new_n714), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G106gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT53), .B1(new_n722), .B2(new_n745), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1339gat));
  NOR2_X1   g553(.A1(KEYINPUT117), .A2(G113gat), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n608), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(KEYINPUT55), .A3(new_n614), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n597), .A2(new_n605), .A3(new_n606), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n556), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n760), .B1(new_n522), .B2(new_n514), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n592), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n596), .A2(new_n607), .A3(new_n593), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(KEYINPUT54), .A3(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n596), .A2(new_n607), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n756), .B1(new_n767), .B2(new_n592), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(KEYINPUT114), .A3(new_n763), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n758), .B1(new_n766), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n617), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n614), .ZN(new_n773));
  INV_X1    g572(.A(new_n773), .ZN(new_n774));
  AND4_X1   g573(.A1(KEYINPUT114), .A2(new_n762), .A3(KEYINPUT54), .A4(new_n763), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT114), .B1(new_n768), .B2(new_n763), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n775), .A2(new_n776), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT115), .B1(new_n780), .B2(new_n758), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n772), .A2(new_n779), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n772), .A2(new_n781), .A3(KEYINPUT116), .A4(new_n779), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n249), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n237), .A2(new_n238), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n244), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n248), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n644), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n646), .B1(new_n786), .B2(new_n791), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n541), .A2(new_n543), .A3(new_n790), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n793), .A3(new_n785), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n697), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n697), .B1(new_n543), .B2(new_n541), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n797), .A2(new_n798), .A3(new_n250), .A4(new_n618), .ZN(new_n799));
  OAI21_X1  g598(.A(KEYINPUT113), .B1(new_n619), .B2(new_n249), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n477), .B1(new_n796), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n490), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n379), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n755), .B1(new_n806), .B2(new_n249), .ZN(new_n807));
  NAND2_X1  g606(.A1(KEYINPUT117), .A2(G113gat), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n807), .B(new_n808), .Z(G1340gat));
  NOR2_X1   g608(.A1(KEYINPUT118), .A2(G120gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n810), .B1(new_n806), .B2(new_n644), .ZN(new_n811));
  NAND2_X1  g610(.A1(KEYINPUT118), .A2(G120gat), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n811), .B(new_n812), .Z(G1341gat));
  NAND2_X1  g612(.A1(new_n806), .A2(new_n591), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(G127gat), .ZN(G1342gat));
  NAND4_X1  g614(.A1(new_n803), .A2(new_n390), .A3(new_n805), .A4(new_n646), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(KEYINPUT119), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n646), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G134gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n817), .A2(KEYINPUT56), .A3(new_n818), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(G1343gat));
  NOR2_X1   g624(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n484), .A2(new_n625), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n673), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n796), .A2(new_n802), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n830), .B2(new_n314), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n487), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n773), .B1(new_n766), .B2(new_n769), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT120), .B1(new_n834), .B2(KEYINPUT55), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n777), .A2(new_n836), .A3(new_n778), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n837), .A3(new_n249), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n772), .A2(new_n781), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n791), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n544), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n591), .B1(new_n841), .B2(new_n794), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n833), .B1(new_n842), .B2(new_n801), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT121), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845));
  OAI211_X1 g644(.A(new_n845), .B(new_n833), .C1(new_n842), .C2(new_n801), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n249), .B(new_n829), .C1(new_n831), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(G141gat), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n673), .A2(new_n487), .A3(new_n379), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n250), .A2(G141gat), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n830), .A2(new_n625), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n827), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n826), .B(new_n854), .C1(new_n848), .C2(G141gat), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(G1344gat));
  AND2_X1   g657(.A1(new_n803), .A2(new_n850), .ZN(new_n859));
  INV_X1    g658(.A(G148gat), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n644), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(G148gat), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n829), .B1(new_n831), .B2(new_n847), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n865), .B2(new_n644), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n620), .A2(new_n621), .A3(new_n249), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n793), .A2(new_n779), .A3(new_n781), .A4(new_n772), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n591), .B1(new_n841), .B2(new_n868), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n832), .B(new_n314), .C1(new_n867), .C2(new_n869), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n673), .A2(new_n618), .A3(new_n828), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n487), .B1(new_n796), .B2(new_n802), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n832), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n862), .B1(new_n873), .B2(G148gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n861), .B1(new_n866), .B2(new_n874), .ZN(G1345gat));
  OAI21_X1  g674(.A(G155gat), .B1(new_n864), .B2(new_n697), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n266), .A3(new_n591), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n859), .B2(new_n646), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n544), .A2(new_n267), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n865), .B2(new_n880), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n484), .A2(new_n625), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n804), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n830), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n250), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n830), .A2(KEYINPUT123), .A3(new_n884), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT123), .B1(new_n830), .B2(new_n884), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n249), .A2(new_n349), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1348gat));
  NOR3_X1   g690(.A1(new_n885), .A2(new_n350), .A3(new_n618), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  OAI211_X1 g692(.A(new_n893), .B(new_n350), .C1(new_n889), .C2(new_n618), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n887), .A2(new_n888), .A3(new_n618), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT124), .B1(new_n895), .B2(G176gat), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n892), .B1(new_n894), .B2(new_n896), .ZN(G1349gat));
  OAI21_X1  g696(.A(new_n325), .B1(new_n885), .B2(new_n697), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n830), .A2(new_n343), .A3(new_n591), .A4(new_n884), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XOR2_X1   g699(.A(new_n900), .B(KEYINPUT60), .Z(G1350gat));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n902));
  OAI221_X1 g701(.A(G190gat), .B1(KEYINPUT125), .B2(new_n902), .C1(new_n885), .C2(new_n544), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(KEYINPUT125), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n889), .A2(G190gat), .A3(new_n544), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1351gat));
  NOR2_X1   g706(.A1(new_n673), .A2(new_n883), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n870), .B(new_n908), .C1(new_n872), .C2(new_n832), .ZN(new_n909));
  OAI21_X1  g708(.A(G197gat), .B1(new_n909), .B2(new_n250), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n872), .A2(new_n908), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n250), .A2(G197gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT126), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n910), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1352gat));
  INV_X1    g717(.A(G204gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n911), .A2(new_n919), .A3(new_n644), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n921));
  OAI21_X1  g720(.A(G204gat), .B1(new_n909), .B2(new_n618), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT62), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1353gat));
  INV_X1    g723(.A(G211gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n911), .A2(new_n925), .A3(new_n591), .ZN(new_n926));
  INV_X1    g725(.A(new_n909), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n591), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT63), .B(G211gat), .C1(new_n909), .C2(new_n697), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(G1354gat));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n646), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n909), .A2(KEYINPUT127), .ZN(new_n935));
  OAI21_X1  g734(.A(G218gat), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(G218gat), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n911), .A2(new_n937), .A3(new_n646), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1355gat));
endmodule


