

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n797), .A2(n746), .ZN(n514) );
  INV_X1 U553 ( .A(KEYINPUT30), .ZN(n680) );
  XNOR2_X1 U554 ( .A(n680), .B(KEYINPUT93), .ZN(n681) );
  XNOR2_X1 U555 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U556 ( .A1(n719), .A2(n718), .ZN(n733) );
  NAND2_X1 U557 ( .A1(n677), .A2(n753), .ZN(n723) );
  NAND2_X1 U558 ( .A1(G8), .A2(n723), .ZN(n797) );
  NOR2_X1 U559 ( .A1(G651), .A2(n616), .ZN(n634) );
  XNOR2_X1 U560 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n516) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XNOR2_X1 U562 ( .A(n516), .B(n515), .ZN(n593) );
  NAND2_X1 U563 ( .A1(G137), .A2(n593), .ZN(n518) );
  AND2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n877) );
  NAND2_X1 U565 ( .A1(G113), .A2(n877), .ZN(n517) );
  NAND2_X1 U566 ( .A1(n518), .A2(n517), .ZN(n520) );
  INV_X1 U567 ( .A(KEYINPUT68), .ZN(n519) );
  XNOR2_X1 U568 ( .A(n520), .B(n519), .ZN(n522) );
  INV_X1 U569 ( .A(G2105), .ZN(n523) );
  NOR2_X1 U570 ( .A1(G2104), .A2(n523), .ZN(n876) );
  NAND2_X1 U571 ( .A1(n876), .A2(G125), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n527) );
  AND2_X1 U573 ( .A1(G2104), .A2(n523), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n524), .B(KEYINPUT66), .ZN(n669) );
  NAND2_X1 U575 ( .A1(G101), .A2(n669), .ZN(n525) );
  XNOR2_X1 U576 ( .A(KEYINPUT23), .B(n525), .ZN(n526) );
  NOR2_X2 U577 ( .A1(n527), .A2(n526), .ZN(G160) );
  AND2_X1 U578 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U579 ( .A(G82), .ZN(G220) );
  INV_X1 U580 ( .A(G120), .ZN(G236) );
  INV_X1 U581 ( .A(G651), .ZN(n534) );
  XOR2_X1 U582 ( .A(G543), .B(KEYINPUT0), .Z(n528) );
  XNOR2_X1 U583 ( .A(KEYINPUT70), .B(n528), .ZN(n616) );
  NOR2_X1 U584 ( .A1(n534), .A2(n616), .ZN(n630) );
  NAND2_X1 U585 ( .A1(n630), .A2(G76), .ZN(n529) );
  XNOR2_X1 U586 ( .A(KEYINPUT78), .B(n529), .ZN(n532) );
  NOR2_X1 U587 ( .A1(G543), .A2(G651), .ZN(n633) );
  NAND2_X1 U588 ( .A1(n633), .A2(G89), .ZN(n530) );
  XNOR2_X1 U589 ( .A(KEYINPUT4), .B(n530), .ZN(n531) );
  NAND2_X1 U590 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U591 ( .A(n533), .B(KEYINPUT5), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G51), .A2(n634), .ZN(n538) );
  NOR2_X1 U593 ( .A1(G543), .A2(n534), .ZN(n535) );
  XOR2_X1 U594 ( .A(KEYINPUT72), .B(n535), .Z(n536) );
  XNOR2_X1 U595 ( .A(KEYINPUT1), .B(n536), .ZN(n639) );
  NAND2_X1 U596 ( .A1(G63), .A2(n639), .ZN(n537) );
  NAND2_X1 U597 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U598 ( .A(KEYINPUT6), .B(n539), .Z(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U600 ( .A(n542), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U601 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U602 ( .A1(G7), .A2(G661), .ZN(n543) );
  XNOR2_X1 U603 ( .A(n543), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U604 ( .A(G223), .ZN(n823) );
  NAND2_X1 U605 ( .A1(n823), .A2(G567), .ZN(n544) );
  XOR2_X1 U606 ( .A(KEYINPUT11), .B(n544), .Z(G234) );
  NAND2_X1 U607 ( .A1(n639), .A2(G56), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT14), .B(n545), .Z(n552) );
  NAND2_X1 U609 ( .A1(n630), .A2(G68), .ZN(n546) );
  XNOR2_X1 U610 ( .A(KEYINPUT75), .B(n546), .ZN(n549) );
  NAND2_X1 U611 ( .A1(n633), .A2(G81), .ZN(n547) );
  XOR2_X1 U612 ( .A(KEYINPUT12), .B(n547), .Z(n548) );
  NOR2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n550), .B(KEYINPUT13), .ZN(n551) );
  NOR2_X1 U615 ( .A1(n552), .A2(n551), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n634), .A2(G43), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n921) );
  INV_X1 U618 ( .A(G860), .ZN(n582) );
  OR2_X1 U619 ( .A1(n921), .A2(n582), .ZN(G153) );
  NAND2_X1 U620 ( .A1(G77), .A2(n630), .ZN(n556) );
  NAND2_X1 U621 ( .A1(G90), .A2(n633), .ZN(n555) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(KEYINPUT9), .B(n557), .ZN(n562) );
  NAND2_X1 U624 ( .A1(G52), .A2(n634), .ZN(n559) );
  NAND2_X1 U625 ( .A1(G64), .A2(n639), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT73), .B(n560), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(G301) );
  NAND2_X1 U629 ( .A1(G301), .A2(G868), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT76), .ZN(n572) );
  NAND2_X1 U631 ( .A1(G79), .A2(n630), .ZN(n565) );
  NAND2_X1 U632 ( .A1(G92), .A2(n633), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U634 ( .A1(G54), .A2(n634), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G66), .A2(n639), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U638 ( .A(KEYINPUT15), .B(n570), .Z(n916) );
  OR2_X1 U639 ( .A1(G868), .A2(n916), .ZN(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT77), .B(n573), .Z(G284) );
  NAND2_X1 U642 ( .A1(G78), .A2(n630), .ZN(n575) );
  NAND2_X1 U643 ( .A1(G91), .A2(n633), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G53), .A2(n634), .ZN(n577) );
  NAND2_X1 U646 ( .A1(G65), .A2(n639), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n924) );
  INV_X1 U649 ( .A(n924), .ZN(G299) );
  INV_X1 U650 ( .A(G868), .ZN(n642) );
  NOR2_X1 U651 ( .A1(G286), .A2(n642), .ZN(n581) );
  NOR2_X1 U652 ( .A1(G868), .A2(G299), .ZN(n580) );
  NOR2_X1 U653 ( .A1(n581), .A2(n580), .ZN(G297) );
  NAND2_X1 U654 ( .A1(n582), .A2(G559), .ZN(n583) );
  NAND2_X1 U655 ( .A1(n583), .A2(n916), .ZN(n584) );
  XNOR2_X1 U656 ( .A(n584), .B(KEYINPUT16), .ZN(n585) );
  XOR2_X1 U657 ( .A(KEYINPUT79), .B(n585), .Z(G148) );
  NAND2_X1 U658 ( .A1(n916), .A2(G868), .ZN(n586) );
  NOR2_X1 U659 ( .A1(G559), .A2(n586), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n587), .B(KEYINPUT80), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n921), .A2(G868), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G282) );
  NAND2_X1 U663 ( .A1(n876), .A2(G123), .ZN(n590) );
  XNOR2_X1 U664 ( .A(n590), .B(KEYINPUT18), .ZN(n592) );
  NAND2_X1 U665 ( .A1(G111), .A2(n877), .ZN(n591) );
  NAND2_X1 U666 ( .A1(n592), .A2(n591), .ZN(n597) );
  BUF_X1 U667 ( .A(n593), .Z(n882) );
  NAND2_X1 U668 ( .A1(G135), .A2(n882), .ZN(n595) );
  BUF_X1 U669 ( .A(n669), .Z(n880) );
  NAND2_X1 U670 ( .A1(G99), .A2(n880), .ZN(n594) );
  NAND2_X1 U671 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U672 ( .A1(n597), .A2(n596), .ZN(n976) );
  XNOR2_X1 U673 ( .A(G2096), .B(n976), .ZN(n599) );
  INV_X1 U674 ( .A(G2100), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(G156) );
  NAND2_X1 U676 ( .A1(G80), .A2(n630), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G93), .A2(n633), .ZN(n600) );
  NAND2_X1 U678 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U679 ( .A1(G55), .A2(n634), .ZN(n602) );
  XNOR2_X1 U680 ( .A(KEYINPUT81), .B(n602), .ZN(n603) );
  NOR2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U682 ( .A1(G67), .A2(n639), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n644) );
  NAND2_X1 U684 ( .A1(n916), .A2(G559), .ZN(n651) );
  XNOR2_X1 U685 ( .A(n921), .B(n651), .ZN(n607) );
  NOR2_X1 U686 ( .A1(G860), .A2(n607), .ZN(n608) );
  XOR2_X1 U687 ( .A(n644), .B(n608), .Z(G145) );
  NAND2_X1 U688 ( .A1(G75), .A2(n630), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G50), .A2(n634), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U691 ( .A1(G88), .A2(n633), .ZN(n611) );
  XNOR2_X1 U692 ( .A(KEYINPUT83), .B(n611), .ZN(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G62), .A2(n639), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G303) );
  INV_X1 U696 ( .A(G303), .ZN(G166) );
  NAND2_X1 U697 ( .A1(G49), .A2(n634), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G87), .A2(n616), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n639), .A2(n619), .ZN(n621) );
  NAND2_X1 U701 ( .A1(G651), .A2(G74), .ZN(n620) );
  NAND2_X1 U702 ( .A1(n621), .A2(n620), .ZN(G288) );
  NAND2_X1 U703 ( .A1(G47), .A2(n634), .ZN(n623) );
  NAND2_X1 U704 ( .A1(G60), .A2(n639), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G72), .A2(n630), .ZN(n624) );
  XNOR2_X1 U707 ( .A(KEYINPUT71), .B(n624), .ZN(n625) );
  NOR2_X1 U708 ( .A1(n626), .A2(n625), .ZN(n629) );
  NAND2_X1 U709 ( .A1(n633), .A2(G85), .ZN(n627) );
  XOR2_X1 U710 ( .A(KEYINPUT69), .B(n627), .Z(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(G290) );
  XOR2_X1 U712 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n632) );
  NAND2_X1 U713 ( .A1(G73), .A2(n630), .ZN(n631) );
  XNOR2_X1 U714 ( .A(n632), .B(n631), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G86), .A2(n633), .ZN(n636) );
  NAND2_X1 U716 ( .A1(G48), .A2(n634), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U719 ( .A1(G61), .A2(n639), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U721 ( .A1(n642), .A2(n644), .ZN(n643) );
  XNOR2_X1 U722 ( .A(n643), .B(KEYINPUT84), .ZN(n654) );
  XNOR2_X1 U723 ( .A(KEYINPUT19), .B(G288), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U725 ( .A(G166), .B(n646), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n921), .B(n924), .ZN(n647) );
  XNOR2_X1 U727 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n649), .B(G290), .ZN(n650) );
  XNOR2_X1 U729 ( .A(n650), .B(G305), .ZN(n895) );
  XOR2_X1 U730 ( .A(n895), .B(n651), .Z(n652) );
  NAND2_X1 U731 ( .A1(G868), .A2(n652), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2084), .A2(G2078), .ZN(n655) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U736 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XOR2_X1 U738 ( .A(KEYINPUT85), .B(G44), .Z(n659) );
  XNOR2_X1 U739 ( .A(KEYINPUT3), .B(n659), .ZN(G218) );
  XOR2_X1 U740 ( .A(KEYINPUT74), .B(G132), .Z(G219) );
  NAND2_X1 U741 ( .A1(G69), .A2(G108), .ZN(n660) );
  NOR2_X1 U742 ( .A1(G236), .A2(n660), .ZN(n661) );
  NAND2_X1 U743 ( .A1(G57), .A2(n661), .ZN(n827) );
  NAND2_X1 U744 ( .A1(n827), .A2(G567), .ZN(n667) );
  NOR2_X1 U745 ( .A1(G219), .A2(G220), .ZN(n662) );
  XNOR2_X1 U746 ( .A(KEYINPUT22), .B(n662), .ZN(n663) );
  NAND2_X1 U747 ( .A1(n663), .A2(G96), .ZN(n664) );
  NOR2_X1 U748 ( .A1(G218), .A2(n664), .ZN(n665) );
  XOR2_X1 U749 ( .A(KEYINPUT86), .B(n665), .Z(n828) );
  NAND2_X1 U750 ( .A1(G2106), .A2(n828), .ZN(n666) );
  NAND2_X1 U751 ( .A1(n667), .A2(n666), .ZN(n829) );
  NAND2_X1 U752 ( .A1(G661), .A2(G483), .ZN(n668) );
  NOR2_X1 U753 ( .A1(n829), .A2(n668), .ZN(n826) );
  NAND2_X1 U754 ( .A1(n826), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(G138), .A2(n882), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G102), .A2(n669), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G126), .A2(n876), .ZN(n673) );
  NAND2_X1 U759 ( .A1(G114), .A2(n877), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U761 ( .A1(n675), .A2(n674), .ZN(G164) );
  INV_X1 U762 ( .A(G301), .ZN(G171) );
  NAND2_X1 U763 ( .A1(G40), .A2(G160), .ZN(n676) );
  XOR2_X1 U764 ( .A(n676), .B(KEYINPUT87), .Z(n752) );
  INV_X1 U765 ( .A(n752), .ZN(n677) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n753) );
  NOR2_X1 U767 ( .A1(G1966), .A2(n797), .ZN(n732) );
  NOR2_X1 U768 ( .A1(G2084), .A2(n723), .ZN(n734) );
  NOR2_X1 U769 ( .A1(n732), .A2(n734), .ZN(n678) );
  XNOR2_X1 U770 ( .A(n678), .B(KEYINPUT92), .ZN(n679) );
  NAND2_X1 U771 ( .A1(n679), .A2(G8), .ZN(n682) );
  NOR2_X1 U772 ( .A1(G168), .A2(n683), .ZN(n687) );
  XNOR2_X1 U773 ( .A(G2078), .B(KEYINPUT25), .ZN(n951) );
  NOR2_X1 U774 ( .A1(n723), .A2(n951), .ZN(n685) );
  INV_X1 U775 ( .A(n723), .ZN(n690) );
  INV_X1 U776 ( .A(G1961), .ZN(n1000) );
  NOR2_X1 U777 ( .A1(n690), .A2(n1000), .ZN(n684) );
  NOR2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n715) );
  NOR2_X1 U779 ( .A1(G171), .A2(n715), .ZN(n686) );
  NOR2_X1 U780 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n688), .B(KEYINPUT94), .ZN(n689) );
  XNOR2_X1 U782 ( .A(n689), .B(KEYINPUT31), .ZN(n719) );
  NAND2_X1 U783 ( .A1(n690), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U784 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  AND2_X1 U785 ( .A1(G1956), .A2(n723), .ZN(n692) );
  NOR2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n695) );
  NOR2_X1 U787 ( .A1(n695), .A2(n924), .ZN(n694) );
  XOR2_X1 U788 ( .A(n694), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U789 ( .A1(n695), .A2(n924), .ZN(n711) );
  INV_X1 U790 ( .A(G1996), .ZN(n948) );
  NOR2_X1 U791 ( .A1(n723), .A2(n948), .ZN(n697) );
  XOR2_X1 U792 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n696) );
  XNOR2_X1 U793 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n723), .A2(G1341), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U796 ( .A(KEYINPUT91), .B(n700), .Z(n701) );
  NOR2_X1 U797 ( .A1(n921), .A2(n701), .ZN(n702) );
  XNOR2_X1 U798 ( .A(KEYINPUT65), .B(n702), .ZN(n706) );
  AND2_X1 U799 ( .A1(n723), .A2(G1348), .ZN(n704) );
  INV_X1 U800 ( .A(G2067), .ZN(n943) );
  NOR2_X1 U801 ( .A1(n723), .A2(n943), .ZN(n703) );
  NOR2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n916), .A2(n707), .ZN(n705) );
  NAND2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n709) );
  OR2_X1 U805 ( .A1(n916), .A2(n707), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U809 ( .A(n714), .B(KEYINPUT29), .ZN(n717) );
  AND2_X1 U810 ( .A1(G171), .A2(n715), .ZN(n716) );
  NOR2_X1 U811 ( .A1(n717), .A2(n716), .ZN(n718) );
  INV_X1 U812 ( .A(n733), .ZN(n721) );
  AND2_X1 U813 ( .A1(G286), .A2(G8), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n730) );
  INV_X1 U815 ( .A(G8), .ZN(n728) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n797), .ZN(n722) );
  XNOR2_X1 U817 ( .A(n722), .B(KEYINPUT96), .ZN(n725) );
  NOR2_X1 U818 ( .A1(n723), .A2(G2090), .ZN(n724) );
  NOR2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U820 ( .A1(n726), .A2(G303), .ZN(n727) );
  OR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  AND2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n731), .B(KEYINPUT32), .ZN(n740) );
  INV_X1 U824 ( .A(KEYINPUT95), .ZN(n738) );
  NOR2_X1 U825 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U826 ( .A1(G8), .A2(n734), .ZN(n735) );
  NAND2_X1 U827 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U828 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n796) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n741) );
  XNOR2_X1 U831 ( .A(n741), .B(KEYINPUT97), .ZN(n742) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n750) );
  INV_X1 U833 ( .A(n750), .ZN(n928) );
  AND2_X1 U834 ( .A1(n742), .A2(n928), .ZN(n744) );
  INV_X1 U835 ( .A(KEYINPUT33), .ZN(n743) );
  AND2_X1 U836 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U837 ( .A1(n796), .A2(n745), .ZN(n748) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n927) );
  INV_X1 U839 ( .A(n927), .ZN(n746) );
  OR2_X1 U840 ( .A1(KEYINPUT33), .A2(n514), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n749), .B(KEYINPUT98), .ZN(n788) );
  NAND2_X1 U843 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  OR2_X1 U844 ( .A1(n797), .A2(n751), .ZN(n786) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n934) );
  XNOR2_X1 U846 ( .A(G1986), .B(G290), .ZN(n918) );
  NOR2_X1 U847 ( .A1(n753), .A2(n752), .ZN(n816) );
  AND2_X1 U848 ( .A1(n918), .A2(n816), .ZN(n783) );
  NAND2_X1 U849 ( .A1(G131), .A2(n882), .ZN(n755) );
  NAND2_X1 U850 ( .A1(G95), .A2(n880), .ZN(n754) );
  NAND2_X1 U851 ( .A1(n755), .A2(n754), .ZN(n759) );
  NAND2_X1 U852 ( .A1(G119), .A2(n876), .ZN(n757) );
  NAND2_X1 U853 ( .A1(G107), .A2(n877), .ZN(n756) );
  NAND2_X1 U854 ( .A1(n757), .A2(n756), .ZN(n758) );
  NOR2_X1 U855 ( .A1(n759), .A2(n758), .ZN(n873) );
  INV_X1 U856 ( .A(G1991), .ZN(n949) );
  NOR2_X1 U857 ( .A1(n873), .A2(n949), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G129), .A2(n876), .ZN(n761) );
  NAND2_X1 U859 ( .A1(G117), .A2(n877), .ZN(n760) );
  NAND2_X1 U860 ( .A1(n761), .A2(n760), .ZN(n764) );
  NAND2_X1 U861 ( .A1(G105), .A2(n880), .ZN(n762) );
  XOR2_X1 U862 ( .A(KEYINPUT38), .B(n762), .Z(n763) );
  NOR2_X1 U863 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U864 ( .A(n765), .B(KEYINPUT90), .ZN(n767) );
  NAND2_X1 U865 ( .A1(G141), .A2(n882), .ZN(n766) );
  NAND2_X1 U866 ( .A1(n767), .A2(n766), .ZN(n888) );
  AND2_X1 U867 ( .A1(n888), .A2(G1996), .ZN(n768) );
  NOR2_X1 U868 ( .A1(n769), .A2(n768), .ZN(n978) );
  INV_X1 U869 ( .A(n978), .ZN(n770) );
  NAND2_X1 U870 ( .A1(n770), .A2(n816), .ZN(n803) );
  NAND2_X1 U871 ( .A1(G140), .A2(n882), .ZN(n772) );
  NAND2_X1 U872 ( .A1(G104), .A2(n880), .ZN(n771) );
  NAND2_X1 U873 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U874 ( .A(KEYINPUT34), .B(n773), .ZN(n780) );
  NAND2_X1 U875 ( .A1(n877), .A2(G116), .ZN(n774) );
  XNOR2_X1 U876 ( .A(KEYINPUT89), .B(n774), .ZN(n777) );
  NAND2_X1 U877 ( .A1(n876), .A2(G128), .ZN(n775) );
  XOR2_X1 U878 ( .A(KEYINPUT88), .B(n775), .Z(n776) );
  NOR2_X1 U879 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U880 ( .A(n778), .B(KEYINPUT35), .ZN(n779) );
  NOR2_X1 U881 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U882 ( .A(KEYINPUT36), .B(n781), .ZN(n891) );
  XNOR2_X1 U883 ( .A(KEYINPUT37), .B(G2067), .ZN(n814) );
  NOR2_X1 U884 ( .A1(n891), .A2(n814), .ZN(n973) );
  NAND2_X1 U885 ( .A1(n816), .A2(n973), .ZN(n811) );
  NAND2_X1 U886 ( .A1(n803), .A2(n811), .ZN(n782) );
  OR2_X1 U887 ( .A1(n783), .A2(n782), .ZN(n802) );
  INV_X1 U888 ( .A(n802), .ZN(n784) );
  AND2_X1 U889 ( .A1(n934), .A2(n784), .ZN(n785) );
  NAND2_X1 U890 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U891 ( .A1(n788), .A2(n787), .ZN(n821) );
  NOR2_X1 U892 ( .A1(G2090), .A2(G303), .ZN(n789) );
  XOR2_X1 U893 ( .A(KEYINPUT99), .B(n789), .Z(n790) );
  NAND2_X1 U894 ( .A1(n790), .A2(G8), .ZN(n794) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XOR2_X1 U896 ( .A(n791), .B(KEYINPUT24), .Z(n792) );
  NOR2_X1 U897 ( .A1(n797), .A2(n792), .ZN(n798) );
  INV_X1 U898 ( .A(n798), .ZN(n793) );
  AND2_X1 U899 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U900 ( .A1(n796), .A2(n795), .ZN(n800) );
  OR2_X1 U901 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U902 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U903 ( .A1(n802), .A2(n801), .ZN(n819) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n888), .ZN(n988) );
  INV_X1 U905 ( .A(n803), .ZN(n807) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n805) );
  AND2_X1 U907 ( .A1(n949), .A2(n873), .ZN(n804) );
  XNOR2_X1 U908 ( .A(KEYINPUT100), .B(n804), .ZN(n980) );
  NOR2_X1 U909 ( .A1(n805), .A2(n980), .ZN(n806) );
  NOR2_X1 U910 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U911 ( .A1(n988), .A2(n808), .ZN(n809) );
  XOR2_X1 U912 ( .A(KEYINPUT39), .B(n809), .Z(n810) );
  XNOR2_X1 U913 ( .A(KEYINPUT101), .B(n810), .ZN(n812) );
  NAND2_X1 U914 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U915 ( .A(n813), .B(KEYINPUT102), .ZN(n815) );
  NAND2_X1 U916 ( .A1(n891), .A2(n814), .ZN(n972) );
  NAND2_X1 U917 ( .A1(n815), .A2(n972), .ZN(n817) );
  NAND2_X1 U918 ( .A1(n817), .A2(n816), .ZN(n818) );
  AND2_X1 U919 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U920 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U921 ( .A(n822), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U924 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U926 ( .A1(n826), .A2(n825), .ZN(G188) );
  XOR2_X1 U927 ( .A(G96), .B(KEYINPUT104), .Z(G221) );
  XNOR2_X1 U928 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  XOR2_X1 U929 ( .A(G108), .B(KEYINPUT116), .Z(G238) );
  NOR2_X1 U931 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  INV_X1 U933 ( .A(n829), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT108), .B(G1981), .Z(n831) );
  XNOR2_X1 U935 ( .A(G1961), .B(G1956), .ZN(n830) );
  XNOR2_X1 U936 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U937 ( .A(n832), .B(KEYINPUT41), .Z(n834) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n833) );
  XNOR2_X1 U939 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n836) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1966), .ZN(n835) );
  XNOR2_X1 U942 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U943 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U944 ( .A(KEYINPUT107), .B(G2474), .ZN(n839) );
  XNOR2_X1 U945 ( .A(n840), .B(n839), .ZN(G229) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U947 ( .A(G2090), .B(G2678), .ZN(n841) );
  XNOR2_X1 U948 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U949 ( .A(n843), .B(KEYINPUT106), .Z(n845) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U951 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U952 ( .A(KEYINPUT42), .B(G2100), .Z(n847) );
  XNOR2_X1 U953 ( .A(G2084), .B(G2078), .ZN(n846) );
  XNOR2_X1 U954 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U955 ( .A(n849), .B(n848), .ZN(G227) );
  NAND2_X1 U956 ( .A1(n876), .A2(G124), .ZN(n850) );
  XNOR2_X1 U957 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U958 ( .A1(G112), .A2(n877), .ZN(n851) );
  NAND2_X1 U959 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U960 ( .A1(G136), .A2(n882), .ZN(n854) );
  NAND2_X1 U961 ( .A1(G100), .A2(n880), .ZN(n853) );
  NAND2_X1 U962 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U963 ( .A1(n856), .A2(n855), .ZN(G162) );
  XOR2_X1 U964 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n858) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n857) );
  XNOR2_X1 U966 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U967 ( .A(n859), .B(G162), .Z(n871) );
  NAND2_X1 U968 ( .A1(n880), .A2(G103), .ZN(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT111), .B(KEYINPUT47), .ZN(n863) );
  NAND2_X1 U970 ( .A1(G127), .A2(n876), .ZN(n861) );
  NAND2_X1 U971 ( .A1(G115), .A2(n877), .ZN(n860) );
  NAND2_X1 U972 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U973 ( .A(n863), .B(n862), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n882), .A2(G139), .ZN(n864) );
  XOR2_X1 U975 ( .A(KEYINPUT110), .B(n864), .Z(n865) );
  NOR2_X1 U976 ( .A1(n866), .A2(n865), .ZN(n867) );
  NAND2_X1 U977 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U978 ( .A(n869), .B(KEYINPUT112), .ZN(n983) );
  XNOR2_X1 U979 ( .A(G164), .B(n983), .ZN(n870) );
  XNOR2_X1 U980 ( .A(n871), .B(n870), .ZN(n872) );
  XOR2_X1 U981 ( .A(n872), .B(n976), .Z(n875) );
  XNOR2_X1 U982 ( .A(G160), .B(n873), .ZN(n874) );
  XNOR2_X1 U983 ( .A(n875), .B(n874), .ZN(n893) );
  NAND2_X1 U984 ( .A1(G130), .A2(n876), .ZN(n879) );
  NAND2_X1 U985 ( .A1(G118), .A2(n877), .ZN(n878) );
  NAND2_X1 U986 ( .A1(n879), .A2(n878), .ZN(n887) );
  NAND2_X1 U987 ( .A1(G106), .A2(n880), .ZN(n881) );
  XOR2_X1 U988 ( .A(KEYINPUT109), .B(n881), .Z(n884) );
  NAND2_X1 U989 ( .A1(n882), .A2(G142), .ZN(n883) );
  NAND2_X1 U990 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U991 ( .A(n885), .B(KEYINPUT45), .Z(n886) );
  NOR2_X1 U992 ( .A1(n887), .A2(n886), .ZN(n889) );
  XNOR2_X1 U993 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U994 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U996 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U997 ( .A(n916), .B(G286), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U999 ( .A(G301), .B(n897), .Z(n898) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n898), .ZN(n899) );
  XOR2_X1 U1001 ( .A(KEYINPUT115), .B(n899), .Z(G397) );
  XOR2_X1 U1002 ( .A(G2454), .B(G2430), .Z(n901) );
  XNOR2_X1 U1003 ( .A(G2451), .B(G2446), .ZN(n900) );
  XNOR2_X1 U1004 ( .A(n901), .B(n900), .ZN(n908) );
  XOR2_X1 U1005 ( .A(G2443), .B(G2427), .Z(n903) );
  XNOR2_X1 U1006 ( .A(G2438), .B(KEYINPUT103), .ZN(n902) );
  XNOR2_X1 U1007 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1008 ( .A(n904), .B(G2435), .Z(n906) );
  XNOR2_X1 U1009 ( .A(G1348), .B(G1341), .ZN(n905) );
  XNOR2_X1 U1010 ( .A(n906), .B(n905), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(n908), .B(n907), .ZN(n909) );
  NAND2_X1 U1012 ( .A1(n909), .A2(G14), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1016 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1018 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  INV_X1 U1021 ( .A(n915), .ZN(G401) );
  XNOR2_X1 U1022 ( .A(n916), .B(G1348), .ZN(n920) );
  XNOR2_X1 U1023 ( .A(G1961), .B(G301), .ZN(n917) );
  NOR2_X1 U1024 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1025 ( .A1(n920), .A2(n919), .ZN(n923) );
  XNOR2_X1 U1026 ( .A(G1341), .B(n921), .ZN(n922) );
  NOR2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(G166), .B(G1971), .ZN(n926) );
  XNOR2_X1 U1029 ( .A(n924), .B(G1956), .ZN(n925) );
  NAND2_X1 U1030 ( .A1(n926), .A2(n925), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1033 ( .A(KEYINPUT123), .B(n931), .Z(n932) );
  NAND2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(G1966), .B(G168), .ZN(n935) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(n936), .B(KEYINPUT57), .ZN(n937) );
  XOR2_X1 U1038 ( .A(KEYINPUT122), .B(n937), .Z(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G16), .B(KEYINPUT56), .ZN(n940) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n971) );
  XNOR2_X1 U1043 ( .A(n943), .B(G26), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G2072), .B(G33), .ZN(n944) );
  XNOR2_X1 U1045 ( .A(n944), .B(KEYINPUT117), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n947), .B(KEYINPUT118), .ZN(n957) );
  XNOR2_X1 U1048 ( .A(G32), .B(n948), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G25), .B(n949), .ZN(n950) );
  NAND2_X1 U1050 ( .A1(n950), .A2(G28), .ZN(n953) );
  XOR2_X1 U1051 ( .A(G27), .B(n951), .Z(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT53), .B(n958), .Z(n962) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(G34), .ZN(n959) );
  XNOR2_X1 U1057 ( .A(n959), .B(KEYINPUT119), .ZN(n960) );
  XNOR2_X1 U1058 ( .A(G2084), .B(n960), .ZN(n961) );
  NAND2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(G35), .B(G2090), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(KEYINPUT55), .B(n965), .ZN(n967) );
  INV_X1 U1063 ( .A(G29), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n968), .A2(G11), .ZN(n969) );
  XNOR2_X1 U1066 ( .A(KEYINPUT120), .B(n969), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n999) );
  INV_X1 U1068 ( .A(n972), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n982) );
  XOR2_X1 U1070 ( .A(G2084), .B(G160), .Z(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n993) );
  XOR2_X1 U1075 ( .A(G164), .B(G2078), .Z(n985) );
  XNOR2_X1 U1076 ( .A(G2072), .B(n983), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT50), .B(n986), .ZN(n991) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n987) );
  NOR2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n989), .Z(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(KEYINPUT52), .B(n994), .ZN(n996) );
  INV_X1 U1085 ( .A(KEYINPUT55), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(G29), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1027) );
  XNOR2_X1 U1089 ( .A(n1000), .B(G5), .ZN(n1021) );
  XOR2_X1 U1090 ( .A(G1966), .B(G21), .Z(n1011) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(G4), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1956), .B(G20), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(KEYINPUT125), .B(G1341), .Z(n1006) );
  XNOR2_X1 U1098 ( .A(G19), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1009), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  XNOR2_X1 U1102 ( .A(G1986), .B(G24), .ZN(n1013) );
  XNOR2_X1 U1103 ( .A(G1971), .B(G22), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(G1976), .B(KEYINPUT126), .Z(n1014) );
  XNOR2_X1 U1106 ( .A(G23), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(n1022), .B(KEYINPUT61), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1023), .Z(n1025) );
  XNOR2_X1 U1113 ( .A(KEYINPUT124), .B(G16), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(n1028), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

