//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1211, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G13), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  NAND2_X1  g0009(.A1(G107), .A2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G50), .B2(G226), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G97), .A2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G116), .ZN(new_n219));
  INV_X1    g0019(.A(G270), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n218), .A2(new_n221), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G77), .A2(G244), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n204), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n216), .A2(new_n211), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n209), .B(new_n228), .C1(new_n231), .C2(new_n234), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G264), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n220), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(KEYINPUT66), .B(G107), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(G116), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  XNOR2_X1  g0052(.A(KEYINPUT3), .B(G33), .ZN(new_n253));
  INV_X1    g0053(.A(G1698), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G222), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  OAI211_X1 g0056(.A(new_n253), .B(new_n255), .C1(new_n256), .C2(new_n254), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n229), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n257), .B(new_n259), .C1(G77), .C2(new_n253), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n261), .A2(G1), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT67), .A2(G41), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT67), .A2(G41), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR3_X1   g0066(.A1(new_n258), .A2(KEYINPUT68), .A3(new_n229), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT68), .ZN(new_n268));
  AND2_X1   g0068(.A1(G1), .A2(G13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G41), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n262), .B(new_n266), .C1(new_n267), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G226), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1), .B1(new_n274), .B2(new_n263), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT68), .B1(new_n258), .B2(new_n229), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n269), .A2(new_n268), .A3(new_n270), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n260), .B(new_n272), .C1(new_n273), .C2(new_n279), .ZN(new_n280));
  OR2_X1    g0080(.A1(new_n280), .A2(G179), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT69), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT69), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n284), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n283), .A2(new_n229), .A3(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(G20), .B1(new_n232), .B2(G50), .ZN(new_n287));
  INV_X1    g0087(.A(G150), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n230), .A2(G33), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT8), .B(G58), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n287), .B1(new_n288), .B2(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G1), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n286), .B1(new_n294), .B2(G20), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n286), .A2(new_n293), .B1(new_n295), .B2(G50), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(G13), .A3(G20), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n296), .B1(G50), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G169), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n280), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n281), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n298), .B1(KEYINPUT72), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n304));
  XOR2_X1   g0104(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n280), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(G200), .B2(new_n280), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n301), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G33), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT3), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT7), .B1(new_n317), .B2(new_n230), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  AOI211_X1 g0119(.A(new_n319), .B(G20), .C1(new_n314), .C2(new_n316), .ZN(new_n320));
  OAI21_X1  g0120(.A(G68), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n289), .A2(G159), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G58), .A2(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n232), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G20), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n321), .A2(KEYINPUT16), .A3(new_n322), .A4(new_n325), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n328), .A2(new_n286), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n256), .A2(new_n254), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n273), .A2(G1698), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n314), .A2(new_n331), .A3(new_n316), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(G33), .A2(G87), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n259), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n276), .A2(new_n277), .ZN(new_n337));
  INV_X1    g0137(.A(new_n275), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G232), .A3(new_n338), .ZN(new_n339));
  AND3_X1   g0139(.A1(new_n336), .A2(new_n272), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G190), .ZN(new_n341));
  INV_X1    g0141(.A(new_n297), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n292), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n292), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n295), .A2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n330), .A2(new_n341), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT17), .B1(new_n349), .B2(KEYINPUT75), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT17), .ZN(new_n352));
  NOR4_X1   g0152(.A1(new_n346), .A2(new_n351), .A3(new_n352), .A4(new_n348), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G50), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n290), .A2(new_n355), .B1(new_n230), .B2(G68), .ZN(new_n356));
  INV_X1    g0156(.A(G77), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n291), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n286), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT11), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n283), .A2(new_n285), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n229), .C1(G1), .C2(new_n230), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n360), .B1(new_n211), .B2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n294), .A2(new_n211), .A3(G13), .A4(G20), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT73), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT12), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n365), .ZN(new_n367));
  XOR2_X1   g0167(.A(new_n366), .B(new_n367), .Z(new_n368));
  NOR2_X1   g0168(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n217), .A2(G1698), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n370), .B1(G226), .B2(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G97), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n371), .A2(new_n317), .B1(new_n313), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n259), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n278), .A2(G238), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n375), .A3(new_n272), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT13), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(KEYINPUT13), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n369), .B1(new_n379), .B2(new_n306), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n347), .B1(new_n377), .B2(new_n378), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(G169), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n377), .A2(G179), .A3(new_n378), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT14), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n379), .A2(new_n386), .A3(G169), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n369), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n330), .A2(new_n343), .A3(new_n345), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT67), .B(G41), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n276), .A2(new_n277), .B1(new_n392), .B2(new_n263), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n262), .A2(new_n393), .B1(new_n278), .B2(G232), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n299), .B1(new_n394), .B2(new_n336), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n336), .A2(new_n339), .A3(G179), .A4(new_n272), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT74), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT74), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n399), .B(new_n396), .C1(new_n340), .C2(new_n299), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n391), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n391), .A2(new_n401), .A3(KEYINPUT18), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n354), .A2(new_n390), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n297), .A2(G77), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n362), .A2(new_n357), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n292), .A2(new_n290), .B1(new_n230), .B2(new_n357), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT70), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g0212(.A(KEYINPUT15), .B(G87), .Z(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n230), .A3(G33), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n408), .B(new_n409), .C1(new_n416), .C2(new_n286), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G238), .A2(G1698), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n253), .B(new_n418), .C1(new_n217), .C2(G1698), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n419), .B(new_n259), .C1(G107), .C2(new_n253), .ZN(new_n420));
  INV_X1    g0220(.A(G244), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n272), .C1(new_n421), .C2(new_n279), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n299), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(KEYINPUT71), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n409), .B1(new_n416), .B2(new_n286), .ZN(new_n426));
  INV_X1    g0226(.A(new_n408), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT71), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n422), .A2(G179), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n422), .A2(G200), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n306), .B2(new_n422), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n312), .A2(new_n407), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n254), .A2(G257), .ZN(new_n437));
  NAND2_X1  g0237(.A1(G264), .A2(G1698), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n253), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G303), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n317), .A2(new_n440), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n439), .A2(new_n259), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n264), .A2(new_n265), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT5), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n263), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT78), .B(KEYINPUT5), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT79), .B1(new_n446), .B2(G41), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n444), .A2(KEYINPUT78), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT78), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT79), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n451), .A2(new_n452), .A3(new_n274), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n445), .A2(new_n447), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n272), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n442), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n447), .A2(new_n453), .ZN(new_n457));
  OAI211_X1 g0257(.A(new_n294), .B(G45), .C1(new_n392), .C2(KEYINPUT5), .ZN(new_n458));
  OAI211_X1 g0258(.A(G270), .B(new_n337), .C1(new_n457), .C2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n299), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(G20), .B1(G33), .B2(G283), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(G33), .B2(new_n372), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n219), .A2(G20), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n286), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT20), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n286), .A2(KEYINPUT20), .A3(new_n462), .A4(new_n463), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n463), .A2(G1), .A3(new_n205), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n294), .A2(G33), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n297), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n286), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n472), .B2(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT21), .B1(new_n460), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n452), .B1(new_n451), .B2(new_n274), .ZN(new_n476));
  AOI211_X1 g0276(.A(KEYINPUT79), .B(G41), .C1(new_n448), .C2(new_n450), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n455), .A2(new_n478), .A3(new_n445), .ZN(new_n479));
  INV_X1    g0279(.A(new_n442), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n459), .A3(new_n480), .ZN(new_n481));
  AND4_X1   g0281(.A1(KEYINPUT21), .A2(new_n481), .A3(G169), .A4(new_n474), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n475), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT82), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n474), .A2(new_n456), .A3(G179), .A4(new_n459), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n481), .A2(G200), .ZN(new_n486));
  INV_X1    g0286(.A(new_n474), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n456), .A2(G190), .A3(new_n459), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n483), .A2(new_n484), .A3(new_n485), .A4(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n481), .A2(G169), .A3(new_n474), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT21), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n460), .A2(KEYINPUT21), .A3(new_n474), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n489), .A2(new_n493), .A3(new_n485), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(KEYINPUT82), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n314), .A2(new_n316), .A3(new_n230), .A4(G87), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n499));
  NAND2_X1  g0299(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n253), .A2(new_n230), .A3(G87), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n230), .A2(G107), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT23), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT84), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT24), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n502), .A2(KEYINPUT24), .A3(new_n504), .A4(new_n507), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n286), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n471), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n361), .A2(new_n513), .A3(G107), .A4(new_n229), .ZN(new_n514));
  AND2_X1   g0314(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(new_n297), .B2(G107), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT85), .A2(KEYINPUT25), .ZN(new_n517));
  OR4_X1    g0317(.A1(G107), .A2(new_n297), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n514), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT86), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n514), .A2(KEYINPUT86), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(G264), .B(new_n337), .C1(new_n457), .C2(new_n458), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n253), .B1(G257), .B2(new_n254), .ZN(new_n526));
  NOR2_X1   g0326(.A1(G250), .A2(G1698), .ZN(new_n527));
  INV_X1    g0327(.A(G294), .ZN(new_n528));
  OAI22_X1  g0328(.A1(new_n526), .A2(new_n527), .B1(new_n313), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n259), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n479), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n299), .ZN(new_n532));
  INV_X1    g0332(.A(G179), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n479), .A2(new_n525), .A3(new_n533), .A4(new_n530), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n524), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n531), .A2(G200), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n479), .A2(new_n525), .A3(G190), .A4(new_n530), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n512), .A3(new_n537), .A4(new_n523), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n223), .B1(new_n263), .B2(G1), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n263), .A2(G1), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n261), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n337), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n212), .A2(new_n254), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n421), .A2(G1698), .ZN(new_n544));
  AND2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n545), .A2(new_n253), .B1(G33), .B2(G116), .ZN(new_n546));
  INV_X1    g0346(.A(new_n259), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n548), .A2(new_n306), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n230), .ZN(new_n552));
  INV_X1    g0352(.A(G107), .ZN(new_n553));
  AND4_X1   g0353(.A1(KEYINPUT81), .A2(new_n222), .A3(new_n372), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(G87), .A2(G97), .ZN(new_n555));
  AOI21_X1  g0355(.A(KEYINPUT81), .B1(new_n555), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT19), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n291), .B2(new_n372), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n253), .A2(new_n230), .A3(G68), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n413), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n286), .B1(new_n342), .B2(new_n562), .ZN(new_n563));
  AND3_X1   g0363(.A1(new_n337), .A2(new_n539), .A3(new_n541), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n253), .A2(new_n543), .A3(new_n544), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n547), .B1(new_n565), .B2(new_n505), .ZN(new_n566));
  OAI21_X1  g0366(.A(G200), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n472), .A2(G87), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n472), .A2(new_n413), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n563), .A2(new_n570), .B1(new_n548), .B2(new_n299), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n564), .A2(new_n566), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n533), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n550), .A2(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n535), .A2(new_n538), .A3(new_n574), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n314), .A2(new_n316), .A3(G244), .A4(new_n254), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(KEYINPUT77), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n253), .A2(G244), .A3(new_n579), .A4(new_n254), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n582));
  INV_X1    g0382(.A(G283), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n582), .B1(new_n313), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n259), .B1(new_n581), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(G257), .B(new_n337), .C1(new_n457), .C2(new_n458), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n479), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n319), .B1(new_n253), .B2(G20), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n317), .A2(KEYINPUT7), .A3(new_n230), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n553), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g0392(.A(G97), .B(G107), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n594), .A2(new_n372), .A3(G107), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n598), .A2(G20), .B1(G77), .B2(new_n289), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n592), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(G97), .B1(new_n286), .B2(new_n471), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n297), .A2(new_n372), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT76), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT76), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n601), .A2(new_n605), .A3(new_n602), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n600), .A2(new_n286), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n585), .A2(new_n479), .A3(new_n586), .A4(G190), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n588), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n587), .A2(new_n299), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n604), .A2(new_n606), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n596), .B1(new_n594), .B2(new_n593), .ZN(new_n612));
  OAI22_X1  g0412(.A1(new_n612), .A2(new_n230), .B1(new_n357), .B2(new_n290), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n286), .B1(new_n613), .B2(new_n591), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n585), .A2(new_n479), .A3(new_n586), .A4(new_n533), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n610), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n609), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT80), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n609), .A2(new_n617), .A3(KEYINPUT80), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n575), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n436), .A2(new_n497), .A3(new_n622), .ZN(G372));
  NAND3_X1  g0423(.A1(new_n493), .A2(new_n485), .A3(new_n494), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT89), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT89), .A4(new_n485), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n535), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n609), .A2(new_n617), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT88), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n549), .B1(new_n632), .B2(KEYINPUT88), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n548), .A2(new_n299), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT87), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n636), .A2(new_n637), .B1(new_n563), .B2(new_n570), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n635), .A2(KEYINPUT87), .B1(new_n572), .B2(new_n533), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n633), .A2(new_n634), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n631), .A2(new_n538), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n629), .A2(new_n630), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT91), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n617), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n617), .A2(new_n645), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n640), .B(new_n644), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n574), .ZN(new_n649));
  OAI21_X1  g0449(.A(KEYINPUT26), .B1(new_n649), .B2(new_n617), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n638), .A2(new_n639), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n648), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n535), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n653), .B1(new_n626), .B2(new_n627), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT90), .B1(new_n654), .B2(new_n641), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n643), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n436), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n301), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n395), .A2(new_n397), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n391), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n403), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n391), .A2(new_n660), .A3(KEYINPUT18), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT92), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n432), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n425), .A2(new_n430), .A3(KEYINPUT92), .A4(new_n431), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n382), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n668), .B1(new_n389), .B2(new_n388), .ZN(new_n669));
  INV_X1    g0469(.A(new_n354), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n309), .B(KEYINPUT10), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n658), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n657), .A2(new_n673), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n294), .A2(new_n230), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n474), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n497), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n628), .B2(new_n681), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n524), .A2(new_n680), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n653), .B1(new_n538), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n535), .A2(new_n680), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(G330), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT93), .ZN(new_n689));
  INV_X1    g0489(.A(new_n686), .ZN(new_n690));
  INV_X1    g0490(.A(new_n680), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n687), .A2(new_n624), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n690), .A3(new_n692), .ZN(G399));
  NOR2_X1   g0493(.A1(new_n206), .A2(new_n443), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  OR3_X1    g0496(.A1(new_n554), .A2(new_n556), .A3(G116), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n696), .A2(new_n697), .B1(new_n233), .B2(new_n695), .ZN(new_n698));
  XOR2_X1   g0498(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n699));
  XNOR2_X1  g0499(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n656), .A2(new_n691), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n653), .A2(new_n624), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n641), .A2(new_n704), .ZN(new_n705));
  NOR3_X1   g0505(.A1(new_n649), .A2(KEYINPUT26), .A3(new_n617), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n706), .B1(new_n638), .B2(new_n639), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT26), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(KEYINPUT29), .A3(new_n691), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n497), .A2(new_n622), .A3(new_n691), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT96), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n587), .A2(new_n481), .A3(new_n533), .A4(new_n548), .ZN(new_n717));
  INV_X1    g0517(.A(new_n531), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n525), .A2(new_n530), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n587), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n481), .A2(new_n533), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n572), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n587), .A2(new_n720), .A3(new_n548), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n722), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n719), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n680), .B1(new_n728), .B2(KEYINPUT95), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT95), .ZN(new_n730));
  AOI211_X1 g0530(.A(new_n730), .B(new_n719), .C1(new_n724), .C2(new_n727), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n716), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n497), .A2(new_n622), .A3(KEYINPUT96), .A4(new_n691), .ZN(new_n733));
  INV_X1    g0533(.A(new_n727), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n726), .B1(new_n725), .B2(new_n722), .ZN(new_n735));
  OAI22_X1  g0535(.A1(new_n734), .A2(new_n735), .B1(new_n718), .B2(new_n717), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n715), .A2(new_n732), .A3(new_n733), .A4(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n712), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n700), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n683), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(G20), .B1(KEYINPUT99), .B2(G169), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(KEYINPUT99), .A2(G169), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n229), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n533), .A2(new_n347), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n230), .A2(G190), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n211), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n347), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n553), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G159), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT32), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n230), .A2(new_n306), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n751), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n755), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n764), .A2(new_n355), .B1(new_n765), .B2(new_n222), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n230), .B1(new_n758), .B2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n533), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n752), .A2(new_n768), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n253), .B1(new_n767), .B2(new_n372), .C1(new_n357), .C2(new_n769), .ZN(new_n770));
  OR4_X1    g0570(.A1(new_n757), .A2(new_n762), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n763), .A2(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n754), .B(new_n771), .C1(G58), .C2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n753), .ZN(new_n775));
  INV_X1    g0575(.A(G317), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(KEYINPUT33), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n760), .A2(G329), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n583), .C2(new_n756), .ZN(new_n781));
  INV_X1    g0581(.A(new_n764), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n781), .B1(G326), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n765), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(G303), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n253), .B1(new_n773), .B2(G322), .ZN(new_n786));
  INV_X1    g0586(.A(new_n767), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G294), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n783), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n769), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G311), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n750), .B1(new_n774), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(G355), .B(KEYINPUT98), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n207), .A2(new_n253), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n206), .A2(new_n253), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(G45), .B2(new_n233), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n251), .A2(G45), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n794), .B1(G116), .B2(new_n207), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n750), .A2(new_n744), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n230), .A2(G13), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT97), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n294), .B1(new_n802), .B2(G45), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n804), .A2(new_n694), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n746), .A2(new_n792), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n683), .A2(G330), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n683), .A2(G330), .ZN(new_n808));
  INV_X1    g0608(.A(new_n805), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n806), .B1(new_n807), .B2(new_n810), .ZN(G396));
  OAI21_X1  g0611(.A(new_n435), .B1(new_n417), .B2(new_n691), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n666), .A2(new_n428), .A3(new_n667), .A4(new_n680), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n701), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n814), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n656), .A2(new_n691), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(new_n739), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n809), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n814), .A2(new_n742), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n750), .A2(new_n742), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(new_n357), .ZN(new_n823));
  INV_X1    g0623(.A(G311), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n756), .A2(new_n222), .B1(new_n759), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT100), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n253), .B(new_n826), .C1(G294), .C2(new_n773), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n784), .A2(G107), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n775), .A2(G283), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n764), .A2(new_n440), .B1(new_n769), .B2(new_n219), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G97), .B2(new_n787), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n765), .A2(new_n355), .B1(new_n756), .B2(new_n211), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n317), .B(new_n833), .C1(G58), .C2(new_n787), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n835), .B2(new_n759), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT101), .Z(new_n837));
  AOI22_X1  g0637(.A1(G143), .A2(new_n773), .B1(new_n790), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n764), .C1(new_n288), .C2(new_n753), .ZN(new_n840));
  XOR2_X1   g0640(.A(new_n840), .B(KEYINPUT34), .Z(new_n841));
  OAI21_X1  g0641(.A(new_n832), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n750), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n821), .A2(new_n805), .A3(new_n823), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n820), .A2(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n432), .A2(new_n680), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n817), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(new_n678), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n391), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(new_n354), .B2(new_n406), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n330), .A2(new_n343), .A3(new_n345), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n853), .A2(new_n659), .B1(new_n346), .B2(new_n348), .ZN(new_n854));
  INV_X1    g0654(.A(new_n851), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n348), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n853), .A2(new_n857), .A3(new_n341), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(new_n402), .A4(new_n851), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n849), .B1(new_n852), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n853), .A2(KEYINPUT75), .A3(new_n857), .A4(new_n341), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n352), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n349), .A2(KEYINPUT75), .A3(KEYINPUT17), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n865), .A2(new_n406), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n855), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n863), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n388), .A2(new_n389), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n691), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n389), .A2(new_n680), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n390), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n848), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n664), .A2(new_n850), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT102), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n870), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n860), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT103), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n854), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n858), .A2(KEYINPUT103), .A3(new_n661), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n886), .A2(new_n887), .A3(new_n851), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n884), .B1(new_n888), .B2(KEYINPUT37), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n851), .B1(new_n354), .B2(new_n664), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n849), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(KEYINPUT39), .B1(new_n891), .B2(new_n869), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n871), .A2(new_n680), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n876), .A2(KEYINPUT102), .A3(new_n878), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n881), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n703), .A2(new_n711), .A3(new_n436), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n673), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n736), .A2(new_n730), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n728), .A2(KEYINPUT95), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT31), .A4(new_n680), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n715), .A2(new_n732), .A3(new_n733), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n874), .A2(new_n814), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI221_X4 g0707(.A(new_n849), .B1(new_n856), .B2(new_n860), .C1(new_n867), .C2(new_n855), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT38), .B1(new_n868), .B2(new_n861), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n901), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n851), .B1(new_n854), .B2(new_n885), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT103), .B1(new_n858), .B2(new_n661), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT37), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n865), .A2(new_n664), .A3(new_n866), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n914), .A2(new_n860), .B1(new_n855), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n869), .B1(new_n916), .B2(KEYINPUT38), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n905), .A4(new_n906), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n911), .A2(G330), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n436), .A2(G330), .A3(new_n905), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n911), .A2(new_n918), .A3(new_n436), .A4(new_n905), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n900), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n294), .B2(new_n802), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n219), .B1(new_n598), .B2(KEYINPUT35), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n926), .B(new_n231), .C1(KEYINPUT35), .C2(new_n598), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT36), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n323), .A2(G77), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n233), .A2(new_n929), .B1(G50), .B2(new_n211), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n930), .A2(G1), .A3(new_n205), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n925), .A2(new_n928), .A3(new_n931), .ZN(G367));
  OAI21_X1  g0732(.A(new_n631), .B1(new_n607), .B2(new_n691), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n617), .A2(new_n691), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT105), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n653), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n617), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n691), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n692), .A2(new_n618), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n563), .A2(new_n568), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n680), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n640), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n651), .A2(new_n944), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n948));
  XNOR2_X1  g0748(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT107), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n942), .A2(new_n950), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT106), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n936), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n689), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n955), .B(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n740), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n692), .A2(new_n690), .ZN(new_n960));
  INV_X1    g0760(.A(new_n935), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT44), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT110), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT44), .B1(new_n960), .B2(new_n961), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n960), .A2(new_n961), .ZN(new_n967));
  XNOR2_X1  g0767(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT109), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n964), .A2(new_n965), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n966), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(new_n689), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n624), .A2(new_n691), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n687), .B(new_n974), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(new_n808), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n959), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n694), .B(KEYINPUT41), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n803), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n958), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n795), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n799), .B1(new_n207), .B2(new_n562), .C1(new_n243), .C2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n355), .A2(new_n769), .B1(new_n756), .B2(new_n357), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G150), .A2(new_n773), .B1(new_n760), .B2(G137), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n211), .B2(new_n767), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n987), .C1(G159), .C2(new_n775), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n988), .B(new_n253), .C1(new_n216), .C2(new_n765), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G143), .B2(new_n782), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n775), .A2(G294), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n765), .A2(new_n219), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n992), .A2(KEYINPUT46), .B1(new_n440), .B2(new_n772), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(KEYINPUT46), .B2(new_n992), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n769), .A2(new_n583), .B1(new_n767), .B2(new_n553), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n995), .A2(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n756), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(G97), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n1000), .B(new_n317), .C1(new_n776), .C2(new_n759), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT112), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n998), .B(new_n1002), .C1(G311), .C2(new_n782), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n990), .B1(new_n991), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT47), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n750), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n805), .B(new_n984), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n947), .A2(new_n745), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n982), .A2(new_n1010), .ZN(G387));
  NAND2_X1  g0811(.A1(new_n959), .A2(new_n976), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n740), .A2(new_n977), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n694), .A3(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT113), .B(G150), .Z(new_n1015));
  AOI21_X1  g0815(.A(new_n317), .B1(new_n760), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n784), .A2(G77), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n292), .C2(new_n753), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G68), .B2(new_n790), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n773), .A2(G50), .B1(new_n787), .B2(new_n413), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n782), .A2(G159), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1019), .A2(new_n1021), .A3(new_n1000), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(G322), .A2(new_n782), .B1(new_n775), .B2(G311), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(new_n440), .B2(new_n769), .C1(new_n776), .C2(new_n772), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT48), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n583), .B2(new_n767), .C1(new_n528), .C2(new_n765), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT49), .Z(new_n1028));
  AOI21_X1  g0828(.A(new_n253), .B1(new_n760), .B2(G326), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n219), .B2(new_n756), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1023), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n750), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n344), .A2(new_n355), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT50), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n211), .A2(new_n357), .ZN(new_n1035));
  NOR4_X1   g0835(.A1(new_n1034), .A2(G45), .A3(new_n1035), .A4(new_n697), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n240), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n795), .B1(new_n1037), .B2(new_n263), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n207), .A2(new_n253), .A3(new_n697), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1036), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n207), .A2(G107), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n799), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n744), .B1(new_n685), .B2(new_n686), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1032), .A2(new_n805), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1014), .B(new_n1044), .C1(new_n803), .C2(new_n976), .ZN(G393));
  NAND2_X1  g0845(.A1(new_n973), .A2(new_n804), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n799), .B1(new_n207), .B2(new_n372), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n248), .B2(new_n795), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(G283), .A2(new_n784), .B1(new_n760), .B2(G322), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT115), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n753), .A2(new_n440), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n317), .B1(new_n769), .B2(new_n528), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1050), .A2(new_n757), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n219), .B2(new_n767), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n764), .A2(new_n776), .B1(new_n772), .B2(new_n824), .ZN(new_n1055));
  XOR2_X1   g0855(.A(new_n1055), .B(KEYINPUT52), .Z(new_n1056));
  OAI22_X1  g0856(.A1(new_n765), .A2(new_n211), .B1(new_n769), .B2(new_n292), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(G50), .B2(new_n775), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n787), .A2(G77), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G87), .A2(new_n999), .B1(new_n760), .B2(G143), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1058), .A2(new_n253), .A3(new_n1059), .A4(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(G159), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n764), .A2(new_n288), .B1(new_n772), .B2(new_n1062), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT51), .Z(new_n1064));
  OAI22_X1  g0864(.A1(new_n1054), .A2(new_n1056), .B1(new_n1061), .B2(new_n1064), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n809), .B(new_n1048), .C1(new_n1065), .C2(new_n750), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n936), .B2(new_n745), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1013), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n973), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n694), .B1(new_n973), .B2(new_n1068), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1046), .B(new_n1067), .C1(new_n1070), .C2(new_n1071), .ZN(G390));
  AOI21_X1  g0872(.A(new_n874), .B1(new_n817), .B2(new_n847), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n892), .A2(new_n883), .B1(new_n1073), .B2(new_n894), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n894), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n816), .A2(new_n691), .A3(new_n710), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n847), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n917), .B(new_n1075), .C1(new_n1078), .C2(new_n874), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1074), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n905), .A2(new_n906), .A3(G330), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n738), .A2(G330), .A3(new_n816), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1083), .A2(new_n874), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1074), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n803), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT116), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n764), .A2(new_n583), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n765), .A2(new_n222), .B1(new_n756), .B2(new_n211), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1059), .A2(new_n317), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G107), .C2(new_n775), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n372), .B2(new_n769), .C1(new_n528), .C2(new_n759), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1088), .B(new_n1092), .C1(G116), .C2(new_n773), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n753), .A2(new_n839), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n784), .A2(new_n1015), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT53), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n253), .B1(new_n759), .B2(new_n1097), .C1(new_n835), .C2(new_n772), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n782), .A2(G128), .B1(new_n999), .B2(G50), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1099), .B(new_n1100), .C1(new_n1062), .C2(new_n767), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  AOI211_X1 g0902(.A(new_n1094), .B(new_n1101), .C1(new_n790), .C2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n750), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n805), .B(new_n1104), .C1(new_n893), .C2(new_n743), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n292), .B2(new_n822), .ZN(new_n1106));
  OR3_X1    g0906(.A1(new_n1086), .A2(new_n1087), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1087), .B1(new_n1086), .B2(new_n1106), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1083), .A2(new_n874), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n1081), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n848), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n905), .A2(G330), .A3(new_n816), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n874), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n1078), .C1(new_n874), .C2(new_n1083), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n898), .A2(new_n673), .A3(new_n920), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1116), .B1(new_n1111), .B2(new_n1114), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1074), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1081), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1120), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n694), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1107), .A2(new_n1108), .A3(new_n1125), .ZN(G378));
  XOR2_X1   g0926(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1127));
  NAND2_X1  g0927(.A1(new_n312), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1127), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n672), .A2(new_n301), .A3(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n298), .A2(new_n850), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1130), .A2(new_n1128), .A3(new_n298), .A4(new_n850), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1135), .A2(new_n743), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n443), .A2(new_n253), .ZN(new_n1137));
  AOI211_X1 g0937(.A(G50), .B(new_n1137), .C1(new_n313), .C2(new_n274), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n769), .A2(new_n839), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n764), .A2(new_n1097), .B1(new_n767), .B2(new_n288), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT117), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(new_n784), .C2(new_n1102), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n835), .B2(new_n753), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G128), .B2(new_n773), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT59), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G159), .A2(new_n999), .B1(new_n760), .B2(G124), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1146), .A2(new_n313), .A3(new_n274), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1138), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n999), .A2(G58), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1017), .B(new_n1149), .C1(new_n583), .C2(new_n759), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n413), .B2(new_n790), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G116), .A2(new_n782), .B1(new_n775), .B2(G97), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n773), .A2(G107), .B1(new_n787), .B2(G68), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n1137), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT58), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1006), .B1(new_n1148), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n822), .A2(new_n355), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(new_n1136), .A2(new_n809), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1160), .A2(new_n911), .A3(G330), .A4(new_n918), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n919), .A2(new_n1135), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n897), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1161), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n880), .B(new_n877), .C1(new_n1073), .C2(new_n870), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT102), .B1(new_n876), .B2(new_n878), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1164), .A2(new_n895), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1159), .B1(new_n1169), .B2(new_n804), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1124), .A2(new_n1117), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n695), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1174), .B1(new_n1124), .B2(new_n1117), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT118), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1163), .A2(new_n1168), .A3(new_n1177), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n897), .A2(KEYINPUT118), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1171), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(G375));
  NOR2_X1   g0982(.A1(new_n767), .A2(new_n355), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1149), .B1(new_n835), .B2(new_n764), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G137), .C2(new_n773), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n775), .A2(new_n1102), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n760), .A2(G128), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n253), .B1(new_n769), .B2(new_n288), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G159), .B2(new_n784), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n765), .A2(new_n372), .B1(new_n756), .B2(new_n357), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n562), .A2(new_n767), .B1(new_n759), .B2(new_n440), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n317), .B1(new_n769), .B2(new_n553), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n764), .A2(new_n528), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n219), .B2(new_n753), .C1(new_n583), .C2(new_n772), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1006), .B1(new_n1190), .B2(new_n1196), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n809), .B(new_n1197), .C1(new_n211), .C2(new_n822), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n875), .A2(new_n743), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT119), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1115), .A2(new_n804), .B1(new_n1198), .B2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1111), .A2(new_n1116), .A3(new_n1114), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n979), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1201), .B1(new_n1203), .B2(new_n1120), .ZN(G381));
  NOR3_X1   g1004(.A1(G387), .A2(G384), .A3(G390), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(G375), .A2(G378), .ZN(new_n1206));
  INV_X1    g1006(.A(G381), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(G393), .A2(G396), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT120), .ZN(G407));
  NAND2_X1  g1010(.A1(new_n1206), .A2(new_n679), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(G407), .A2(G213), .A3(new_n1211), .ZN(G409));
  INV_X1    g1012(.A(G378), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1178), .A2(new_n804), .A3(new_n1179), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1159), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1214), .B(new_n1215), .C1(new_n980), .C2(new_n1173), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1213), .A2(new_n1216), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n1163), .A2(new_n1168), .B1(new_n1124), .B2(new_n1117), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n694), .B1(new_n1218), .B2(KEYINPUT57), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G378), .B(new_n1170), .C1(new_n1219), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT121), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n897), .B(new_n1164), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1116), .B1(new_n1225), .B2(new_n1120), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1174), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n1180), .A3(new_n694), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1228), .A2(KEYINPUT121), .A3(G378), .A4(new_n1170), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1217), .B1(new_n1223), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(G213), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G343), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1230), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT60), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1202), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n1118), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT122), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1202), .A2(new_n1234), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT122), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1235), .A2(new_n1239), .A3(new_n1118), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1237), .A2(new_n694), .A3(new_n1238), .A4(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1201), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT123), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(G384), .B(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n820), .A2(new_n844), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1241), .A2(new_n1243), .A3(new_n1246), .A4(new_n1201), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1233), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT62), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT61), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1232), .A2(G2897), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1245), .A2(new_n1247), .A3(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1253), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1230), .B2(new_n1232), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1233), .A2(new_n1258), .A3(new_n1248), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1250), .A2(new_n1251), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1009), .B1(new_n958), .B2(new_n981), .ZN(new_n1261));
  AND2_X1   g1061(.A1(G393), .A2(G396), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n1261), .A2(KEYINPUT124), .B1(new_n1208), .B2(new_n1262), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1208), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(G387), .A2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1263), .A2(new_n1265), .A3(G390), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G390), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1251), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1257), .A2(KEYINPUT63), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1249), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1217), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT121), .B1(new_n1181), .B2(G378), .ZN(new_n1274));
  AND4_X1   g1074(.A1(KEYINPUT121), .A2(new_n1228), .A3(G378), .A4(new_n1170), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1232), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1277), .A4(new_n1248), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT125), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1233), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1248), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1272), .A2(new_n1282), .A3(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1272), .B2(new_n1282), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1269), .B1(new_n1284), .B2(new_n1285), .ZN(G405));
  OAI22_X1  g1086(.A1(new_n1274), .A2(new_n1275), .B1(G378), .B2(new_n1181), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1248), .B1(new_n1287), .B2(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(KEYINPUT127), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1288), .B(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1268), .ZN(G402));
endmodule


