

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U549 ( .A(n692), .B(n691), .ZN(n695) );
  XNOR2_X1 U550 ( .A(n714), .B(n713), .ZN(n718) );
  INV_X1 U551 ( .A(KEYINPUT29), .ZN(n713) );
  NOR2_X1 U552 ( .A1(n733), .A2(n732), .ZN(n735) );
  NOR2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XNOR2_X2 U554 ( .A(KEYINPUT66), .B(n516), .ZN(n517) );
  OR2_X1 U555 ( .A1(G301), .A2(n719), .ZN(n513) );
  AND2_X1 U556 ( .A1(n808), .A2(n819), .ZN(n514) );
  INV_X1 U557 ( .A(KEYINPUT94), .ZN(n691) );
  OR2_X1 U558 ( .A1(n702), .A2(n962), .ZN(n708) );
  XNOR2_X1 U559 ( .A(n723), .B(KEYINPUT97), .ZN(n725) );
  AND2_X1 U560 ( .A1(n725), .A2(n724), .ZN(n726) );
  INV_X1 U561 ( .A(KEYINPUT31), .ZN(n728) );
  INV_X1 U562 ( .A(KEYINPUT99), .ZN(n734) );
  AND2_X1 U563 ( .A1(n966), .A2(n762), .ZN(n752) );
  NOR2_X1 U564 ( .A1(G543), .A2(n522), .ZN(n515) );
  NAND2_X1 U565 ( .A1(n514), .A2(n809), .ZN(n810) );
  XNOR2_X1 U566 ( .A(n595), .B(KEYINPUT15), .ZN(n962) );
  OR2_X1 U567 ( .A1(n811), .A2(n810), .ZN(n826) );
  NOR2_X1 U568 ( .A1(G651), .A2(n635), .ZN(n652) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n635) );
  NAND2_X1 U570 ( .A1(G51), .A2(n652), .ZN(n519) );
  INV_X1 U571 ( .A(G651), .ZN(n522) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n515), .Z(n516) );
  NAND2_X1 U573 ( .A1(G63), .A2(n517), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U575 ( .A(KEYINPUT6), .B(n520), .ZN(n527) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U577 ( .A1(n648), .A2(G89), .ZN(n521) );
  XNOR2_X1 U578 ( .A(n521), .B(KEYINPUT4), .ZN(n524) );
  NOR2_X1 U579 ( .A1(n635), .A2(n522), .ZN(n649) );
  NAND2_X1 U580 ( .A1(G76), .A2(n649), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U582 ( .A(n525), .B(KEYINPUT5), .Z(n526) );
  NOR2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U584 ( .A(KEYINPUT73), .B(n528), .Z(n529) );
  XOR2_X1 U585 ( .A(KEYINPUT7), .B(n529), .Z(G168) );
  INV_X1 U586 ( .A(G2105), .ZN(n532) );
  AND2_X1 U587 ( .A1(n532), .A2(G2104), .ZN(n883) );
  NAND2_X1 U588 ( .A1(G102), .A2(n883), .ZN(n531) );
  AND2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U590 ( .A1(G114), .A2(n879), .ZN(n530) );
  AND2_X1 U591 ( .A1(n531), .A2(n530), .ZN(n535) );
  NOR2_X1 U592 ( .A1(G2104), .A2(n532), .ZN(n551) );
  BUF_X1 U593 ( .A(n551), .Z(n878) );
  NAND2_X1 U594 ( .A1(n878), .A2(G126), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(KEYINPUT84), .ZN(n534) );
  AND2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n538) );
  XOR2_X2 U597 ( .A(KEYINPUT17), .B(n536), .Z(n882) );
  NAND2_X1 U598 ( .A1(n882), .A2(G138), .ZN(n537) );
  AND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(G164) );
  XOR2_X1 U600 ( .A(G2446), .B(G2430), .Z(n540) );
  XNOR2_X1 U601 ( .A(G2451), .B(G2454), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U603 ( .A(n541), .B(G2427), .Z(n543) );
  XNOR2_X1 U604 ( .A(G1348), .B(G1341), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(n547) );
  XOR2_X1 U606 ( .A(G2443), .B(KEYINPUT104), .Z(n545) );
  XNOR2_X1 U607 ( .A(G2438), .B(G2435), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U609 ( .A(n547), .B(n546), .Z(n548) );
  AND2_X1 U610 ( .A1(G14), .A2(n548), .ZN(G401) );
  NAND2_X1 U611 ( .A1(G135), .A2(n882), .ZN(n550) );
  NAND2_X1 U612 ( .A1(G111), .A2(n879), .ZN(n549) );
  NAND2_X1 U613 ( .A1(n550), .A2(n549), .ZN(n554) );
  BUF_X1 U614 ( .A(n551), .Z(n869) );
  NAND2_X1 U615 ( .A1(n869), .A2(G123), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT18), .B(n552), .Z(n553) );
  NOR2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n883), .A2(G99), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n999) );
  XNOR2_X1 U620 ( .A(G2096), .B(n999), .ZN(n557) );
  OR2_X1 U621 ( .A1(G2100), .A2(n557), .ZN(G156) );
  NAND2_X1 U622 ( .A1(G101), .A2(n883), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT23), .B(n558), .Z(n561) );
  NAND2_X1 U624 ( .A1(G125), .A2(n869), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT65), .B(n559), .Z(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G137), .A2(n882), .ZN(n563) );
  NAND2_X1 U628 ( .A1(G113), .A2(n879), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n686) );
  BUF_X1 U631 ( .A(n686), .Z(G160) );
  INV_X1 U632 ( .A(G108), .ZN(G238) );
  INV_X1 U633 ( .A(G132), .ZN(G219) );
  INV_X1 U634 ( .A(G82), .ZN(G220) );
  NAND2_X1 U635 ( .A1(G52), .A2(n652), .ZN(n567) );
  NAND2_X1 U636 ( .A1(G64), .A2(n517), .ZN(n566) );
  NAND2_X1 U637 ( .A1(n567), .A2(n566), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n648), .A2(G90), .ZN(n568) );
  XNOR2_X1 U639 ( .A(n568), .B(KEYINPUT68), .ZN(n570) );
  NAND2_X1 U640 ( .A1(G77), .A2(n649), .ZN(n569) );
  NAND2_X1 U641 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n571), .Z(n572) );
  NOR2_X1 U643 ( .A1(n573), .A2(n572), .ZN(G171) );
  NAND2_X1 U644 ( .A1(G94), .A2(G452), .ZN(n574) );
  XNOR2_X1 U645 ( .A(n574), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n575) );
  XNOR2_X1 U647 ( .A(n575), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n829) );
  NAND2_X1 U649 ( .A1(n829), .A2(G567), .ZN(n576) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n576), .Z(G234) );
  NAND2_X1 U651 ( .A1(n648), .A2(G81), .ZN(n577) );
  XNOR2_X1 U652 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U653 ( .A1(G68), .A2(n649), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n580), .B(KEYINPUT13), .ZN(n582) );
  NAND2_X1 U656 ( .A1(G43), .A2(n652), .ZN(n581) );
  NAND2_X1 U657 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n517), .A2(G56), .ZN(n583) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n583), .Z(n584) );
  NOR2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U661 ( .A(KEYINPUT71), .B(n586), .ZN(n972) );
  INV_X1 U662 ( .A(n972), .ZN(n587) );
  NAND2_X1 U663 ( .A1(n587), .A2(G860), .ZN(G153) );
  INV_X1 U664 ( .A(G171), .ZN(G301) );
  NAND2_X1 U665 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U666 ( .A1(G79), .A2(n649), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G54), .A2(n652), .ZN(n589) );
  NAND2_X1 U668 ( .A1(G92), .A2(n648), .ZN(n588) );
  NAND2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n517), .A2(G66), .ZN(n590) );
  XOR2_X1 U671 ( .A(KEYINPUT72), .B(n590), .Z(n591) );
  NOR2_X1 U672 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U674 ( .A(n962), .ZN(n608) );
  INV_X1 U675 ( .A(G868), .ZN(n612) );
  NAND2_X1 U676 ( .A1(n608), .A2(n612), .ZN(n596) );
  NAND2_X1 U677 ( .A1(n597), .A2(n596), .ZN(G284) );
  XOR2_X1 U678 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U679 ( .A1(G91), .A2(n648), .ZN(n599) );
  NAND2_X1 U680 ( .A1(G78), .A2(n649), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G53), .A2(n652), .ZN(n601) );
  NAND2_X1 U683 ( .A1(G65), .A2(n517), .ZN(n600) );
  NAND2_X1 U684 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U685 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U686 ( .A(KEYINPUT70), .B(n604), .Z(G299) );
  NOR2_X1 U687 ( .A1(G286), .A2(n612), .ZN(n606) );
  NOR2_X1 U688 ( .A1(G299), .A2(G868), .ZN(n605) );
  NOR2_X1 U689 ( .A1(n606), .A2(n605), .ZN(G297) );
  INV_X1 U690 ( .A(G559), .ZN(n610) );
  NOR2_X1 U691 ( .A1(G860), .A2(n610), .ZN(n607) );
  NOR2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U693 ( .A(KEYINPUT16), .B(n609), .Z(G148) );
  NAND2_X1 U694 ( .A1(n610), .A2(n962), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n611), .A2(G868), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n972), .A2(n612), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(G282) );
  NAND2_X1 U698 ( .A1(G559), .A2(n962), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n615), .B(KEYINPUT74), .ZN(n665) );
  XNOR2_X1 U700 ( .A(n665), .B(n972), .ZN(n616) );
  NOR2_X1 U701 ( .A1(n616), .A2(G860), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n652), .A2(G55), .ZN(n617) );
  XOR2_X1 U703 ( .A(KEYINPUT75), .B(n617), .Z(n619) );
  NAND2_X1 U704 ( .A1(G67), .A2(n517), .ZN(n618) );
  NAND2_X1 U705 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U706 ( .A(KEYINPUT76), .B(n620), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G93), .A2(n648), .ZN(n622) );
  NAND2_X1 U708 ( .A1(G80), .A2(n649), .ZN(n621) );
  NAND2_X1 U709 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n663) );
  XNOR2_X1 U711 ( .A(n625), .B(n663), .ZN(G145) );
  NAND2_X1 U712 ( .A1(n649), .A2(G73), .ZN(n627) );
  XNOR2_X1 U713 ( .A(KEYINPUT78), .B(KEYINPUT2), .ZN(n626) );
  XNOR2_X1 U714 ( .A(n627), .B(n626), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G48), .A2(n652), .ZN(n629) );
  NAND2_X1 U716 ( .A1(G86), .A2(n648), .ZN(n628) );
  NAND2_X1 U717 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U718 ( .A1(G61), .A2(n517), .ZN(n630) );
  XNOR2_X1 U719 ( .A(KEYINPUT77), .B(n630), .ZN(n631) );
  NOR2_X1 U720 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U722 ( .A1(G87), .A2(n635), .ZN(n637) );
  NAND2_X1 U723 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U725 ( .A1(n517), .A2(n638), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n652), .A2(G49), .ZN(n639) );
  NAND2_X1 U727 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U728 ( .A1(G85), .A2(n648), .ZN(n642) );
  NAND2_X1 U729 ( .A1(G72), .A2(n649), .ZN(n641) );
  NAND2_X1 U730 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G47), .A2(n652), .ZN(n643) );
  XNOR2_X1 U732 ( .A(KEYINPUT67), .B(n643), .ZN(n644) );
  NOR2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U734 ( .A1(G60), .A2(n517), .ZN(n646) );
  NAND2_X1 U735 ( .A1(n647), .A2(n646), .ZN(G290) );
  NAND2_X1 U736 ( .A1(G88), .A2(n648), .ZN(n651) );
  NAND2_X1 U737 ( .A1(G75), .A2(n649), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(n656) );
  NAND2_X1 U739 ( .A1(G50), .A2(n652), .ZN(n654) );
  NAND2_X1 U740 ( .A1(G62), .A2(n517), .ZN(n653) );
  NAND2_X1 U741 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U742 ( .A1(n656), .A2(n655), .ZN(G166) );
  NOR2_X1 U743 ( .A1(G868), .A2(n663), .ZN(n657) );
  XNOR2_X1 U744 ( .A(n657), .B(KEYINPUT79), .ZN(n668) );
  XNOR2_X1 U745 ( .A(KEYINPUT19), .B(G305), .ZN(n658) );
  XNOR2_X1 U746 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U747 ( .A(G299), .B(n659), .ZN(n661) );
  XNOR2_X1 U748 ( .A(G290), .B(G166), .ZN(n660) );
  XNOR2_X1 U749 ( .A(n661), .B(n660), .ZN(n662) );
  XOR2_X1 U750 ( .A(n663), .B(n662), .Z(n664) );
  XNOR2_X1 U751 ( .A(n972), .B(n664), .ZN(n853) );
  XNOR2_X1 U752 ( .A(n853), .B(n665), .ZN(n666) );
  NAND2_X1 U753 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U754 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n670), .ZN(n671) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n671), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n672), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n673) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n673), .Z(n674) );
  NOR2_X1 U763 ( .A1(G218), .A2(n674), .ZN(n675) );
  XNOR2_X1 U764 ( .A(KEYINPUT80), .B(n675), .ZN(n676) );
  NAND2_X1 U765 ( .A1(n676), .A2(G96), .ZN(n834) );
  NAND2_X1 U766 ( .A1(G2106), .A2(n834), .ZN(n677) );
  XOR2_X1 U767 ( .A(KEYINPUT81), .B(n677), .Z(n682) );
  NAND2_X1 U768 ( .A1(G69), .A2(G120), .ZN(n678) );
  XNOR2_X1 U769 ( .A(KEYINPUT82), .B(n678), .ZN(n679) );
  NOR2_X1 U770 ( .A1(G238), .A2(n679), .ZN(n680) );
  NAND2_X1 U771 ( .A1(G57), .A2(n680), .ZN(n835) );
  NAND2_X1 U772 ( .A1(G567), .A2(n835), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U774 ( .A(KEYINPUT83), .B(n683), .ZN(G319) );
  INV_X1 U775 ( .A(G319), .ZN(n906) );
  NAND2_X1 U776 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U777 ( .A1(n906), .A2(n684), .ZN(n833) );
  NAND2_X1 U778 ( .A1(n833), .A2(G36), .ZN(G176) );
  INV_X1 U779 ( .A(G166), .ZN(G303) );
  NOR2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n757) );
  NOR2_X1 U781 ( .A1(G1971), .A2(G303), .ZN(n685) );
  NOR2_X1 U782 ( .A1(n757), .A2(n685), .ZN(n966) );
  INV_X1 U783 ( .A(G299), .ZN(n969) );
  AND2_X1 U784 ( .A1(n686), .A2(G40), .ZN(n792) );
  NOR2_X1 U785 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NAND2_X1 U786 ( .A1(n792), .A2(n794), .ZN(n720) );
  INV_X1 U787 ( .A(n720), .ZN(n687) );
  INV_X1 U788 ( .A(n687), .ZN(n740) );
  NAND2_X1 U789 ( .A1(G1956), .A2(n740), .ZN(n690) );
  NAND2_X1 U790 ( .A1(n687), .A2(G2072), .ZN(n688) );
  XOR2_X1 U791 ( .A(KEYINPUT27), .B(n688), .Z(n689) );
  NAND2_X1 U792 ( .A1(n690), .A2(n689), .ZN(n692) );
  NOR2_X1 U793 ( .A1(n969), .A2(n695), .ZN(n694) );
  XNOR2_X1 U794 ( .A(KEYINPUT95), .B(KEYINPUT28), .ZN(n693) );
  XNOR2_X1 U795 ( .A(n694), .B(n693), .ZN(n712) );
  NAND2_X1 U796 ( .A1(n969), .A2(n695), .ZN(n710) );
  INV_X1 U797 ( .A(G1996), .ZN(n789) );
  NOR2_X1 U798 ( .A1(n720), .A2(n789), .ZN(n697) );
  XOR2_X1 U799 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n696) );
  XNOR2_X1 U800 ( .A(n697), .B(n696), .ZN(n699) );
  NAND2_X1 U801 ( .A1(n740), .A2(G1341), .ZN(n698) );
  NAND2_X1 U802 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U803 ( .A(KEYINPUT96), .B(n700), .ZN(n701) );
  NOR2_X1 U804 ( .A1(n701), .A2(n972), .ZN(n702) );
  NAND2_X1 U805 ( .A1(n702), .A2(n962), .ZN(n706) );
  NOR2_X1 U806 ( .A1(n687), .A2(G1348), .ZN(n704) );
  NOR2_X1 U807 ( .A1(G2067), .A2(n740), .ZN(n703) );
  NOR2_X1 U808 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U809 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U810 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U811 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U812 ( .A1(n712), .A2(n711), .ZN(n714) );
  XOR2_X1 U813 ( .A(G1961), .B(KEYINPUT92), .Z(n927) );
  NAND2_X1 U814 ( .A1(n927), .A2(n740), .ZN(n715) );
  XNOR2_X1 U815 ( .A(n715), .B(KEYINPUT93), .ZN(n717) );
  XOR2_X1 U816 ( .A(G2078), .B(KEYINPUT25), .Z(n946) );
  NOR2_X1 U817 ( .A1(n740), .A2(n946), .ZN(n716) );
  NOR2_X1 U818 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U819 ( .A1(n718), .A2(n513), .ZN(n731) );
  AND2_X1 U820 ( .A1(G301), .A2(n719), .ZN(n727) );
  NAND2_X1 U821 ( .A1(G8), .A2(n720), .ZN(n768) );
  NOR2_X1 U822 ( .A1(G1966), .A2(n768), .ZN(n732) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n740), .ZN(n736) );
  NOR2_X1 U824 ( .A1(n732), .A2(n736), .ZN(n721) );
  NAND2_X1 U825 ( .A1(G8), .A2(n721), .ZN(n722) );
  XNOR2_X1 U826 ( .A(KEYINPUT30), .B(n722), .ZN(n723) );
  INV_X1 U827 ( .A(G168), .ZN(n724) );
  NOR2_X1 U828 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U829 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U830 ( .A1(n731), .A2(n730), .ZN(n739) );
  XOR2_X1 U831 ( .A(KEYINPUT98), .B(n739), .Z(n733) );
  XNOR2_X1 U832 ( .A(n735), .B(n734), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n736), .A2(G8), .ZN(n737) );
  NAND2_X1 U834 ( .A1(n738), .A2(n737), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n739), .A2(G286), .ZN(n745) );
  NOR2_X1 U836 ( .A1(G1971), .A2(n768), .ZN(n742) );
  NOR2_X1 U837 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U838 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U840 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U841 ( .A1(n746), .A2(G8), .ZN(n747) );
  XNOR2_X1 U842 ( .A(n747), .B(KEYINPUT100), .ZN(n748) );
  XNOR2_X1 U843 ( .A(KEYINPUT32), .B(n748), .ZN(n749) );
  NAND2_X1 U844 ( .A1(n750), .A2(n749), .ZN(n762) );
  INV_X1 U845 ( .A(KEYINPUT101), .ZN(n751) );
  XNOR2_X1 U846 ( .A(n752), .B(n751), .ZN(n755) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n961) );
  INV_X1 U848 ( .A(n768), .ZN(n753) );
  NAND2_X1 U849 ( .A1(n961), .A2(n753), .ZN(n754) );
  NOR2_X1 U850 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U851 ( .A1(n756), .A2(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n757), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U853 ( .A1(n758), .A2(n768), .ZN(n759) );
  NOR2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n977) );
  AND2_X1 U856 ( .A1(n761), .A2(n977), .ZN(n773) );
  NOR2_X1 U857 ( .A1(G2090), .A2(G303), .ZN(n763) );
  NAND2_X1 U858 ( .A1(G8), .A2(n763), .ZN(n764) );
  NAND2_X1 U859 ( .A1(n762), .A2(n764), .ZN(n765) );
  NAND2_X1 U860 ( .A1(n765), .A2(n768), .ZN(n771) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XNOR2_X1 U862 ( .A(n766), .B(KEYINPUT24), .ZN(n767) );
  XNOR2_X1 U863 ( .A(n767), .B(KEYINPUT91), .ZN(n769) );
  OR2_X1 U864 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X1 U866 ( .A1(n773), .A2(n772), .ZN(n811) );
  NAND2_X1 U867 ( .A1(n883), .A2(G95), .ZN(n774) );
  XNOR2_X1 U868 ( .A(n774), .B(KEYINPUT88), .ZN(n776) );
  NAND2_X1 U869 ( .A1(G107), .A2(n879), .ZN(n775) );
  NAND2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U871 ( .A1(G119), .A2(n878), .ZN(n778) );
  NAND2_X1 U872 ( .A1(G131), .A2(n882), .ZN(n777) );
  NAND2_X1 U873 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n890) );
  AND2_X1 U875 ( .A1(n890), .A2(G1991), .ZN(n791) );
  NAND2_X1 U876 ( .A1(G117), .A2(n879), .ZN(n787) );
  NAND2_X1 U877 ( .A1(G129), .A2(n878), .ZN(n782) );
  NAND2_X1 U878 ( .A1(G141), .A2(n882), .ZN(n781) );
  NAND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n883), .A2(G105), .ZN(n783) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U883 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U884 ( .A(n788), .B(KEYINPUT89), .ZN(n894) );
  NOR2_X1 U885 ( .A1(n894), .A2(n789), .ZN(n790) );
  NOR2_X1 U886 ( .A1(n791), .A2(n790), .ZN(n991) );
  INV_X1 U887 ( .A(n792), .ZN(n793) );
  NOR2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n823) );
  INV_X1 U889 ( .A(n823), .ZN(n795) );
  NOR2_X1 U890 ( .A1(n991), .A2(n795), .ZN(n814) );
  XOR2_X1 U891 ( .A(KEYINPUT90), .B(n814), .Z(n808) );
  XNOR2_X1 U892 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NAND2_X1 U893 ( .A1(n883), .A2(G104), .ZN(n796) );
  XOR2_X1 U894 ( .A(KEYINPUT85), .B(n796), .Z(n798) );
  NAND2_X1 U895 ( .A1(n882), .A2(G140), .ZN(n797) );
  NAND2_X1 U896 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U897 ( .A(KEYINPUT34), .B(n799), .ZN(n806) );
  NAND2_X1 U898 ( .A1(n879), .A2(G116), .ZN(n800) );
  XNOR2_X1 U899 ( .A(n800), .B(KEYINPUT86), .ZN(n802) );
  NAND2_X1 U900 ( .A1(G128), .A2(n869), .ZN(n801) );
  NAND2_X1 U901 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U902 ( .A(KEYINPUT35), .B(n803), .ZN(n804) );
  XNOR2_X1 U903 ( .A(KEYINPUT87), .B(n804), .ZN(n805) );
  NOR2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n807), .ZN(n901) );
  NOR2_X1 U906 ( .A1(n821), .A2(n901), .ZN(n1005) );
  NAND2_X1 U907 ( .A1(n823), .A2(n1005), .ZN(n819) );
  XNOR2_X1 U908 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U909 ( .A1(n968), .A2(n823), .ZN(n809) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n890), .ZN(n1002) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U912 ( .A1(n1002), .A2(n812), .ZN(n813) );
  NOR2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n817) );
  INV_X1 U914 ( .A(n894), .ZN(n815) );
  NOR2_X1 U915 ( .A1(n815), .A2(G1996), .ZN(n816) );
  XNOR2_X1 U916 ( .A(n816), .B(KEYINPUT102), .ZN(n993) );
  NOR2_X1 U917 ( .A1(n817), .A2(n993), .ZN(n818) );
  XNOR2_X1 U918 ( .A(n818), .B(KEYINPUT39), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n821), .A2(n901), .ZN(n990) );
  NAND2_X1 U921 ( .A1(n822), .A2(n990), .ZN(n824) );
  NAND2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(n828) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n829), .ZN(G217) );
  NAND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n830) );
  XNOR2_X1 U928 ( .A(KEYINPUT105), .B(n830), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n831), .A2(G661), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U931 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U932 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  XNOR2_X1 U933 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n837) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2072), .Z(n839) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U944 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1976), .B(G1981), .Z(n845) );
  XNOR2_X1 U948 ( .A(G1971), .B(G1966), .ZN(n844) );
  XNOR2_X1 U949 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U950 ( .A(n846), .B(G2474), .Z(n848) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1956), .Z(n850) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1961), .ZN(n849) );
  XNOR2_X1 U955 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(G229) );
  XOR2_X1 U957 ( .A(KEYINPUT114), .B(n853), .Z(n855) );
  XNOR2_X1 U958 ( .A(G171), .B(n962), .ZN(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n856), .B(G286), .ZN(n857) );
  NOR2_X1 U961 ( .A1(G37), .A2(n857), .ZN(G397) );
  NAND2_X1 U962 ( .A1(G100), .A2(n883), .ZN(n859) );
  NAND2_X1 U963 ( .A1(G112), .A2(n879), .ZN(n858) );
  NAND2_X1 U964 ( .A1(n859), .A2(n858), .ZN(n867) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n861) );
  NAND2_X1 U966 ( .A1(G124), .A2(n869), .ZN(n860) );
  XNOR2_X1 U967 ( .A(n861), .B(n860), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n882), .A2(G136), .ZN(n862) );
  XNOR2_X1 U969 ( .A(KEYINPUT109), .B(n862), .ZN(n863) );
  NOR2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U971 ( .A(KEYINPUT110), .B(n865), .Z(n866) );
  NOR2_X1 U972 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U973 ( .A1(n879), .A2(G115), .ZN(n868) );
  XNOR2_X1 U974 ( .A(n868), .B(KEYINPUT112), .ZN(n871) );
  NAND2_X1 U975 ( .A1(G127), .A2(n869), .ZN(n870) );
  NAND2_X1 U976 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U977 ( .A(n872), .B(KEYINPUT47), .ZN(n874) );
  NAND2_X1 U978 ( .A1(G139), .A2(n882), .ZN(n873) );
  NAND2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G103), .A2(n883), .ZN(n875) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n875), .ZN(n876) );
  NOR2_X1 U982 ( .A1(n877), .A2(n876), .ZN(n995) );
  NAND2_X1 U983 ( .A1(G130), .A2(n878), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G118), .A2(n879), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U986 ( .A1(G142), .A2(n882), .ZN(n885) );
  NAND2_X1 U987 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U988 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U989 ( .A(KEYINPUT45), .B(n886), .Z(n887) );
  NOR2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U991 ( .A(n995), .B(n889), .ZN(n900) );
  XNOR2_X1 U992 ( .A(G164), .B(G162), .ZN(n898) );
  XOR2_X1 U993 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n892) );
  XOR2_X1 U994 ( .A(n890), .B(KEYINPUT113), .Z(n891) );
  XNOR2_X1 U995 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U996 ( .A(n999), .B(n893), .ZN(n896) );
  XNOR2_X1 U997 ( .A(G160), .B(n894), .ZN(n895) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n902), .B(n901), .Z(n903) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n903), .ZN(G395) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n905), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G397), .A2(n906), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(n909), .A2(G395), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(n910), .B(KEYINPUT115), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U1012 ( .A(G1971), .B(G22), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(G23), .B(G1976), .ZN(n911) );
  NOR2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1015 ( .A(KEYINPUT126), .B(n913), .Z(n915) );
  XNOR2_X1 U1016 ( .A(G1986), .B(G24), .ZN(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(KEYINPUT58), .B(n916), .ZN(n932) );
  XNOR2_X1 U1019 ( .A(G1348), .B(KEYINPUT59), .ZN(n917) );
  XNOR2_X1 U1020 ( .A(n917), .B(G4), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(G1956), .B(G20), .ZN(n919) );
  XNOR2_X1 U1022 ( .A(G6), .B(G1981), .ZN(n918) );
  NOR2_X1 U1023 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1024 ( .A1(n921), .A2(n920), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G19), .B(G1341), .ZN(n922) );
  XNOR2_X1 U1026 ( .A(KEYINPUT124), .B(n922), .ZN(n923) );
  NOR2_X1 U1027 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1028 ( .A(n925), .B(KEYINPUT60), .ZN(n926) );
  XNOR2_X1 U1029 ( .A(n926), .B(KEYINPUT125), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(n927), .B(G5), .ZN(n928) );
  XNOR2_X1 U1031 ( .A(KEYINPUT123), .B(n928), .ZN(n929) );
  NOR2_X1 U1032 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(G21), .B(G1966), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1036 ( .A(KEYINPUT61), .B(n935), .Z(n936) );
  NOR2_X1 U1037 ( .A1(G16), .A2(n936), .ZN(n988) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n956) );
  XOR2_X1 U1039 ( .A(G2084), .B(G34), .Z(n937) );
  XNOR2_X1 U1040 ( .A(KEYINPUT54), .B(n937), .ZN(n953) );
  XNOR2_X1 U1041 ( .A(G2090), .B(G35), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n939) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n938) );
  NOR2_X1 U1044 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1045 ( .A(G2067), .B(G26), .Z(n940) );
  NAND2_X1 U1046 ( .A1(n940), .A2(G28), .ZN(n943) );
  XNOR2_X1 U1047 ( .A(G25), .B(G1991), .ZN(n941) );
  XNOR2_X1 U1048 ( .A(KEYINPUT118), .B(n941), .ZN(n942) );
  NOR2_X1 U1049 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1050 ( .A1(n945), .A2(n944), .ZN(n948) );
  XNOR2_X1 U1051 ( .A(G27), .B(n946), .ZN(n947) );
  NOR2_X1 U1052 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n949), .ZN(n950) );
  NOR2_X1 U1054 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1055 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1056 ( .A(n954), .B(KEYINPUT119), .ZN(n955) );
  XNOR2_X1 U1057 ( .A(n956), .B(n955), .ZN(n957) );
  INV_X1 U1058 ( .A(G29), .ZN(n1016) );
  NAND2_X1 U1059 ( .A1(n957), .A2(n1016), .ZN(n958) );
  NAND2_X1 U1060 ( .A1(G11), .A2(n958), .ZN(n959) );
  XNOR2_X1 U1061 ( .A(n959), .B(KEYINPUT121), .ZN(n986) );
  NAND2_X1 U1062 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NAND2_X1 U1063 ( .A1(n961), .A2(n960), .ZN(n964) );
  XOR2_X1 U1064 ( .A(G1348), .B(n962), .Z(n963) );
  NOR2_X1 U1065 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  NOR2_X1 U1067 ( .A1(n968), .A2(n967), .ZN(n976) );
  XNOR2_X1 U1068 ( .A(G171), .B(G1961), .ZN(n971) );
  XNOR2_X1 U1069 ( .A(n969), .B(G1956), .ZN(n970) );
  NAND2_X1 U1070 ( .A1(n971), .A2(n970), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n972), .ZN(n973) );
  NOR2_X1 U1072 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G168), .B(G1966), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n979), .Z(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1078 ( .A(KEYINPUT122), .B(n982), .Z(n984) );
  XNOR2_X1 U1079 ( .A(G16), .B(KEYINPUT56), .ZN(n983) );
  NAND2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1081 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n989), .B(KEYINPUT127), .ZN(n1018) );
  NAND2_X1 U1084 ( .A1(n991), .A2(n990), .ZN(n1012) );
  XOR2_X1 U1085 ( .A(G2090), .B(G162), .Z(n992) );
  NOR2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1087 ( .A(KEYINPUT51), .B(n994), .Z(n1010) );
  XOR2_X1 U1088 ( .A(G2072), .B(n995), .Z(n997) );
  XOR2_X1 U1089 ( .A(G164), .B(G2078), .Z(n996) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1091 ( .A(KEYINPUT50), .B(n998), .Z(n1008) );
  XNOR2_X1 U1092 ( .A(G160), .B(G2084), .ZN(n1000) );
  NAND2_X1 U1093 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1095 ( .A(KEYINPUT116), .B(n1003), .Z(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT117), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(KEYINPUT52), .B(n1013), .Z(n1014) );
  NOR2_X1 U1102 ( .A1(KEYINPUT55), .A2(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1019), .ZN(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

