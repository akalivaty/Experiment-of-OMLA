//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(new_n202));
  XNOR2_X1  g0002(.A(new_n202), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0003(.A1(G1), .A2(G20), .ZN(new_n204));
  INV_X1    g0004(.A(G87), .ZN(new_n205));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G257), .ZN(new_n208));
  OAI22_X1  g0008(.A1(new_n205), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g0009(.A(new_n209), .B1(G68), .B2(G238), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n213), .B1(G116), .B2(G270), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  INV_X1    g0015(.A(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n214), .B1(new_n215), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n204), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n204), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT65), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT0), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n224), .A2(new_n230), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G226), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(new_n212), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G270), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  OAI21_X1  g0051(.A(G20), .B1(new_n226), .B2(G50), .ZN(new_n252));
  INV_X1    g0052(.A(G150), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n228), .A2(G33), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n252), .B1(new_n253), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n229), .ZN(new_n260));
  INV_X1    g0060(.A(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n261), .A2(new_n228), .A3(G1), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n258), .A2(new_n260), .B1(new_n215), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n270));
  INV_X1    g0070(.A(G274), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n278), .A2(new_n279), .A3(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  OAI21_X1  g0081(.A(KEYINPUT67), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(G223), .A3(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G222), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n281), .ZN(new_n285));
  OAI221_X1 g0085(.A(new_n283), .B1(new_n217), .B2(new_n278), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n272), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n287), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n270), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n290), .A2(new_n216), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n269), .B1(new_n293), .B2(G200), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  AOI211_X1 g0096(.A(new_n272), .B(new_n291), .C1(new_n286), .C2(new_n287), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n296), .B1(new_n297), .B2(G190), .ZN(new_n298));
  AND4_X1   g0098(.A1(new_n296), .A2(new_n288), .A3(G190), .A4(new_n292), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n294), .B(new_n295), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G200), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(KEYINPUT10), .A3(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT10), .B1(new_n302), .B2(KEYINPUT72), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT71), .B1(new_n293), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n297), .A2(new_n296), .A3(G190), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n305), .A2(new_n309), .A3(new_n295), .A4(new_n294), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  OAI22_X1  g0111(.A1(new_n257), .A2(new_n255), .B1(new_n228), .B2(new_n217), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n256), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n260), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT69), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n265), .A2(G77), .ZN(new_n317));
  INV_X1    g0117(.A(new_n262), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(G77), .C2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n320), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n280), .A2(G238), .A3(new_n282), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n324), .B1(new_n211), .B2(new_n278), .C1(new_n221), .C2(new_n285), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n287), .ZN(new_n326));
  INV_X1    g0126(.A(new_n272), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n289), .A2(G244), .A3(new_n270), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n323), .B1(G190), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n267), .B1(new_n297), .B2(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT68), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n297), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT68), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n267), .C1(new_n297), .C2(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n335), .A2(new_n337), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G169), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n329), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n330), .A2(new_n336), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n323), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n311), .A2(new_n333), .A3(new_n340), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT73), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n255), .A2(new_n215), .B1(new_n228), .B2(G68), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n256), .A2(new_n217), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n260), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT11), .ZN(new_n350));
  INV_X1    g0150(.A(new_n265), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n262), .A2(new_n225), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n352), .A2(KEYINPUT12), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(KEYINPUT12), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n350), .B1(new_n225), .B2(new_n351), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(G33), .A2(G97), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n221), .A2(G1698), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G226), .B2(G1698), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(new_n277), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n272), .B1(new_n359), .B2(new_n287), .ZN(new_n360));
  INV_X1    g0160(.A(G238), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n290), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(KEYINPUT13), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n341), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  XOR2_X1   g0166(.A(new_n366), .B(KEYINPUT14), .Z(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(KEYINPUT74), .A3(new_n365), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT74), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n362), .A2(new_n369), .A3(KEYINPUT13), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n336), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n355), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n301), .B1(new_n364), .B2(new_n365), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n370), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n374), .B(new_n355), .C1(new_n375), .C2(G190), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n340), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n378), .B1(new_n304), .B2(new_n310), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(new_n333), .A4(new_n344), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n228), .B1(new_n226), .B2(new_n382), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n383), .A2(KEYINPUT77), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n254), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n383), .A2(KEYINPUT77), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n273), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT75), .B1(new_n273), .B2(KEYINPUT3), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n276), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n391), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n395), .B1(new_n275), .B2(G33), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n273), .A2(KEYINPUT75), .A3(KEYINPUT3), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n393), .B1(new_n398), .B2(G20), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n392), .A2(new_n399), .A3(KEYINPUT76), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT76), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n393), .C1(new_n398), .C2(G20), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G68), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT16), .B(new_n388), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT78), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n277), .B2(new_n228), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n393), .B(G20), .C1(new_n274), .C2(new_n276), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT79), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT79), .B(G68), .C1(new_n406), .C2(new_n407), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n388), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n402), .A2(G68), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n392), .A2(new_n399), .A3(KEYINPUT76), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT78), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(new_n418), .A3(KEYINPUT16), .A4(new_n388), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n405), .A2(new_n260), .A3(new_n414), .A4(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n327), .B1(new_n290), .B2(new_n221), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n216), .A2(G1698), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n398), .B(new_n424), .C1(G223), .C2(G1698), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n289), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(new_n421), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n429), .A2(G190), .B1(G200), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n318), .A2(new_n257), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n432), .B1(new_n265), .B2(new_n257), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n420), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT17), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n420), .A2(new_n433), .ZN(new_n437));
  OAI22_X1  g0237(.A1(new_n429), .A2(G179), .B1(G169), .B2(new_n430), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT18), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n346), .A2(new_n377), .A3(new_n381), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n398), .A2(KEYINPUT22), .A3(G87), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G33), .A2(G116), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n228), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n277), .A2(G20), .A3(new_n205), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(KEYINPUT22), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n228), .A2(G107), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n452), .B(KEYINPUT23), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT24), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n448), .A2(KEYINPUT24), .A3(new_n451), .A4(new_n453), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(new_n260), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n262), .A2(new_n211), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT25), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n398), .B1(G257), .B2(new_n281), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G250), .A2(G1698), .ZN(new_n464));
  INV_X1    g0264(.A(G294), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n463), .A2(new_n464), .B1(new_n273), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(G45), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(G1), .ZN(new_n468));
  AND2_X1   g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n289), .A2(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n466), .A2(new_n287), .B1(G264), .B2(new_n472), .ZN(new_n473));
  OR2_X1    g0273(.A1(new_n471), .A2(new_n271), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G200), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(G190), .ZN(new_n478));
  INV_X1    g0278(.A(new_n260), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n318), .B(new_n479), .C1(G1), .C2(new_n273), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G107), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n462), .A2(new_n477), .A3(new_n478), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n207), .A2(new_n211), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n211), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n489), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n490));
  OAI21_X1  g0290(.A(G107), .B1(new_n406), .B2(new_n407), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n479), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n480), .A2(new_n207), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n318), .A2(G97), .ZN(new_n494));
  OR3_X1    g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n391), .B2(new_n218), .ZN(new_n497));
  OAI21_X1  g0297(.A(KEYINPUT4), .B1(new_n277), .B2(new_n206), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n278), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n497), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n287), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n472), .A2(G257), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n503), .A2(new_n336), .A3(new_n474), .A4(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n503), .A2(new_n474), .A3(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n495), .B(new_n505), .C1(new_n506), .C2(G169), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n503), .A2(G190), .A3(new_n474), .A4(new_n504), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n509), .C1(new_n506), .C2(new_n301), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n208), .A2(new_n281), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n212), .A2(G1698), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n398), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n277), .A2(G303), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT87), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(KEYINPUT87), .A3(new_n516), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n287), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n474), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(G270), .B2(new_n472), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(G190), .A3(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n500), .B(new_n228), .C1(G33), .C2(new_n207), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n525), .B(new_n260), .C1(new_n228), .C2(G116), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT20), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n526), .B(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n481), .A2(G116), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(new_n529), .C1(G116), .C2(new_n318), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n301), .B1(new_n521), .B2(new_n523), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT88), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n533), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT88), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n524), .A4(new_n531), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n483), .A2(new_n512), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n458), .A2(new_n482), .A3(new_n461), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n476), .A2(new_n341), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n475), .A2(new_n336), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n521), .A2(new_n523), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n531), .A2(new_n544), .A3(new_n336), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(G169), .A3(new_n530), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT21), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT21), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n544), .A2(new_n548), .A3(G169), .A4(new_n530), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n545), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n287), .B1(G274), .B2(new_n468), .ZN(new_n553));
  OAI21_X1  g0353(.A(G250), .B1(new_n467), .B2(G1), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n446), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n396), .A2(new_n397), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n557), .A2(G244), .A3(G1698), .A4(new_n276), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT82), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT82), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n398), .A2(new_n560), .A3(G244), .A4(G1698), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n556), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n557), .A2(G238), .A3(new_n281), .A4(new_n276), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(KEYINPUT81), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT81), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n398), .A2(new_n565), .A3(G238), .A4(new_n281), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n562), .A2(KEYINPUT83), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT83), .B1(new_n562), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n555), .B1(new_n570), .B2(new_n287), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT86), .B1(new_n571), .B2(new_n306), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n559), .A2(new_n561), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n567), .A3(new_n446), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n562), .A2(KEYINPUT83), .A3(new_n567), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n287), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n555), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(G200), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n398), .A2(new_n228), .A3(G68), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n228), .B1(new_n356), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n486), .A2(new_n205), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n582), .B1(new_n256), .B2(new_n207), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(new_n260), .B1(new_n262), .B2(new_n313), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n481), .A2(G87), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n580), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n578), .A2(new_n579), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT86), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n593), .A3(G190), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n572), .A2(new_n591), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT84), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n578), .A2(G169), .A3(new_n579), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n336), .B1(new_n578), .B2(new_n579), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n578), .A2(G169), .A3(new_n579), .ZN(new_n600));
  OAI211_X1 g0400(.A(KEYINPUT84), .B(new_n600), .C1(new_n571), .C2(new_n336), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n588), .B1(new_n313), .B2(new_n480), .ZN(new_n602));
  XOR2_X1   g0402(.A(new_n602), .B(KEYINPUT85), .Z(new_n603));
  NAND3_X1  g0403(.A1(new_n599), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AND4_X1   g0404(.A1(new_n539), .A2(new_n552), .A3(new_n595), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n444), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT89), .ZN(G372));
  AOI21_X1  g0407(.A(new_n438), .B1(new_n420), .B2(new_n433), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n608), .B(KEYINPUT18), .ZN(new_n609));
  INV_X1    g0409(.A(new_n376), .ZN(new_n610));
  INV_X1    g0410(.A(new_n344), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n373), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n612), .B2(new_n436), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n378), .B1(new_n613), .B2(new_n311), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n478), .A2(new_n482), .A3(new_n461), .A4(new_n458), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n511), .B1(new_n615), .B2(new_n477), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n603), .B1(new_n597), .B2(new_n598), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n595), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n595), .A2(new_n616), .A3(KEYINPUT90), .A4(new_n617), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n551), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n507), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n604), .A2(new_n623), .A3(new_n595), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT26), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT26), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n595), .A2(new_n626), .A3(new_n623), .A4(new_n617), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n617), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n614), .B1(new_n443), .B2(new_n629), .ZN(G369));
  INV_X1    g0430(.A(new_n550), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n261), .A2(G20), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n264), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(KEYINPUT27), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(G213), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G343), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n530), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g0439(.A(new_n639), .B(KEYINPUT91), .Z(new_n640));
  NOR2_X1   g0440(.A1(new_n631), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n538), .A2(new_n550), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(G330), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n543), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n540), .A2(new_n638), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n483), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n543), .A2(new_n638), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n550), .A2(new_n638), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(new_n649), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n651), .A2(new_n655), .ZN(G399));
  INV_X1    g0456(.A(new_n231), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(G41), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n584), .A2(G116), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G1), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n227), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT29), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n595), .A2(new_n623), .A3(new_n617), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n604), .A2(new_n626), .A3(new_n595), .A4(new_n623), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n595), .A2(new_n616), .A3(new_n551), .A4(new_n617), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n666), .A2(new_n617), .A3(new_n667), .A4(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n638), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n627), .A2(new_n617), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(KEYINPUT26), .B2(new_n624), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n620), .A2(new_n551), .A3(new_n621), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n638), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n675), .B2(new_n664), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n571), .A2(KEYINPUT92), .A3(new_n336), .A4(new_n544), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n475), .A2(new_n506), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n578), .A2(new_n336), .A3(new_n544), .A4(new_n579), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT92), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n503), .A2(new_n474), .A3(new_n504), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n544), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n592), .A2(G179), .A3(new_n473), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n598), .A2(KEYINPUT30), .A3(new_n473), .A4(new_n684), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT31), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n689), .A2(new_n690), .A3(new_n638), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n689), .B2(new_n638), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n539), .A2(new_n552), .A3(new_n595), .A4(new_n604), .ZN(new_n693));
  OAI22_X1  g0493(.A1(new_n691), .A2(new_n692), .B1(new_n693), .B2(new_n638), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G330), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n676), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n663), .B1(new_n697), .B2(G1), .ZN(G364));
  NAND2_X1  g0498(.A1(new_n632), .A2(G45), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n659), .A2(G1), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n643), .A2(G330), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n645), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G13), .A2(G33), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G20), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n701), .B1(new_n643), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n229), .B1(G20), .B2(new_n341), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n228), .A2(G190), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G179), .A2(G200), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n278), .B1(new_n714), .B2(G329), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n336), .A2(new_n301), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n711), .ZN(new_n717));
  XOR2_X1   g0517(.A(KEYINPUT33), .B(G317), .Z(new_n718));
  OAI21_X1  g0518(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n336), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n711), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G311), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n228), .B1(new_n712), .B2(G190), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n721), .A2(new_n722), .B1(new_n723), .B2(new_n465), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n228), .A2(new_n306), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n716), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n724), .B1(G326), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT94), .Z(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n720), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n719), .B(new_n729), .C1(G322), .C2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G283), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n301), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n711), .ZN(new_n735));
  INV_X1    g0535(.A(G303), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n725), .A2(new_n734), .ZN(new_n737));
  OAI221_X1 g0537(.A(new_n732), .B1(new_n733), .B2(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n737), .A2(new_n205), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n726), .A2(new_n215), .B1(new_n723), .B2(new_n207), .ZN(new_n740));
  AOI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(G58), .C2(new_n731), .ZN(new_n741));
  INV_X1    g0541(.A(new_n717), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G68), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n278), .B1(new_n721), .B2(new_n217), .ZN(new_n744));
  INV_X1    g0544(.A(new_n735), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n744), .B1(G107), .B2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G159), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n713), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n741), .A2(new_n743), .A3(new_n746), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n710), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g0552(.A1(G355), .A2(new_n231), .A3(new_n278), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n247), .A2(new_n467), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n398), .A2(new_n657), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(G45), .B2(new_n227), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n753), .B1(G116), .B2(new_n231), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n706), .A2(new_n709), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n708), .A2(new_n752), .A3(new_n759), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n703), .A2(new_n760), .ZN(G396));
  NOR2_X1   g0561(.A1(new_n344), .A2(new_n638), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n323), .A2(new_n638), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n333), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n762), .B1(new_n764), .B2(new_n344), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n675), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n670), .B(new_n765), .C1(new_n622), .C2(new_n628), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OR3_X1    g0568(.A1(new_n766), .A2(new_n768), .A3(new_n695), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n695), .B1(new_n766), .B2(new_n768), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n769), .A2(new_n700), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n762), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n331), .A2(new_n332), .B1(new_n323), .B2(new_n638), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n772), .B1(new_n773), .B2(new_n611), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n704), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n709), .A2(new_n704), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n217), .ZN(new_n777));
  INV_X1    g0577(.A(new_n721), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G143), .A2(new_n731), .B1(new_n778), .B2(G159), .ZN(new_n779));
  INV_X1    g0579(.A(G137), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n779), .B1(new_n780), .B2(new_n726), .C1(new_n253), .C2(new_n717), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT34), .Z(new_n782));
  NOR2_X1   g0582(.A1(new_n735), .A2(new_n225), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n737), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n391), .B1(G50), .B2(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n784), .B(new_n786), .C1(new_n220), .C2(new_n723), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G132), .B2(new_n714), .ZN(new_n788));
  INV_X1    g0588(.A(G116), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n726), .A2(new_n736), .B1(new_n721), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n790), .B1(G283), .B2(new_n742), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT95), .Z(new_n792));
  OAI22_X1  g0592(.A1(new_n730), .A2(new_n465), .B1(new_n735), .B2(new_n205), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n723), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n278), .B1(new_n795), .B2(G97), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n794), .B(new_n796), .C1(new_n211), .C2(new_n737), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(G311), .B2(new_n714), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n709), .B1(new_n788), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n775), .A2(new_n701), .A3(new_n777), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n771), .A2(new_n800), .ZN(G384));
  AOI21_X1  g0601(.A(new_n789), .B1(new_n489), .B2(KEYINPUT35), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n229), .A2(new_n228), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(KEYINPUT35), .C2(new_n489), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT36), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n382), .A2(G77), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n227), .A2(new_n806), .B1(G50), .B2(new_n225), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G1), .A3(new_n261), .ZN(new_n808));
  AND3_X1   g0608(.A1(new_n420), .A2(new_n431), .A3(new_n433), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n636), .B1(new_n420), .B2(new_n433), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n440), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n812), .A2(KEYINPUT37), .ZN(new_n813));
  INV_X1    g0613(.A(new_n636), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n437), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n440), .A2(new_n815), .A3(new_n816), .A4(new_n434), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT98), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n818), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n813), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n810), .B1(new_n436), .B2(new_n441), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT38), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n817), .A2(new_n818), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n811), .A2(KEYINPUT98), .A3(new_n816), .A4(new_n440), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n387), .B1(new_n415), .B2(new_n416), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n413), .B1(new_n826), .B2(KEYINPUT97), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n827), .B1(KEYINPUT97), .B2(new_n826), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n405), .A2(new_n260), .A3(new_n419), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n433), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n814), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n439), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n831), .A2(new_n832), .A3(new_n434), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n824), .A2(new_n825), .B1(new_n833), .B2(KEYINPUT37), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n831), .B1(new_n609), .B2(new_n435), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n823), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n373), .A2(new_n638), .ZN(new_n839));
  INV_X1    g0639(.A(new_n355), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT96), .B1(new_n840), .B2(new_n670), .ZN(new_n841));
  OR3_X1    g0641(.A1(new_n840), .A2(KEYINPUT96), .A3(new_n670), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n372), .A2(new_n610), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  AND3_X1   g0644(.A1(new_n694), .A2(new_n765), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n838), .A2(KEYINPUT40), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n819), .B2(new_n820), .ZN(new_n848));
  INV_X1    g0648(.A(new_n836), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT38), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT99), .B1(new_n850), .B2(new_n837), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n848), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT99), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n851), .A2(new_n845), .A3(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT100), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  OAI211_X1 g0660(.A(G330), .B(new_n846), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(G330), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n677), .A2(new_n678), .A3(new_n681), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n687), .A2(new_n688), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n638), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT31), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n689), .A2(new_n690), .A3(new_n638), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n605), .A2(new_n670), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n862), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n444), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n861), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g0672(.A(new_n872), .B(KEYINPUT101), .Z(new_n873));
  INV_X1    g0673(.A(new_n846), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n856), .A2(new_n858), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT100), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND3_X1   g0678(.A1(new_n878), .A2(new_n444), .A3(new_n694), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n851), .A2(new_n855), .ZN(new_n880));
  INV_X1    g0680(.A(new_n844), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n767), .B2(new_n772), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n880), .A2(new_n882), .B1(new_n441), .B2(new_n636), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT39), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n884), .B1(new_n823), .B2(new_n837), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n372), .A2(new_n638), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n852), .A2(new_n853), .A3(KEYINPUT39), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n676), .A2(new_n443), .ZN(new_n890));
  INV_X1    g0690(.A(new_n614), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n889), .B(new_n892), .Z(new_n893));
  INV_X1    g0693(.A(KEYINPUT102), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n873), .A2(new_n879), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n632), .A2(new_n264), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n805), .B(new_n808), .C1(new_n897), .C2(new_n898), .ZN(G367));
  OAI21_X1  g0699(.A(new_n512), .B1(new_n509), .B2(new_n670), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n654), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT103), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n902), .A2(KEYINPUT42), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n507), .B1(new_n900), .B2(new_n543), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n670), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n595), .B(new_n617), .C1(new_n590), .C2(new_n670), .ZN(new_n909));
  OR3_X1    g0709(.A1(new_n617), .A2(new_n590), .A3(new_n670), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT43), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT104), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n912), .A3(new_n910), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n908), .A2(KEYINPUT104), .A3(new_n913), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT105), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n916), .A2(new_n918), .A3(KEYINPUT105), .A4(new_n919), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n651), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n623), .A2(new_n638), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n900), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n699), .A2(G1), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n655), .A2(new_n927), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT45), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT106), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(KEYINPUT44), .C1(new_n655), .C2(new_n927), .ZN(new_n936));
  XOR2_X1   g0736(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n937));
  OR3_X1    g0737(.A1(new_n655), .A2(new_n927), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n939), .A2(KEYINPUT107), .A3(new_n925), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n925), .B1(new_n939), .B2(KEYINPUT107), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n650), .B(new_n652), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n644), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n696), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n658), .B(KEYINPUT41), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n931), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n922), .A2(new_n925), .A3(new_n927), .A4(new_n923), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n929), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n755), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n758), .B1(new_n231), .B2(new_n313), .C1(new_n243), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n398), .B1(new_n745), .B2(G97), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n954), .B1(new_n465), .B2(new_n717), .C1(new_n736), .C2(new_n730), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(G283), .B2(new_n778), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n737), .A2(new_n789), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n957), .A2(KEYINPUT46), .B1(new_n722), .B2(new_n726), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(KEYINPUT46), .B2(new_n957), .ZN(new_n959));
  AND2_X1   g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(G317), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n211), .B2(new_n723), .C1(new_n961), .C2(new_n713), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n730), .A2(new_n253), .B1(new_n723), .B2(new_n225), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n965));
  INV_X1    g0765(.A(G143), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n726), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT109), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n278), .B1(new_n735), .B2(new_n217), .C1(new_n220), .C2(new_n737), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n215), .B2(new_n721), .C1(new_n780), .C2(new_n713), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n717), .A2(new_n747), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n962), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT110), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT47), .Z(new_n977));
  OAI211_X1 g0777(.A(new_n701), .B(new_n953), .C1(new_n977), .C2(new_n710), .ZN(new_n978));
  INV_X1    g0778(.A(new_n911), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n978), .B1(new_n706), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n951), .A2(new_n981), .ZN(G387));
  NAND2_X1  g0782(.A1(new_n696), .A2(new_n944), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n659), .B1(new_n983), .B2(KEYINPUT111), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n696), .A2(new_n944), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n984), .B(new_n986), .C1(KEYINPUT111), .C2(new_n983), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n945), .A2(new_n930), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n952), .B1(new_n240), .B2(G45), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n660), .A2(new_n277), .A3(new_n657), .ZN(new_n990));
  INV_X1    g0790(.A(new_n660), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n257), .A2(G50), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT50), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n467), .C1(new_n225), .C2(new_n217), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n989), .A2(new_n990), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n657), .A2(new_n211), .ZN(new_n996));
  AOI211_X1 g0796(.A(new_n709), .B(new_n706), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G322), .A2(new_n727), .B1(new_n742), .B2(G311), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n736), .B2(new_n721), .C1(new_n961), .C2(new_n730), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n733), .B2(new_n723), .C1(new_n465), .C2(new_n737), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT49), .Z(new_n1002));
  INV_X1    g0802(.A(G326), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n391), .B1(new_n789), .B2(new_n735), .C1(new_n1003), .C2(new_n713), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n727), .A2(G159), .B1(new_n778), .B2(G68), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n785), .A2(G77), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n313), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n795), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1006), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n713), .A2(new_n253), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n398), .B1(new_n215), .B2(new_n730), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n717), .A2(new_n257), .B1(new_n735), .B2(new_n207), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n709), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n701), .C1(new_n650), .C2(new_n707), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n987), .B(new_n988), .C1(new_n997), .C2(new_n1016), .ZN(G393));
  OR2_X1    g0817(.A1(new_n939), .A2(new_n925), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n939), .A2(new_n925), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(new_n931), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n758), .B1(new_n207), .B2(new_n231), .C1(new_n250), .C2(new_n952), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n742), .A2(G50), .B1(new_n795), .B2(G77), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n257), .B2(new_n721), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n735), .A2(new_n205), .B1(new_n713), .B2(new_n966), .ZN(new_n1025));
  NOR3_X1   g0825(.A1(new_n1024), .A2(new_n391), .A3(new_n1025), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n726), .A2(new_n253), .B1(new_n730), .B2(new_n747), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT51), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(new_n225), .C2(new_n737), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G283), .A2(new_n785), .B1(new_n714), .B2(G322), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT112), .Z(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n211), .B2(new_n735), .C1(new_n736), .C2(new_n717), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n726), .A2(new_n961), .B1(new_n730), .B2(new_n722), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT52), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n278), .B1(new_n778), .B2(G294), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n789), .C2(new_n723), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1029), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT113), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n709), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n900), .A2(new_n706), .A3(new_n926), .ZN(new_n1040));
  AND3_X1   g0840(.A1(new_n1039), .A2(new_n1040), .A3(new_n701), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1021), .B1(new_n1022), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n942), .A2(new_n985), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1020), .A2(new_n986), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1043), .A2(new_n658), .A3(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1042), .A2(new_n1045), .ZN(G390));
  NAND2_X1  g0846(.A1(new_n764), .A2(new_n344), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n669), .A2(new_n670), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n772), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n844), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n886), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n1051), .A3(new_n838), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT114), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n885), .A2(new_n887), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n882), .B2(new_n886), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1050), .A2(new_n838), .A3(KEYINPUT114), .A4(new_n1051), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  AND4_X1   g0858(.A1(G330), .A2(new_n694), .A3(new_n765), .A4(new_n844), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(KEYINPUT115), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1054), .A2(new_n1056), .A3(new_n1060), .A4(new_n1057), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n694), .A2(G330), .A3(new_n765), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n881), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n774), .B1(new_n843), .B2(new_n839), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n870), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(KEYINPUT116), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n767), .A2(new_n772), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT116), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1065), .A2(new_n1071), .A3(new_n881), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1065), .A2(new_n881), .B1(new_n870), .B2(new_n1067), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n772), .A3(new_n1048), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n871), .B(new_n614), .C1(new_n676), .C2(new_n443), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1064), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1077), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1062), .A2(new_n1081), .A3(new_n1063), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n658), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1062), .A2(new_n930), .A3(new_n1063), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT117), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1055), .A2(new_n704), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n776), .A2(new_n257), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT54), .B(G143), .Z(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n721), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n785), .A2(G150), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT53), .ZN(new_n1092));
  INV_X1    g0892(.A(G132), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n278), .B1(new_n730), .B2(new_n1093), .C1(new_n780), .C2(new_n717), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(G50), .A2(new_n745), .B1(new_n714), .B2(G125), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1095), .B(new_n1096), .C1(new_n747), .C2(new_n723), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1090), .B(new_n1097), .C1(G128), .C2(new_n727), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n783), .B(new_n739), .C1(G107), .C2(new_n742), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n778), .A2(G97), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n278), .B1(new_n795), .B2(G77), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n727), .A2(G283), .B1(new_n714), .B2(G294), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G116), .B2(new_n731), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n709), .B1(new_n1098), .B2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1086), .A2(new_n701), .A3(new_n1087), .A4(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1084), .A2(new_n1085), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1085), .B1(new_n1084), .B2(new_n1106), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1083), .B1(new_n1107), .B2(new_n1108), .ZN(G378));
  XOR2_X1   g0909(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1110));
  XNOR2_X1  g0910(.A(new_n379), .B(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n267), .A2(new_n814), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n878), .B2(G330), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n861), .A2(new_n1113), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n889), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1082), .B2(new_n1078), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n878), .A2(G330), .A3(new_n1114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n861), .A2(new_n1113), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n888), .A4(new_n883), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1124), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1120), .A2(new_n1126), .A3(new_n1121), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1125), .A2(new_n1127), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n658), .B(new_n1123), .C1(new_n1128), .C2(KEYINPUT57), .ZN(new_n1129));
  AOI21_X1  g0929(.A(G41), .B1(new_n398), .B2(G33), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1130), .A2(G50), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G41), .B1(new_n714), .B2(G124), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n721), .A2(new_n780), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n1089), .A2(new_n737), .B1(new_n253), .B2(new_n723), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G128), .C2(new_n731), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n727), .A2(G125), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n1093), .C2(new_n717), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n273), .B(new_n1132), .C1(new_n1137), .C2(KEYINPUT59), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G159), .B2(new_n745), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(KEYINPUT59), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1131), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g0941(.A(G41), .B1(new_n727), .B2(G116), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1142), .A2(new_n391), .A3(new_n1007), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n735), .A2(new_n220), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(G283), .B2(new_n714), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n225), .B2(new_n723), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1143), .B(new_n1146), .C1(new_n1008), .C2(new_n778), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(new_n207), .B2(new_n717), .C1(new_n211), .C2(new_n730), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT58), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n710), .B1(new_n1141), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n700), .B1(new_n215), .B2(new_n776), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n1150), .B(new_n1153), .C1(new_n1114), .C2(new_n704), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1155), .B2(new_n930), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1129), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(G375));
  OAI21_X1  g0958(.A(new_n1009), .B1(new_n465), .B2(new_n726), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n713), .A2(new_n736), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n217), .A2(new_n735), .B1(new_n721), .B2(new_n211), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n277), .B1(new_n737), .B2(new_n207), .ZN(new_n1162));
  NOR4_X1   g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n789), .B2(new_n717), .C1(new_n733), .C2(new_n730), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n723), .A2(new_n215), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n726), .A2(new_n1093), .B1(new_n737), .B2(new_n747), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G150), .C2(new_n778), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n714), .A2(G128), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n742), .A2(new_n1088), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n391), .B(new_n1144), .C1(G137), .C2(new_n731), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n710), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n700), .B(new_n1172), .C1(new_n225), .C2(new_n776), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n844), .A2(new_n705), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT120), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1076), .A2(new_n930), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1073), .A2(new_n1077), .A3(new_n1075), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n947), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1178), .B2(new_n1081), .ZN(G381));
  AND2_X1   g0979(.A1(new_n1084), .A2(new_n1106), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1083), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1157), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(G390), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n951), .A2(new_n1184), .A3(new_n981), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1186));
  XOR2_X1   g0986(.A(new_n1186), .B(KEYINPUT121), .Z(new_n1187));
  OR4_X1    g0987(.A1(G381), .A2(new_n1183), .A3(new_n1185), .A4(new_n1187), .ZN(G407));
  OAI211_X1 g0988(.A(G407), .B(G213), .C1(G343), .C2(new_n1183), .ZN(G409));
  NAND2_X1  g0989(.A1(new_n1082), .A2(new_n1078), .ZN(new_n1190));
  AOI21_X1  g0990(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1123), .A2(new_n658), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G378), .B(new_n1156), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1120), .A2(new_n1126), .A3(new_n1121), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1126), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n947), .B(new_n1190), .C1(new_n1194), .C2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1154), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1117), .A2(new_n930), .A3(new_n1122), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n1182), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1193), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n637), .A2(G213), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G384), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT60), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1177), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  AND3_X1   g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1079), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1207), .B1(new_n1206), .B2(new_n1079), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n658), .B1(new_n1177), .B2(new_n1205), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1176), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n844), .B1(new_n870), .B2(new_n765), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1214), .A2(new_n1059), .A3(new_n1049), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n762), .B1(new_n675), .B2(new_n765), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1074), .B2(KEYINPUT116), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1215), .B1(new_n1217), .B2(new_n1072), .ZN(new_n1218));
  AOI21_X1  g1018(.A(KEYINPUT60), .B1(new_n1218), .B2(new_n1077), .ZN(new_n1219));
  OAI21_X1  g1019(.A(KEYINPUT122), .B1(new_n1219), .B2(new_n1081), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1210), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1206), .A2(new_n1207), .A3(new_n1079), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(G384), .A3(new_n1176), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1213), .A2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n637), .A2(G213), .A3(G2897), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(KEYINPUT125), .B1(new_n1225), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1229), .B(new_n1226), .C1(new_n1213), .C2(new_n1224), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT123), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1223), .A2(G384), .A3(new_n1176), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1223), .B2(new_n1176), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1213), .A2(KEYINPUT123), .A3(new_n1224), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1226), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1235), .A2(new_n1236), .A3(KEYINPUT124), .A4(new_n1226), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1203), .A2(new_n1231), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1233), .A2(new_n1234), .A3(new_n1232), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT123), .B1(new_n1213), .B2(new_n1224), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1201), .A2(new_n1244), .A3(new_n1202), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1201), .A2(new_n1244), .A3(new_n1248), .A4(new_n1202), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1241), .A2(new_n1246), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  XOR2_X1   g1050(.A(G393), .B(G396), .Z(new_n1251));
  NAND2_X1  g1051(.A1(new_n1185), .A2(KEYINPUT126), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1184), .B1(new_n951), .B2(new_n981), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G387), .A2(G390), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1251), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1255), .A2(new_n1256), .A3(KEYINPUT126), .A4(new_n1185), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT63), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1258), .B1(new_n1260), .B2(new_n1245), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1201), .A2(new_n1244), .A3(KEYINPUT63), .A4(new_n1202), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1261), .A2(new_n1247), .A3(new_n1241), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1259), .A2(new_n1263), .ZN(G405));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1265), .B(new_n1193), .C1(new_n1157), .C2(new_n1181), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1193), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1181), .B1(new_n1129), .B2(new_n1156), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT127), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1269), .A3(new_n1244), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1193), .B(new_n1225), .C1(new_n1157), .C2(new_n1181), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1258), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1270), .A2(new_n1257), .A3(new_n1254), .A4(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(G402));
endmodule


