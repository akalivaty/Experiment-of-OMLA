//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT66), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n465), .A2(new_n467), .A3(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n465), .A2(new_n467), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n475), .A2(new_n463), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n475), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  OR2_X1    g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n480), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n464), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G102), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G126), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n486), .B1(new_n490), .B2(new_n463), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n463), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n489), .A2(KEYINPUT4), .A3(G138), .A4(new_n463), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n484), .B1(new_n491), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n486), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n487), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n498), .B1(new_n500), .B2(G2105), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(KEYINPUT68), .A3(new_n494), .A4(new_n495), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n497), .A2(new_n502), .ZN(G164));
  AND2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .A3(G50), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g090(.A(KEYINPUT5), .B(G543), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g098(.A(KEYINPUT70), .B1(new_n523), .B2(new_n506), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n511), .A3(new_n525), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT71), .B(G88), .Z(new_n527));
  NAND3_X1  g102(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n515), .A2(new_n519), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND2_X1   g105(.A1(new_n524), .A2(new_n526), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n508), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n532), .A2(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  AOI22_X1  g114(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n541), .A2(G651), .B1(new_n508), .B2(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n524), .A2(new_n526), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  NAND2_X1  g121(.A1(new_n531), .A2(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n523), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n550), .A2(G651), .B1(new_n508), .B2(G43), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n508), .A2(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n560), .B2(KEYINPUT73), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n508), .A2(KEYINPUT72), .A3(G53), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(KEYINPUT9), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n531), .A2(G91), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n559), .B(new_n565), .C1(new_n560), .C2(KEYINPUT73), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n518), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n563), .A2(new_n564), .A3(new_n566), .A4(new_n568), .ZN(G299));
  OAI21_X1  g144(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n508), .A2(G49), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n570), .B(new_n571), .C1(new_n544), .C2(new_n572), .ZN(G288));
  NAND3_X1  g148(.A1(new_n524), .A2(G86), .A3(new_n526), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n508), .A2(G48), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n520), .A2(new_n522), .A3(G61), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n516), .A2(KEYINPUT74), .A3(G61), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n576), .A2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n508), .A2(G47), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  OAI221_X1 g162(.A(new_n585), .B1(new_n518), .B2(new_n586), .C1(new_n544), .C2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  OR3_X1    g164(.A1(G171), .A2(KEYINPUT75), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT75), .B1(G171), .B2(new_n589), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OR3_X1    g167(.A1(new_n544), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n523), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(new_n508), .B2(G54), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT10), .B1(new_n544), .B2(new_n592), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n590), .B(new_n591), .C1(G868), .C2(new_n600), .ZN(G284));
  OAI211_X1 g176(.A(new_n590), .B(new_n591), .C1(G868), .C2(new_n600), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  XNOR2_X1  g181(.A(KEYINPUT76), .B(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(G860), .B2(new_n607), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n552), .ZN(G323));
  XOR2_X1   g186(.A(G323), .B(KEYINPUT77), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n489), .A2(new_n485), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2100), .ZN(new_n617));
  INV_X1    g192(.A(new_n476), .ZN(new_n618));
  INV_X1    g193(.A(G123), .ZN(new_n619));
  OR3_X1    g194(.A1(new_n618), .A2(KEYINPUT78), .A3(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT78), .B1(new_n618), .B2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n478), .A2(G135), .ZN(new_n622));
  OR2_X1    g197(.A1(G99), .A2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n624));
  NAND4_X1  g199(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n625), .A2(G2096), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(G2096), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n617), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT79), .Z(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2443), .B(G2446), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT80), .ZN(G401));
  INV_X1    g218(.A(KEYINPUT18), .ZN(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(G2096), .Z(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  AOI21_X1  g228(.A(new_n653), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT81), .B(G2100), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G227));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT82), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  AND2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n665), .A2(new_n666), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n662), .A2(new_n667), .A3(new_n664), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n668), .B(new_n669), .C1(new_n666), .C2(new_n665), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(G1986), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G1991), .B(G1996), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G1981), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G229));
  INV_X1    g252(.A(G1971), .ZN(new_n678));
  NAND2_X1  g253(.A1(G166), .A2(G16), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n680));
  OR2_X1    g255(.A1(G16), .A2(G22), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n680), .B1(new_n679), .B2(new_n681), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n678), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n679), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(KEYINPUT85), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(G1971), .A3(new_n682), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(G6), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G305), .B2(G16), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT32), .B(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n685), .A2(new_n688), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n689), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n689), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT33), .ZN(new_n698));
  INV_X1    g273(.A(G1976), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n697), .A2(KEYINPUT33), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(KEYINPUT33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n701), .A2(G1976), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT34), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n689), .A2(G24), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G290), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n710), .A2(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(G1986), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT83), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G119), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n478), .A2(G131), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(G25), .B(new_n718), .S(G29), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT84), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT35), .B(G1991), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n707), .A2(new_n711), .A3(new_n712), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(KEYINPUT86), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n705), .A2(new_n706), .B1(G1986), .B2(new_n710), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT86), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n725), .A2(new_n726), .A3(new_n711), .A4(new_n722), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n705), .A2(new_n706), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n730), .B1(new_n724), .B2(new_n727), .ZN(new_n733));
  NAND2_X1  g308(.A1(KEYINPUT87), .A2(KEYINPUT36), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n732), .A2(KEYINPUT87), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G16), .A2(G19), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n552), .B2(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1341), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n689), .A2(KEYINPUT23), .A3(G20), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n740));
  INV_X1    g315(.A(G20), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n740), .B1(new_n741), .B2(G16), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n739), .B(new_n742), .C1(new_n604), .C2(new_n689), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  NOR2_X1   g319(.A1(G4), .A2(G16), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n600), .B2(G16), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n744), .B1(G1348), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G27), .A2(G29), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G164), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2078), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n485), .A2(G103), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT25), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n478), .A2(G139), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n759), .A2(new_n463), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(new_n751), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT91), .ZN(new_n763));
  INV_X1    g338(.A(G2072), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n750), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(G168), .A2(KEYINPUT93), .A3(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT93), .B1(G16), .B2(G21), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G286), .B2(new_n689), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT94), .ZN(new_n769));
  INV_X1    g344(.A(G1966), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  AND3_X1   g346(.A1(new_n766), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n769), .A2(new_n770), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  OR2_X1    g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  NAND2_X1  g351(.A1(KEYINPUT24), .A2(G34), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n776), .A2(new_n751), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G160), .B2(new_n751), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT92), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G2084), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n774), .A2(new_n775), .A3(new_n782), .ZN(new_n783));
  AND4_X1   g358(.A1(new_n738), .A2(new_n747), .A3(new_n765), .A4(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n625), .A2(new_n751), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n781), .A2(G2084), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G11), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n786), .B(new_n787), .C1(new_n763), .C2(new_n764), .ZN(new_n788));
  OAI21_X1  g363(.A(KEYINPUT96), .B1(G5), .B2(G16), .ZN(new_n789));
  OR3_X1    g364(.A1(KEYINPUT96), .A2(G5), .A3(G16), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n789), .B(new_n790), .C1(G301), .C2(new_n689), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1961), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n751), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n751), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT97), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT29), .ZN(new_n796));
  INV_X1    g371(.A(G2090), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT28), .ZN(new_n799));
  INV_X1    g374(.A(G26), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(G29), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(G29), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n478), .A2(G140), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n476), .A2(G128), .ZN(new_n806));
  OR2_X1    g381(.A1(G104), .A2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n478), .A2(KEYINPUT89), .A3(G140), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n805), .A2(new_n806), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n802), .B1(new_n810), .B2(G29), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n801), .B1(new_n811), .B2(new_n799), .ZN(new_n812));
  INV_X1    g387(.A(G2067), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT95), .B(G28), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT30), .ZN(new_n816));
  OAI221_X1 g391(.A(new_n814), .B1(G29), .B2(new_n816), .C1(G1348), .C2(new_n746), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n788), .A2(new_n798), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n796), .A2(new_n797), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n784), .A2(new_n785), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n737), .A2(G1341), .ZN(new_n821));
  NOR2_X1   g396(.A1(G29), .A2(G32), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n478), .A2(G141), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n476), .A2(G129), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n485), .A2(G105), .ZN(new_n825));
  NAND3_X1  g400(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT26), .Z(new_n827));
  NAND4_X1  g402(.A1(new_n823), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n822), .B1(new_n829), .B2(G29), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT27), .B(G1996), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n820), .A2(new_n821), .A3(new_n832), .ZN(new_n833));
  AOI211_X1 g408(.A(KEYINPUT88), .B(new_n730), .C1(new_n724), .C2(new_n727), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(KEYINPUT36), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n735), .A2(new_n835), .ZN(G311));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n732), .A2(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n733), .A2(new_n734), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT87), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n733), .B2(new_n729), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n838), .B(new_n833), .C1(new_n839), .C2(new_n841), .ZN(G150));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n531), .A2(G93), .ZN(new_n844));
  NAND2_X1  g419(.A1(G80), .A2(G543), .ZN(new_n845));
  INV_X1    g420(.A(G67), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n523), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n847), .A2(G651), .B1(new_n508), .B2(G55), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n547), .A2(new_n551), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n552), .A2(KEYINPUT100), .A3(new_n849), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g429(.A(KEYINPUT101), .B1(new_n552), .B2(new_n849), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n850), .A2(new_n856), .A3(new_n851), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n600), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT99), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n861), .B(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(KEYINPUT102), .Z(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n864), .B2(KEYINPUT39), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n849), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(new_n718), .B(new_n615), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n478), .A2(G142), .ZN(new_n873));
  NOR2_X1   g448(.A1(G106), .A2(G2105), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n876), .B1(G130), .B2(new_n476), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n872), .B(new_n877), .Z(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT103), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n500), .A2(G2105), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n881), .A2(new_n486), .A3(new_n494), .A4(new_n495), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n761), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n810), .B(new_n828), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n879), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n625), .B(G160), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(G162), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n878), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n886), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(new_n849), .A2(new_n589), .ZN(new_n898));
  XNOR2_X1  g473(.A(G305), .B(G288), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(G290), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G303), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT42), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n604), .A2(new_n600), .ZN(new_n903));
  NOR2_X1   g478(.A1(G299), .A2(new_n599), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n903), .A2(new_n904), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT41), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n859), .B(new_n609), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n913), .B1(new_n912), .B2(new_n905), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n902), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n898), .B1(new_n915), .B2(new_n589), .ZN(G295));
  OAI21_X1  g491(.A(new_n898), .B1(new_n915), .B2(new_n589), .ZN(G331));
  NAND3_X1  g492(.A1(new_n854), .A2(new_n858), .A3(G301), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(G301), .B1(new_n854), .B2(new_n858), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n919), .A2(G286), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n859), .A2(G171), .ZN(new_n922));
  AOI21_X1  g497(.A(G168), .B1(new_n922), .B2(new_n918), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n911), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(G286), .B1(new_n919), .B2(new_n920), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(G168), .A3(new_n918), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n908), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n901), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n924), .A2(new_n901), .A3(new_n927), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n905), .A2(new_n909), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n908), .A2(new_n906), .ZN(new_n938));
  OAI211_X1 g513(.A(new_n937), .B(new_n938), .C1(new_n921), .C2(new_n923), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n925), .A2(new_n926), .A3(KEYINPUT105), .A4(new_n908), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n929), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n932), .A2(new_n931), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n934), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n933), .A2(new_n944), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n948), .B1(new_n947), .B2(new_n951), .ZN(G397));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n953));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n491), .B2(new_n496), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n957));
  NOR2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(KEYINPUT107), .B1(G160), .B2(G40), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n468), .A2(new_n469), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G2105), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n471), .A2(new_n472), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n463), .ZN(new_n964));
  AND4_X1   g539(.A1(KEYINPUT107), .A2(new_n962), .A3(new_n964), .A4(G40), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n960), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n953), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n962), .A2(new_n964), .A3(G40), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(G160), .A2(KEYINPUT107), .A3(G40), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n958), .A2(KEYINPUT108), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n967), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(G1996), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  INV_X1    g551(.A(new_n974), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n810), .B(G2067), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n976), .A2(new_n829), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n718), .A2(new_n721), .ZN(new_n980));
  AND2_X1   g555(.A1(new_n718), .A2(new_n721), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(G1996), .A3(new_n828), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT110), .ZN(new_n984));
  XNOR2_X1  g559(.A(G290), .B(G1986), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n979), .A2(new_n982), .A3(new_n984), .A4(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n987), .B(KEYINPUT111), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n955), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT112), .B(new_n954), .C1(new_n491), .C2(new_n496), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n497), .A2(new_n502), .A3(new_n954), .A4(new_n957), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n972), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n770), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n990), .A2(new_n992), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n966), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G2084), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT113), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n497), .A2(new_n502), .A3(new_n954), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n1004), .B2(KEYINPUT50), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1004), .A2(new_n1003), .A3(KEYINPUT50), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1001), .B(new_n1002), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n995), .A2(KEYINPUT117), .A3(new_n770), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n998), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1009), .A2(G8), .A3(G168), .ZN(new_n1010));
  INV_X1    g585(.A(new_n992), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT112), .B1(new_n882), .B2(new_n954), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n972), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n972), .A2(new_n1000), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1013), .A2(KEYINPUT116), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n972), .C1(new_n999), .C2(new_n1000), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1015), .A2(new_n1017), .A3(new_n797), .A4(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n957), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1004), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n956), .A2(KEYINPUT45), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n972), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(new_n678), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G8), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  NAND3_X1  g602(.A1(G303), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1027), .B1(G303), .B2(G8), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1026), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n999), .B2(new_n972), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n696), .A2(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(G288), .B2(new_n699), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n583), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n574), .A2(new_n575), .ZN(new_n1042));
  OAI21_X1  g617(.A(G1981), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1981), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n576), .A2(new_n1044), .A3(new_n583), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1043), .A2(new_n1045), .A3(KEYINPUT49), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT49), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1044), .B1(new_n576), .B2(new_n583), .ZN(new_n1048));
  AND4_X1   g623(.A1(new_n1044), .A2(new_n583), .A3(new_n574), .A4(new_n575), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1036), .A2(new_n1046), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT115), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1036), .A2(new_n1053), .A3(new_n1050), .A4(new_n1046), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1038), .B(new_n1040), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1001), .B(new_n797), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1024), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT114), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1030), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1028), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1010), .A2(new_n1033), .A3(new_n1055), .A4(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT118), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1038), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1040), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1063), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1069), .A2(new_n1070), .A3(new_n1033), .A4(new_n1010), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT63), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1065), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1038), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1067), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1031), .B1(new_n1057), .B2(G8), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1072), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT119), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1063), .A3(new_n1010), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1073), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1076), .A2(new_n1063), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1074), .A2(new_n699), .A3(new_n696), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1045), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n1086), .B2(new_n1036), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT122), .B(G1961), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G2078), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n993), .A2(new_n972), .A3(new_n994), .A4(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1092), .B1(new_n1023), .B2(G2078), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(G171), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n998), .A2(G168), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(G8), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1009), .B2(G286), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1103), .B2(KEYINPUT62), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1031), .B1(new_n1025), .B2(G8), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT125), .B1(new_n1068), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT125), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1033), .A2(new_n1055), .A3(new_n1107), .A4(new_n1063), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1100), .B(new_n1110), .C1(new_n1099), .C2(new_n1102), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1104), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1083), .A2(new_n1087), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n1114));
  OAI21_X1  g689(.A(G2105), .B1(new_n961), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT124), .B1(new_n468), .B2(new_n469), .ZN(new_n1116));
  OAI211_X1 g691(.A(G40), .B(new_n964), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n959), .A2(new_n1022), .A3(new_n1093), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1004), .A2(KEYINPUT50), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT113), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1004), .A2(new_n1003), .A3(KEYINPUT50), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI211_X1 g698(.A(KEYINPUT123), .B(new_n1089), .C1(new_n1123), .C2(new_n1001), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1095), .B(new_n1119), .C1(new_n1124), .C2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1097), .B1(new_n1127), .B2(G171), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(G171), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT126), .B1(new_n1096), .B2(G171), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1133), .A2(new_n1134), .A3(G301), .A4(new_n1095), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1131), .A2(KEYINPUT54), .A3(new_n1132), .A4(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1109), .A2(new_n1130), .A3(new_n1136), .A4(new_n1103), .ZN(new_n1137));
  INV_X1    g712(.A(G1348), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1088), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n999), .A2(new_n813), .A3(new_n972), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n600), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  OR2_X1    g720(.A1(new_n1023), .A2(G1996), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n1013), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1145), .B1(new_n1149), .B2(new_n552), .ZN(new_n1150));
  AOI211_X1 g725(.A(KEYINPUT59), .B(new_n851), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1142), .A2(new_n599), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1141), .A2(new_n600), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1143), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT57), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G299), .B(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(KEYINPUT56), .B(G2072), .Z(new_n1159));
  OR2_X1    g734(.A1(new_n1023), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1161));
  INV_X1    g736(.A(G1956), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT120), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1158), .B(new_n1160), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT121), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1160), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1158), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT120), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1163), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1174), .A2(new_n1175), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1167), .A2(new_n1170), .A3(new_n1176), .A4(KEYINPUT61), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1166), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1158), .B1(new_n1174), .B2(new_n1160), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1178), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1156), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(new_n1154), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1183), .A2(new_n1180), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1137), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n988), .B1(new_n1113), .B2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n979), .A2(new_n982), .A3(new_n984), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n974), .A2(G1986), .A3(G290), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT48), .Z(new_n1191));
  NAND4_X1  g766(.A1(new_n979), .A2(KEYINPUT127), .A3(new_n982), .A4(new_n984), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n977), .B1(new_n828), .B2(new_n978), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n1196));
  AND3_X1   g771(.A1(new_n1195), .A2(KEYINPUT46), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g772(.A(KEYINPUT46), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1194), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1199), .A2(KEYINPUT47), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT47), .ZN(new_n1201));
  OAI211_X1 g776(.A(new_n1201), .B(new_n1194), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  AND3_X1   g778(.A1(new_n979), .A2(new_n980), .A3(new_n984), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n810), .A2(G2067), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n977), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AND3_X1   g781(.A1(new_n1193), .A2(new_n1203), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1186), .A2(new_n1207), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g783(.A1(new_n642), .A2(new_n657), .ZN(new_n1210));
  AOI21_X1  g784(.A(new_n1210), .B1(new_n892), .B2(new_n895), .ZN(new_n1211));
  NAND4_X1  g785(.A1(new_n946), .A2(new_n1211), .A3(G319), .A4(new_n676), .ZN(G225));
  INV_X1    g786(.A(G225), .ZN(G308));
endmodule


