

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G543), .A2(G651), .ZN(n547) );
  INV_X1 U555 ( .A(n920), .ZN(n990) );
  NAND2_X2 U556 ( .A1(n581), .A2(n580), .ZN(n987) );
  NOR2_X2 U557 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U558 ( .A(n746), .B(KEYINPUT32), .ZN(n754) );
  BUF_X1 U559 ( .A(n712), .Z(n738) );
  INV_X1 U560 ( .A(n712), .ZN(n689) );
  NAND2_X1 U561 ( .A1(n754), .A2(n753), .ZN(n768) );
  NOR2_X1 U562 ( .A1(n987), .A2(n717), .ZN(n719) );
  BUF_X1 U563 ( .A(n701), .Z(n709) );
  XNOR2_X1 U564 ( .A(n687), .B(n686), .ZN(n802) );
  NOR2_X1 U565 ( .A1(n544), .A2(n543), .ZN(n685) );
  BUF_X2 U566 ( .A(n537), .Z(n521) );
  NOR2_X1 U567 ( .A1(n706), .A2(n705), .ZN(n725) );
  XNOR2_X1 U568 ( .A(KEYINPUT30), .B(KEYINPUT99), .ZN(n696) );
  INV_X1 U569 ( .A(n994), .ZN(n760) );
  NAND2_X1 U570 ( .A1(n685), .A2(G40), .ZN(n687) );
  INV_X1 U571 ( .A(G2105), .ZN(n533) );
  BUF_X1 U572 ( .A(n685), .Z(G160) );
  XOR2_X1 U573 ( .A(n697), .B(n696), .Z(n520) );
  INV_X1 U574 ( .A(KEYINPUT26), .ZN(n713) );
  INV_X1 U575 ( .A(KEYINPUT64), .ZN(n718) );
  OR2_X1 U576 ( .A1(n990), .A2(n722), .ZN(n721) );
  NOR2_X1 U577 ( .A1(n725), .A2(n984), .ZN(n708) );
  NOR2_X1 U578 ( .A1(n759), .A2(G1966), .ZN(n750) );
  INV_X1 U579 ( .A(KEYINPUT90), .ZN(n686) );
  NOR2_X1 U580 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U581 ( .A1(n763), .A2(n762), .ZN(n767) );
  AND2_X1 U582 ( .A1(G2104), .A2(G101), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U584 ( .A(KEYINPUT104), .ZN(n783) );
  INV_X1 U585 ( .A(KEYINPUT89), .ZN(n525) );
  INV_X1 U586 ( .A(KEYINPUT17), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT15), .B(n595), .Z(n920) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U589 ( .A(KEYINPUT1), .B(n553), .Z(n650) );
  BUF_X1 U590 ( .A(n684), .Z(G164) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n533), .ZN(n537) );
  NAND2_X1 U592 ( .A1(G126), .A2(n521), .ZN(n522) );
  XNOR2_X1 U593 ( .A(n522), .B(KEYINPUT88), .ZN(n528) );
  NOR2_X2 U594 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  XNOR2_X2 U595 ( .A(n524), .B(n523), .ZN(n904) );
  NAND2_X1 U596 ( .A1(n904), .A2(G138), .ZN(n526) );
  NAND2_X1 U597 ( .A1(n528), .A2(n527), .ZN(n532) );
  AND2_X1 U598 ( .A1(n533), .A2(G2104), .ZN(n906) );
  NAND2_X1 U599 ( .A1(G102), .A2(n906), .ZN(n530) );
  AND2_X1 U600 ( .A1(G2104), .A2(G2105), .ZN(n901) );
  NAND2_X1 U601 ( .A1(G114), .A2(n901), .ZN(n529) );
  NAND2_X1 U602 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U603 ( .A1(n532), .A2(n531), .ZN(n684) );
  INV_X1 U604 ( .A(KEYINPUT23), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n537), .A2(G125), .ZN(n538) );
  NAND2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(KEYINPUT66), .B(n540), .ZN(n544) );
  NAND2_X1 U609 ( .A1(n904), .A2(G137), .ZN(n542) );
  NAND2_X1 U610 ( .A1(n901), .A2(G113), .ZN(n541) );
  NAND2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U612 ( .A(G651), .ZN(n552) );
  XOR2_X1 U613 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  OR2_X1 U614 ( .A1(n552), .A2(n628), .ZN(n545) );
  XNOR2_X2 U615 ( .A(KEYINPUT67), .B(n545), .ZN(n654) );
  NAND2_X1 U616 ( .A1(n654), .A2(G76), .ZN(n546) );
  XNOR2_X1 U617 ( .A(KEYINPUT76), .B(n546), .ZN(n550) );
  XOR2_X1 U618 ( .A(KEYINPUT65), .B(n547), .Z(n653) );
  NAND2_X1 U619 ( .A1(n653), .A2(G89), .ZN(n548) );
  XNOR2_X1 U620 ( .A(KEYINPUT4), .B(n548), .ZN(n549) );
  NAND2_X1 U621 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U622 ( .A(n551), .B(KEYINPUT5), .ZN(n559) );
  XNOR2_X1 U623 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n557) );
  NOR2_X1 U624 ( .A1(G651), .A2(n628), .ZN(n649) );
  NAND2_X1 U625 ( .A1(G51), .A2(n649), .ZN(n555) );
  NOR2_X1 U626 ( .A1(G543), .A2(n552), .ZN(n553) );
  NAND2_X1 U627 ( .A1(G63), .A2(n650), .ZN(n554) );
  NAND2_X1 U628 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U629 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U630 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U631 ( .A(KEYINPUT7), .B(n560), .ZN(G168) );
  XOR2_X1 U632 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U633 ( .A1(n650), .A2(G65), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G53), .A2(n649), .ZN(n562) );
  NAND2_X1 U635 ( .A1(G78), .A2(n654), .ZN(n561) );
  NAND2_X1 U636 ( .A1(n562), .A2(n561), .ZN(n565) );
  NAND2_X1 U637 ( .A1(n653), .A2(G91), .ZN(n563) );
  XOR2_X1 U638 ( .A(KEYINPUT70), .B(n563), .Z(n564) );
  NOR2_X1 U639 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U640 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U641 ( .A(KEYINPUT71), .B(n568), .Z(G299) );
  XNOR2_X1 U642 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  AND2_X1 U643 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U644 ( .A(G132), .ZN(G219) );
  NAND2_X1 U645 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U646 ( .A(n569), .B(KEYINPUT10), .ZN(n570) );
  XNOR2_X1 U647 ( .A(KEYINPUT74), .B(n570), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n837) );
  NAND2_X1 U649 ( .A1(n837), .A2(G567), .ZN(n571) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U651 ( .A1(n653), .A2(G81), .ZN(n572) );
  XNOR2_X1 U652 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U653 ( .A1(G68), .A2(n654), .ZN(n573) );
  NAND2_X1 U654 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U655 ( .A(KEYINPUT13), .B(n575), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G43), .A2(n649), .ZN(n576) );
  XNOR2_X1 U657 ( .A(n576), .B(KEYINPUT75), .ZN(n579) );
  NAND2_X1 U658 ( .A1(G56), .A2(n650), .ZN(n577) );
  XOR2_X1 U659 ( .A(KEYINPUT14), .B(n577), .Z(n578) );
  INV_X1 U660 ( .A(G860), .ZN(n601) );
  OR2_X1 U661 ( .A1(n987), .A2(n601), .ZN(G153) );
  NAND2_X1 U662 ( .A1(G90), .A2(n653), .ZN(n583) );
  NAND2_X1 U663 ( .A1(G77), .A2(n654), .ZN(n582) );
  NAND2_X1 U664 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U665 ( .A(KEYINPUT9), .B(n584), .ZN(n588) );
  NAND2_X1 U666 ( .A1(G52), .A2(n649), .ZN(n586) );
  NAND2_X1 U667 ( .A1(G64), .A2(n650), .ZN(n585) );
  AND2_X1 U668 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U669 ( .A1(n588), .A2(n587), .ZN(G301) );
  NAND2_X1 U670 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G92), .A2(n653), .ZN(n590) );
  NAND2_X1 U672 ( .A1(G79), .A2(n654), .ZN(n589) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n594) );
  NAND2_X1 U674 ( .A1(G54), .A2(n649), .ZN(n592) );
  NAND2_X1 U675 ( .A1(G66), .A2(n650), .ZN(n591) );
  NAND2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n593) );
  NOR2_X1 U677 ( .A1(n594), .A2(n593), .ZN(n595) );
  INV_X1 U678 ( .A(G868), .ZN(n667) );
  NAND2_X1 U679 ( .A1(n990), .A2(n667), .ZN(n596) );
  NAND2_X1 U680 ( .A1(n597), .A2(n596), .ZN(G284) );
  NOR2_X1 U681 ( .A1(G286), .A2(n667), .ZN(n599) );
  NOR2_X1 U682 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U683 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U684 ( .A(KEYINPUT78), .B(n600), .ZN(G297) );
  NAND2_X1 U685 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U686 ( .A1(n602), .A2(n920), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n603), .B(KEYINPUT79), .ZN(n604) );
  XOR2_X1 U688 ( .A(KEYINPUT16), .B(n604), .Z(G148) );
  NOR2_X1 U689 ( .A1(G868), .A2(n987), .ZN(n607) );
  NAND2_X1 U690 ( .A1(G868), .A2(n920), .ZN(n605) );
  NOR2_X1 U691 ( .A1(G559), .A2(n605), .ZN(n606) );
  NOR2_X1 U692 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U693 ( .A1(G99), .A2(n906), .ZN(n609) );
  NAND2_X1 U694 ( .A1(G111), .A2(n901), .ZN(n608) );
  NAND2_X1 U695 ( .A1(n609), .A2(n608), .ZN(n615) );
  NAND2_X1 U696 ( .A1(G123), .A2(n521), .ZN(n610) );
  XNOR2_X1 U697 ( .A(n610), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U698 ( .A1(G135), .A2(n904), .ZN(n611) );
  XNOR2_X1 U699 ( .A(n611), .B(KEYINPUT80), .ZN(n612) );
  NAND2_X1 U700 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n938) );
  XNOR2_X1 U702 ( .A(n938), .B(G2096), .ZN(n617) );
  INV_X1 U703 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U704 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U705 ( .A1(G88), .A2(n653), .ZN(n619) );
  NAND2_X1 U706 ( .A1(G75), .A2(n654), .ZN(n618) );
  NAND2_X1 U707 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U708 ( .A1(n649), .A2(G50), .ZN(n620) );
  XOR2_X1 U709 ( .A(KEYINPUT82), .B(n620), .Z(n621) );
  NOR2_X1 U710 ( .A1(n622), .A2(n621), .ZN(n624) );
  NAND2_X1 U711 ( .A1(n650), .A2(G62), .ZN(n623) );
  NAND2_X1 U712 ( .A1(n624), .A2(n623), .ZN(G303) );
  INV_X1 U713 ( .A(G303), .ZN(G166) );
  NAND2_X1 U714 ( .A1(G49), .A2(n649), .ZN(n626) );
  NAND2_X1 U715 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U716 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U717 ( .A1(n650), .A2(n627), .ZN(n630) );
  NAND2_X1 U718 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U719 ( .A1(n630), .A2(n629), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G48), .A2(n649), .ZN(n632) );
  NAND2_X1 U721 ( .A1(G86), .A2(n653), .ZN(n631) );
  NAND2_X1 U722 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U723 ( .A1(n654), .A2(G73), .ZN(n633) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n633), .Z(n634) );
  NOR2_X1 U725 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U726 ( .A1(n650), .A2(G61), .ZN(n636) );
  NAND2_X1 U727 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U728 ( .A1(n654), .A2(G72), .ZN(n639) );
  NAND2_X1 U729 ( .A1(n653), .A2(G85), .ZN(n638) );
  NAND2_X1 U730 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U731 ( .A1(G47), .A2(n649), .ZN(n640) );
  XOR2_X1 U732 ( .A(KEYINPUT68), .B(n640), .Z(n641) );
  NOR2_X1 U733 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U734 ( .A1(n650), .A2(G60), .ZN(n643) );
  NAND2_X1 U735 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U736 ( .A(KEYINPUT69), .B(n645), .Z(G290) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n647) );
  XNOR2_X1 U738 ( .A(G288), .B(KEYINPUT83), .ZN(n646) );
  XNOR2_X1 U739 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U740 ( .A(G166), .B(n648), .ZN(n662) );
  INV_X1 U741 ( .A(G299), .ZN(n984) );
  XNOR2_X1 U742 ( .A(n984), .B(G305), .ZN(n660) );
  NAND2_X1 U743 ( .A1(G55), .A2(n649), .ZN(n652) );
  NAND2_X1 U744 ( .A1(G67), .A2(n650), .ZN(n651) );
  NAND2_X1 U745 ( .A1(n652), .A2(n651), .ZN(n658) );
  NAND2_X1 U746 ( .A1(G93), .A2(n653), .ZN(n656) );
  NAND2_X1 U747 ( .A1(G80), .A2(n654), .ZN(n655) );
  NAND2_X1 U748 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U749 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U750 ( .A(n659), .B(KEYINPUT81), .ZN(n846) );
  XNOR2_X1 U751 ( .A(n660), .B(n846), .ZN(n661) );
  XNOR2_X1 U752 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U753 ( .A(n663), .B(G290), .ZN(n919) );
  NAND2_X1 U754 ( .A1(G559), .A2(n920), .ZN(n664) );
  XNOR2_X1 U755 ( .A(n664), .B(n987), .ZN(n844) );
  XNOR2_X1 U756 ( .A(n919), .B(n844), .ZN(n665) );
  NAND2_X1 U757 ( .A1(n665), .A2(G868), .ZN(n666) );
  XOR2_X1 U758 ( .A(KEYINPUT85), .B(n666), .Z(n669) );
  NAND2_X1 U759 ( .A1(n846), .A2(n667), .ZN(n668) );
  NAND2_X1 U760 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U761 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XOR2_X1 U762 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U763 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U764 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U765 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XOR2_X1 U766 ( .A(KEYINPUT72), .B(G57), .Z(G237) );
  XNOR2_X1 U767 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NAND2_X1 U768 ( .A1(G108), .A2(G120), .ZN(n674) );
  NOR2_X1 U769 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U770 ( .A1(G69), .A2(n675), .ZN(n841) );
  NAND2_X1 U771 ( .A1(G567), .A2(n841), .ZN(n676) );
  XNOR2_X1 U772 ( .A(n676), .B(KEYINPUT87), .ZN(n682) );
  NOR2_X1 U773 ( .A1(G219), .A2(G220), .ZN(n678) );
  XNOR2_X1 U774 ( .A(KEYINPUT86), .B(KEYINPUT22), .ZN(n677) );
  XNOR2_X1 U775 ( .A(n678), .B(n677), .ZN(n679) );
  NAND2_X1 U776 ( .A1(n679), .A2(G96), .ZN(n680) );
  OR2_X1 U777 ( .A1(G218), .A2(n680), .ZN(n842) );
  AND2_X1 U778 ( .A1(G2106), .A2(n842), .ZN(n681) );
  NOR2_X1 U779 ( .A1(n682), .A2(n681), .ZN(G319) );
  INV_X1 U780 ( .A(G319), .ZN(n925) );
  NAND2_X1 U781 ( .A1(G483), .A2(G661), .ZN(n683) );
  NOR2_X1 U782 ( .A1(n925), .A2(n683), .ZN(n840) );
  NAND2_X1 U783 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U784 ( .A(G301), .ZN(G171) );
  NOR2_X1 U785 ( .A1(n684), .A2(G1384), .ZN(n803) );
  NAND2_X1 U786 ( .A1(n803), .A2(n802), .ZN(n712) );
  NOR2_X1 U787 ( .A1(n689), .A2(G1961), .ZN(n688) );
  XNOR2_X1 U788 ( .A(n688), .B(KEYINPUT95), .ZN(n691) );
  XNOR2_X1 U789 ( .A(n689), .B(KEYINPUT96), .ZN(n701) );
  XNOR2_X1 U790 ( .A(KEYINPUT25), .B(G2078), .ZN(n964) );
  NAND2_X1 U791 ( .A1(n709), .A2(n964), .ZN(n690) );
  NAND2_X1 U792 ( .A1(n691), .A2(n690), .ZN(n731) );
  NOR2_X1 U793 ( .A1(G171), .A2(n731), .ZN(n692) );
  XNOR2_X1 U794 ( .A(n692), .B(KEYINPUT100), .ZN(n699) );
  AND2_X1 U795 ( .A1(G8), .A2(n738), .ZN(n694) );
  INV_X1 U796 ( .A(KEYINPUT94), .ZN(n693) );
  XNOR2_X2 U797 ( .A(n694), .B(n693), .ZN(n759) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n738), .ZN(n747) );
  NOR2_X1 U799 ( .A1(n750), .A2(n747), .ZN(n695) );
  NAND2_X1 U800 ( .A1(G8), .A2(n695), .ZN(n697) );
  NOR2_X1 U801 ( .A1(G168), .A2(n520), .ZN(n698) );
  NOR2_X1 U802 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U803 ( .A(KEYINPUT31), .B(n700), .ZN(n736) );
  NAND2_X1 U804 ( .A1(n701), .A2(G2072), .ZN(n703) );
  XOR2_X1 U805 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n702) );
  XNOR2_X1 U806 ( .A(n703), .B(n702), .ZN(n706) );
  INV_X1 U807 ( .A(G1956), .ZN(n704) );
  NOR2_X1 U808 ( .A1(n709), .A2(n704), .ZN(n705) );
  INV_X1 U809 ( .A(KEYINPUT28), .ZN(n707) );
  XNOR2_X1 U810 ( .A(n708), .B(n707), .ZN(n729) );
  NAND2_X1 U811 ( .A1(n709), .A2(G2067), .ZN(n711) );
  NAND2_X1 U812 ( .A1(n738), .A2(G1348), .ZN(n710) );
  NAND2_X1 U813 ( .A1(n711), .A2(n710), .ZN(n722) );
  INV_X1 U814 ( .A(G1996), .ZN(n965) );
  NOR2_X1 U815 ( .A1(n712), .A2(n965), .ZN(n714) );
  XNOR2_X1 U816 ( .A(n714), .B(n713), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n738), .A2(G1341), .ZN(n715) );
  NAND2_X1 U818 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U819 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U820 ( .A1(n721), .A2(n720), .ZN(n724) );
  NAND2_X1 U821 ( .A1(n990), .A2(n722), .ZN(n723) );
  NAND2_X1 U822 ( .A1(n724), .A2(n723), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n984), .A2(n725), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U825 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U826 ( .A(n730), .B(KEYINPUT29), .ZN(n733) );
  AND2_X1 U827 ( .A1(G171), .A2(n731), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U829 ( .A(n734), .B(KEYINPUT98), .ZN(n735) );
  NOR2_X1 U830 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U831 ( .A(n737), .B(KEYINPUT101), .ZN(n748) );
  NAND2_X1 U832 ( .A1(n748), .A2(G286), .ZN(n743) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n738), .ZN(n740) );
  NOR2_X1 U834 ( .A1(n759), .A2(G1971), .ZN(n739) );
  NOR2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U836 ( .A1(n741), .A2(G303), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U838 ( .A(n744), .B(KEYINPUT102), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n745), .A2(G8), .ZN(n746) );
  NAND2_X1 U840 ( .A1(G8), .A2(n747), .ZN(n752) );
  INV_X1 U841 ( .A(n748), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U844 ( .A1(G1976), .A2(G288), .ZN(n756) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n756), .A2(n755), .ZN(n995) );
  NAND2_X1 U847 ( .A1(n768), .A2(n995), .ZN(n763) );
  AND2_X1 U848 ( .A1(n756), .A2(KEYINPUT33), .ZN(n757) );
  INV_X1 U849 ( .A(n759), .ZN(n777) );
  AND2_X1 U850 ( .A1(n757), .A2(n777), .ZN(n758) );
  XNOR2_X1 U851 ( .A(G1981), .B(G305), .ZN(n1003) );
  OR2_X1 U852 ( .A1(n758), .A2(n1003), .ZN(n764) );
  OR2_X1 U853 ( .A1(n759), .A2(n764), .ZN(n761) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n994) );
  INV_X1 U855 ( .A(n764), .ZN(n765) );
  AND2_X1 U856 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n767), .A2(n766), .ZN(n782) );
  INV_X1 U858 ( .A(n768), .ZN(n775) );
  NAND2_X1 U859 ( .A1(G8), .A2(G166), .ZN(n769) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n769), .ZN(n770) );
  XOR2_X1 U861 ( .A(KEYINPUT103), .B(n770), .Z(n773) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U863 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  AND2_X1 U864 ( .A1(n772), .A2(n777), .ZN(n776) );
  OR2_X1 U865 ( .A1(n773), .A2(n776), .ZN(n774) );
  NOR2_X1 U866 ( .A1(n775), .A2(n774), .ZN(n780) );
  INV_X1 U867 ( .A(n776), .ZN(n778) );
  AND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U869 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n784) );
  XNOR2_X1 U871 ( .A(n784), .B(n783), .ZN(n818) );
  XOR2_X1 U872 ( .A(G1986), .B(G290), .Z(n985) );
  NAND2_X1 U873 ( .A1(G95), .A2(n906), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G119), .A2(n521), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n901), .A2(G107), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT92), .B(n787), .Z(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n904), .A2(G131), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n892) );
  NAND2_X1 U881 ( .A1(G1991), .A2(n892), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT93), .ZN(n801) );
  NAND2_X1 U883 ( .A1(n906), .A2(G105), .ZN(n793) );
  XNOR2_X1 U884 ( .A(n793), .B(KEYINPUT38), .ZN(n795) );
  NAND2_X1 U885 ( .A1(G117), .A2(n901), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n799) );
  NAND2_X1 U887 ( .A1(G141), .A2(n904), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G129), .A2(n521), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n896) );
  NOR2_X1 U891 ( .A1(n965), .A2(n896), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n820) );
  NAND2_X1 U893 ( .A1(n985), .A2(n820), .ZN(n805) );
  INV_X1 U894 ( .A(n802), .ZN(n804) );
  NOR2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n831) );
  NAND2_X1 U896 ( .A1(n805), .A2(n831), .ZN(n816) );
  XOR2_X1 U897 ( .A(G2067), .B(KEYINPUT37), .Z(n830) );
  NAND2_X1 U898 ( .A1(G104), .A2(n906), .ZN(n807) );
  NAND2_X1 U899 ( .A1(G140), .A2(n904), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n808) );
  XNOR2_X1 U901 ( .A(KEYINPUT34), .B(n808), .ZN(n814) );
  NAND2_X1 U902 ( .A1(G116), .A2(n901), .ZN(n810) );
  NAND2_X1 U903 ( .A1(G128), .A2(n521), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U905 ( .A(KEYINPUT91), .B(n811), .ZN(n812) );
  XNOR2_X1 U906 ( .A(KEYINPUT35), .B(n812), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XOR2_X1 U908 ( .A(KEYINPUT36), .B(n815), .Z(n916) );
  AND2_X1 U909 ( .A1(n830), .A2(n916), .ZN(n945) );
  NAND2_X1 U910 ( .A1(n945), .A2(n831), .ZN(n819) );
  AND2_X1 U911 ( .A1(n816), .A2(n819), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n835) );
  INV_X1 U913 ( .A(n819), .ZN(n829) );
  AND2_X1 U914 ( .A1(n965), .A2(n896), .ZN(n950) );
  INV_X1 U915 ( .A(n820), .ZN(n941) );
  NOR2_X1 U916 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U917 ( .A1(G1991), .A2(n892), .ZN(n821) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(n821), .Z(n939) );
  NOR2_X1 U919 ( .A1(n822), .A2(n939), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n823), .B(KEYINPUT106), .ZN(n824) );
  NOR2_X1 U921 ( .A1(n941), .A2(n824), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n950), .A2(n825), .ZN(n826) );
  XNOR2_X1 U923 ( .A(KEYINPUT39), .B(n826), .ZN(n827) );
  NAND2_X1 U924 ( .A1(n827), .A2(n831), .ZN(n828) );
  OR2_X1 U925 ( .A1(n829), .A2(n828), .ZN(n833) );
  NOR2_X1 U926 ( .A1(n830), .A2(n916), .ZN(n937) );
  NAND2_X1 U927 ( .A1(n937), .A2(n831), .ZN(n832) );
  AND2_X1 U928 ( .A1(n833), .A2(n832), .ZN(n834) );
  NAND2_X1 U929 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n836), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n837), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U933 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G108), .ZN(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G69), .ZN(G235) );
  NOR2_X1 U941 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT109), .B(n843), .ZN(G261) );
  INV_X1 U943 ( .A(G261), .ZN(G325) );
  NOR2_X1 U944 ( .A1(G860), .A2(n844), .ZN(n845) );
  XOR2_X1 U945 ( .A(n846), .B(n845), .Z(G145) );
  XOR2_X1 U946 ( .A(G2454), .B(G2430), .Z(n848) );
  XNOR2_X1 U947 ( .A(G2451), .B(G2446), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n855) );
  XOR2_X1 U949 ( .A(G2443), .B(G2427), .Z(n850) );
  XNOR2_X1 U950 ( .A(G2438), .B(KEYINPUT107), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n851), .B(G2435), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1348), .B(G1341), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n856), .A2(G14), .ZN(n857) );
  XOR2_X1 U957 ( .A(KEYINPUT108), .B(n857), .Z(G401) );
  XOR2_X1 U958 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT110), .B(G2678), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2090), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(G2096), .B(G2100), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U967 ( .A(G2084), .B(G2078), .Z(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(G227) );
  XOR2_X1 U969 ( .A(G1976), .B(G1971), .Z(n869) );
  XNOR2_X1 U970 ( .A(G1981), .B(G1966), .ZN(n868) );
  XNOR2_X1 U971 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U972 ( .A(n870), .B(KEYINPUT41), .Z(n872) );
  XNOR2_X1 U973 ( .A(G1996), .B(G1991), .ZN(n871) );
  XNOR2_X1 U974 ( .A(n872), .B(n871), .ZN(n876) );
  XOR2_X1 U975 ( .A(G2474), .B(G1956), .Z(n874) );
  XNOR2_X1 U976 ( .A(G1986), .B(G1961), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(n876), .B(n875), .ZN(G229) );
  NAND2_X1 U979 ( .A1(G124), .A2(n521), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n906), .A2(G100), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G136), .A2(n904), .ZN(n881) );
  NAND2_X1 U984 ( .A1(G112), .A2(n901), .ZN(n880) );
  NAND2_X1 U985 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U986 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U987 ( .A1(G103), .A2(n906), .ZN(n885) );
  NAND2_X1 U988 ( .A1(G139), .A2(n904), .ZN(n884) );
  NAND2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n891) );
  NAND2_X1 U990 ( .A1(n521), .A2(G127), .ZN(n886) );
  XNOR2_X1 U991 ( .A(n886), .B(KEYINPUT114), .ZN(n888) );
  NAND2_X1 U992 ( .A1(G115), .A2(n901), .ZN(n887) );
  NAND2_X1 U993 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n889), .Z(n890) );
  NOR2_X1 U995 ( .A1(n891), .A2(n890), .ZN(n931) );
  XNOR2_X1 U996 ( .A(G160), .B(n931), .ZN(n915) );
  XNOR2_X1 U997 ( .A(G164), .B(n938), .ZN(n900) );
  XNOR2_X1 U998 ( .A(KEYINPUT115), .B(KEYINPUT113), .ZN(n894) );
  XNOR2_X1 U999 ( .A(n892), .B(KEYINPUT48), .ZN(n893) );
  XNOR2_X1 U1000 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U1001 ( .A(n895), .B(KEYINPUT46), .Z(n898) );
  XNOR2_X1 U1002 ( .A(n896), .B(G162), .ZN(n897) );
  XNOR2_X1 U1003 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U1004 ( .A(n900), .B(n899), .ZN(n913) );
  NAND2_X1 U1005 ( .A1(G118), .A2(n901), .ZN(n903) );
  NAND2_X1 U1006 ( .A1(G130), .A2(n521), .ZN(n902) );
  NAND2_X1 U1007 ( .A1(n903), .A2(n902), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(n904), .A2(G142), .ZN(n905) );
  XNOR2_X1 U1009 ( .A(n905), .B(KEYINPUT112), .ZN(n908) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n906), .ZN(n907) );
  NAND2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1012 ( .A(n909), .B(KEYINPUT45), .Z(n910) );
  NOR2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1014 ( .A(n913), .B(n912), .Z(n914) );
  XNOR2_X1 U1015 ( .A(n915), .B(n914), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n917), .B(n916), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n918), .ZN(G395) );
  XOR2_X1 U1018 ( .A(n919), .B(G286), .Z(n922) );
  XNOR2_X1 U1019 ( .A(G171), .B(n920), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(n922), .B(n921), .ZN(n923) );
  XNOR2_X1 U1021 ( .A(n923), .B(n987), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G37), .A2(n924), .ZN(G397) );
  OR2_X1 U1023 ( .A1(G401), .A2(n925), .ZN(n928) );
  NOR2_X1 U1024 ( .A1(G227), .A2(G229), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(KEYINPUT49), .B(n926), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1029 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1030 ( .A(G2072), .B(n931), .ZN(n933) );
  XNOR2_X1 U1031 ( .A(G164), .B(G2078), .ZN(n932) );
  NAND2_X1 U1032 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1033 ( .A(n934), .B(KEYINPUT119), .Z(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT50), .B(n935), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n948) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G160), .B(G2084), .Z(n940) );
  NOR2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(n946), .B(KEYINPUT116), .ZN(n947) );
  NAND2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n955) );
  XOR2_X1 U1043 ( .A(G2090), .B(G162), .Z(n949) );
  NOR2_X1 U1044 ( .A1(n950), .A2(n949), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT51), .B(n951), .Z(n953) );
  XNOR2_X1 U1046 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(n953), .B(n952), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(KEYINPUT52), .B(n956), .ZN(n958) );
  INV_X1 U1050 ( .A(KEYINPUT55), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1052 ( .A1(n959), .A2(G29), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT120), .B(n960), .ZN(n1040) );
  XNOR2_X1 U1054 ( .A(G2067), .B(G26), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(G33), .B(G2072), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n971) );
  XOR2_X1 U1057 ( .A(G1991), .B(G25), .Z(n963) );
  NAND2_X1 U1058 ( .A1(n963), .A2(G28), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(n964), .B(G27), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n965), .B(G32), .ZN(n966) );
  NAND2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT53), .B(n972), .ZN(n977) );
  XOR2_X1 U1065 ( .A(KEYINPUT54), .B(KEYINPUT122), .Z(n974) );
  XNOR2_X1 U1066 ( .A(G34), .B(KEYINPUT121), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n974), .B(n973), .ZN(n975) );
  XOR2_X1 U1068 ( .A(G2084), .B(n975), .Z(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(G35), .B(G2090), .ZN(n978) );
  NOR2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(KEYINPUT55), .B(n980), .ZN(n982) );
  INV_X1 U1073 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(G11), .ZN(n1038) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1010) );
  XNOR2_X1 U1077 ( .A(n984), .B(G1956), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n1001) );
  XNOR2_X1 U1079 ( .A(G301), .B(G1961), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(n987), .B(G1341), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n999) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT125), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(n991), .B(n990), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(G1971), .A2(G303), .ZN(n992) );
  NAND2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(G168), .B(G1966), .Z(n1002) );
  NOR2_X1 U1091 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1004), .Z(n1006) );
  XOR2_X1 U1093 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(n1006), .B(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1036) );
  INV_X1 U1097 ( .A(G16), .ZN(n1034) );
  XOR2_X1 U1098 ( .A(G1348), .B(KEYINPUT59), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(G4), .B(n1011), .ZN(n1019) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G6), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G19), .B(G1341), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1014), .Z(n1016) );
  XNOR2_X1 U1104 ( .A(G1956), .B(G20), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT127), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1020), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G21), .ZN(n1022) );
  XNOR2_X1 U1110 ( .A(G5), .B(G1961), .ZN(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1031) );
  XNOR2_X1 U1113 ( .A(G1971), .B(G22), .ZN(n1026) );
  XNOR2_X1 U1114 ( .A(G23), .B(G1976), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1028) );
  XOR2_X1 U1116 ( .A(G1986), .B(G24), .Z(n1027) );
  NAND2_X1 U1117 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(KEYINPUT58), .B(n1029), .ZN(n1030) );
  NOR2_X1 U1119 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1120 ( .A(KEYINPUT61), .B(n1032), .ZN(n1033) );
  NAND2_X1 U1121 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NAND2_X1 U1122 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NOR2_X1 U1123 ( .A1(n1038), .A2(n1037), .ZN(n1039) );
  NAND2_X1 U1124 ( .A1(n1040), .A2(n1039), .ZN(n1041) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1041), .Z(G311) );
  INV_X1 U1126 ( .A(G311), .ZN(G150) );
endmodule

