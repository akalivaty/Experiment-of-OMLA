//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1201,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n205), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n224), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT2), .B(G226), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G50), .B(G68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G351));
  AOI21_X1  g0041(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n242));
  OR2_X1    g0042(.A1(KEYINPUT64), .A2(G1), .ZN(new_n243));
  NAND2_X1  g0043(.A1(KEYINPUT64), .A2(G1), .ZN(new_n244));
  AND2_X1   g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G41), .A2(G45), .ZN(new_n246));
  INV_X1    g0046(.A(new_n246), .ZN(new_n247));
  AOI21_X1  g0047(.A(new_n242), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G226), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  INV_X1    g0050(.A(new_n211), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n253), .A2(new_n254), .A3(new_n247), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(G223), .B1(new_n265), .B2(G77), .ZN(new_n266));
  INV_X1    g0066(.A(G222), .ZN(new_n267));
  AOI21_X1  g0067(.A(G1698), .B1(new_n260), .B2(new_n261), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n256), .B1(new_n270), .B2(new_n242), .ZN(new_n271));
  AND2_X1   g0071(.A1(KEYINPUT65), .A2(G179), .ZN(new_n272));
  NOR2_X1   g0072(.A1(KEYINPUT65), .A2(G179), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G20), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G150), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT8), .B(G58), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n212), .A2(G33), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n277), .B1(new_n201), .B2(new_n212), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n211), .ZN(new_n282));
  INV_X1    g0082(.A(G50), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n243), .A2(G13), .A3(G20), .A4(new_n244), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n280), .A2(new_n282), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n243), .A2(new_n244), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(new_n212), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n286), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n275), .B(new_n293), .C1(G169), .C2(new_n271), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT66), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n248), .A2(G244), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n255), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n262), .A2(G238), .B1(new_n265), .B2(G107), .ZN(new_n298));
  INV_X1    g0098(.A(G232), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n298), .B1(new_n299), .B2(new_n269), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(new_n242), .B2(new_n300), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n301), .A2(G169), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n274), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n288), .A2(new_n290), .A3(new_n202), .ZN(new_n304));
  INV_X1    g0104(.A(new_n278), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n276), .B1(G20), .B2(G77), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT15), .B(G87), .Z(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n306), .B1(new_n279), .B2(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n304), .B1(new_n309), .B2(new_n282), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n285), .A2(new_n202), .ZN(new_n311));
  XNOR2_X1  g0111(.A(new_n311), .B(KEYINPUT67), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n302), .A2(new_n303), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n313), .B1(new_n301), .B2(G190), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n301), .ZN(new_n317));
  AND3_X1   g0117(.A1(new_n295), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n271), .A2(new_n316), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n319), .B1(G190), .B2(new_n271), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT9), .ZN(new_n321));
  OR2_X1    g0121(.A1(new_n293), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n293), .A2(new_n321), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n320), .A2(new_n322), .A3(new_n324), .A4(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n323), .A2(KEYINPUT10), .ZN(new_n327));
  XOR2_X1   g0127(.A(new_n326), .B(new_n327), .Z(new_n328));
  NAND2_X1  g0128(.A1(new_n248), .A2(G238), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n255), .ZN(new_n330));
  NAND2_X1  g0130(.A1(G33), .A2(G97), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n299), .A2(G1698), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G226), .B2(G1698), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n331), .B1(new_n333), .B2(new_n265), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n334), .A2(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n251), .A2(new_n252), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n334), .B2(KEYINPUT69), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n330), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT13), .ZN(new_n339));
  AND2_X1   g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(new_n339), .ZN(new_n341));
  OAI21_X1  g0141(.A(G169), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n338), .A2(new_n339), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n338), .A2(new_n339), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(G169), .A3(new_n343), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(G179), .A3(new_n347), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n276), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n283), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n279), .A2(new_n202), .B1(new_n212), .B2(G68), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n282), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n291), .A2(G68), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n288), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n284), .A2(G68), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT12), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n351), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n348), .A2(G200), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n346), .A2(G190), .A3(new_n347), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n318), .A2(new_n328), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G58), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n216), .ZN(new_n369));
  NOR2_X1   g0169(.A1(G58), .A2(G68), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n371), .B1(new_n372), .B2(new_n352), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT72), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n260), .A2(new_n212), .A3(new_n261), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT7), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n260), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n261), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n380), .A2(KEYINPUT7), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n377), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  AND4_X1   g0184(.A1(new_n376), .A2(new_n382), .A3(G68), .A4(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT7), .B1(new_n265), .B2(new_n212), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n216), .B1(new_n386), .B2(new_n383), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n376), .B1(new_n387), .B2(new_n382), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n375), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n216), .B1(new_n379), .B2(new_n381), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n374), .B1(new_n390), .B2(new_n373), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT73), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT73), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(new_n374), .C1(new_n390), .C2(new_n373), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n389), .A2(new_n282), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n290), .A2(new_n278), .ZN(new_n396));
  OR2_X1    g0196(.A1(new_n396), .A2(KEYINPUT74), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n288), .B1(new_n396), .B2(KEYINPUT74), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n397), .A2(new_n398), .B1(new_n278), .B2(new_n285), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G223), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n257), .ZN(new_n402));
  INV_X1    g0202(.A(G226), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G1698), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(new_n404), .C1(new_n263), .C2(new_n264), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G87), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n336), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI211_X1 g0208(.A(G232), .B(new_n336), .C1(new_n289), .C2(new_n246), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n255), .A3(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n274), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(G169), .B2(new_n410), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n400), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT18), .ZN(new_n415));
  INV_X1    g0215(.A(G190), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n408), .A2(new_n416), .A3(new_n255), .A4(new_n409), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n409), .A2(new_n255), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n316), .B1(new_n418), .B2(new_n407), .ZN(new_n419));
  AND3_X1   g0219(.A1(new_n417), .A2(new_n419), .A3(KEYINPUT75), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT75), .B1(new_n417), .B2(new_n419), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n395), .A2(new_n399), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT17), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT18), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n400), .A2(new_n425), .A3(new_n413), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n395), .A2(new_n422), .A3(new_n399), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n415), .A2(new_n424), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n367), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT5), .B(G41), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n245), .A2(new_n253), .A3(G45), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n243), .A2(G45), .A3(new_n244), .ZN(new_n434));
  AND2_X1   g0234(.A1(KEYINPUT5), .A2(G41), .ZN(new_n435));
  NOR2_X1   g0235(.A1(KEYINPUT5), .A2(G41), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(G257), .B(new_n336), .C1(new_n434), .C2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(G244), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT4), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n439), .A2(KEYINPUT77), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n440), .B1(new_n439), .B2(KEYINPUT77), .ZN(new_n442));
  OAI211_X1 g0242(.A(G250), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n443));
  NAND2_X1  g0243(.A1(G33), .A2(G283), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n441), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n433), .B(new_n438), .C1(new_n446), .C2(new_n336), .ZN(new_n447));
  INV_X1    g0247(.A(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n276), .A2(G77), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT76), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT6), .ZN(new_n451));
  INV_X1    g0251(.A(G97), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n451), .A2(new_n452), .A3(G107), .ZN(new_n453));
  XNOR2_X1  g0253(.A(G97), .B(G107), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n453), .B1(new_n451), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n450), .B1(new_n212), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n379), .B2(new_n381), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n282), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n284), .A2(G97), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n288), .B1(G33), .B2(new_n245), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G97), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n447), .A2(new_n448), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT78), .B1(new_n446), .B2(new_n336), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n439), .A2(KEYINPUT77), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n439), .A2(KEYINPUT77), .A3(new_n440), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n466), .A2(new_n467), .A3(new_n443), .A4(new_n444), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT78), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n468), .A2(new_n469), .A3(new_n242), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n433), .A2(new_n438), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n433), .A2(new_n438), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n464), .A2(new_n470), .A3(new_n274), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n463), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n464), .A2(new_n470), .A3(new_n475), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT80), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n464), .A2(new_n470), .A3(KEYINPUT80), .A4(new_n475), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(G200), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n459), .A2(new_n462), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n471), .B1(new_n468), .B2(new_n242), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(G190), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n478), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n212), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT22), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n260), .A2(new_n261), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n490), .A2(new_n491), .A3(new_n212), .A4(G87), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT83), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G116), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(G20), .ZN(new_n497));
  OR3_X1    g0297(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n212), .A2(KEYINPUT83), .A3(G33), .A4(G116), .ZN(new_n499));
  OAI21_X1  g0299(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n500));
  AND4_X1   g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n493), .A2(new_n494), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n494), .B1(new_n493), .B2(new_n501), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n282), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n284), .A2(G107), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(KEYINPUT25), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(new_n507), .B1(new_n461), .B2(G107), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n268), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT84), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n262), .B2(G257), .ZN(new_n512));
  OAI211_X1 g0312(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(KEYINPUT84), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n242), .ZN(new_n516));
  INV_X1    g0316(.A(G179), .ZN(new_n517));
  OAI211_X1 g0317(.A(G264), .B(new_n336), .C1(new_n434), .C2(new_n437), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n516), .A2(new_n517), .A3(new_n433), .A4(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(G250), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n520), .B1(new_n259), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n262), .A2(new_n511), .A3(G257), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n513), .A2(KEYINPUT84), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n433), .B(new_n518), .C1(new_n525), .C2(new_n336), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n448), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n509), .A2(new_n519), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G200), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n516), .A2(G190), .A3(new_n433), .A4(new_n518), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(new_n504), .A3(new_n508), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT85), .ZN(new_n533));
  XNOR2_X1  g0333(.A(new_n532), .B(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G238), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n535));
  OAI211_X1 g0335(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n496), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n242), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n242), .B1(new_n434), .B2(new_n219), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n243), .A2(G45), .A3(new_n250), .A4(new_n244), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G200), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n242), .A2(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT19), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n212), .B1(new_n331), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n218), .A2(new_n452), .A3(new_n457), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n212), .B(G68), .C1(new_n263), .C2(new_n264), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n546), .B1(new_n279), .B2(new_n452), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n282), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n284), .A2(new_n307), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n243), .A2(G33), .A3(new_n244), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n284), .A2(new_n287), .A3(new_n556), .A4(G87), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n543), .A2(new_n545), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n554), .B1(new_n552), .B2(new_n282), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n284), .A2(new_n307), .A3(new_n287), .A4(new_n556), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n538), .A2(new_n541), .A3(new_n274), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n562), .B(new_n563), .C1(G169), .C2(new_n544), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT81), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G116), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n285), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n284), .A2(new_n287), .A3(new_n556), .A4(G116), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n281), .A2(new_n211), .B1(G20), .B2(new_n567), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n444), .B(new_n212), .C1(G33), .C2(new_n452), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n570), .A2(KEYINPUT20), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(KEYINPUT20), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n568), .B(new_n569), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(G257), .B(new_n257), .C1(new_n263), .C2(new_n264), .ZN(new_n575));
  OAI211_X1 g0375(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n576));
  INV_X1    g0376(.A(G303), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n490), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n242), .ZN(new_n579));
  OAI211_X1 g0379(.A(G270), .B(new_n336), .C1(new_n434), .C2(new_n437), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n433), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n574), .B1(new_n582), .B2(G190), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT82), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT82), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n583), .A2(new_n587), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n559), .A2(new_n564), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT81), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n581), .A2(G169), .A3(new_n574), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n582), .A2(G179), .A3(new_n574), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n581), .A2(KEYINPUT21), .A3(G169), .A4(new_n574), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AND4_X1   g0397(.A1(new_n566), .A2(new_n589), .A3(new_n591), .A4(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n431), .A2(new_n487), .A3(new_n534), .A4(new_n598), .ZN(G372));
  AND2_X1   g0399(.A1(new_n415), .A2(new_n426), .ZN(new_n600));
  INV_X1    g0400(.A(new_n314), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n351), .B2(new_n362), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n366), .A2(new_n429), .A3(new_n424), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT87), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n328), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n608), .A2(new_n295), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n483), .A2(new_n486), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n597), .A2(new_n528), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n560), .A2(new_n612), .A3(new_n557), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n612), .B1(new_n560), .B2(new_n557), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n543), .B(new_n545), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n531), .A2(new_n564), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n610), .A2(new_n477), .A3(new_n611), .A4(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n615), .A2(new_n564), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n618), .B1(new_n477), .B2(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n591), .A2(new_n476), .A3(new_n463), .A4(new_n566), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(new_n618), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n617), .A2(new_n622), .A3(new_n564), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n431), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n609), .A2(new_n624), .ZN(G369));
  INV_X1    g0425(.A(G13), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(G20), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n245), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(KEYINPUT27), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(G213), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G343), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n574), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n589), .A2(new_n597), .A3(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n597), .B2(new_n634), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT88), .Z(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(G330), .ZN(new_n638));
  INV_X1    g0438(.A(new_n633), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n528), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n509), .A2(new_n633), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT89), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n534), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n638), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n597), .A2(new_n633), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n534), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n528), .B2(new_n633), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n644), .A2(new_n647), .ZN(G399));
  INV_X1    g0448(.A(new_n206), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n650), .A2(new_n254), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n548), .A2(G116), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n651), .A2(new_n652), .B1(new_n210), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g0453(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n653), .B(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n564), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n616), .A2(new_n611), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n656), .B1(new_n657), .B2(new_n487), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n477), .A2(new_n619), .ZN(new_n659));
  MUX2_X1   g0459(.A(new_n659), .B(new_n621), .S(new_n618), .Z(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n639), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT29), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n623), .A2(new_n639), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n663), .B1(KEYINPUT29), .B2(new_n664), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n598), .A2(new_n534), .A3(new_n487), .A4(new_n639), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT31), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n516), .A2(new_n518), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n581), .A2(new_n517), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n669), .A3(new_n485), .A4(new_n544), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT30), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n274), .ZN(new_n673));
  NOR3_X1   g0473(.A1(new_n582), .A2(new_n673), .A3(new_n544), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n479), .A2(new_n674), .A3(new_n526), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n668), .A2(new_n544), .A3(new_n669), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT91), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(KEYINPUT30), .A4(new_n485), .ZN(new_n679));
  OAI21_X1  g0479(.A(KEYINPUT91), .B1(new_n670), .B2(new_n671), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n667), .B1(new_n681), .B2(new_n639), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  INV_X1    g0483(.A(new_n676), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n639), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT31), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n666), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n665), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n655), .B1(new_n689), .B2(G1), .ZN(G364));
  XNOR2_X1  g0490(.A(new_n627), .B(KEYINPUT92), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G45), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n651), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n637), .B2(G330), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(G330), .B2(new_n637), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n211), .B1(G20), .B2(new_n448), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n212), .A2(new_n416), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n316), .A2(G179), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n212), .A2(G190), .ZN(new_n703));
  NOR2_X1   g0503(.A1(G179), .A2(G200), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI22_X1  g0506(.A1(G303), .A2(new_n702), .B1(new_n706), .B2(G329), .ZN(new_n707));
  INV_X1    g0507(.A(G283), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n700), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n707), .B(new_n265), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n673), .A2(new_n316), .A3(new_n699), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n710), .B1(G322), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n212), .A2(new_n316), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n673), .A2(G190), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n704), .A2(G190), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G20), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n716), .A2(G326), .B1(G294), .B2(new_n718), .ZN(new_n719));
  OR2_X1    g0519(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(KEYINPUT94), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n673), .A2(new_n316), .A3(new_n703), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n673), .A2(new_n416), .A3(new_n714), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g0525(.A(KEYINPUT33), .B(G317), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n723), .A2(G311), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n713), .A2(new_n720), .A3(new_n721), .A4(new_n727), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n283), .A2(new_n715), .B1(new_n724), .B2(new_n216), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(G58), .B2(new_n712), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n702), .A2(G87), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n731), .B(new_n490), .C1(new_n457), .C2(new_n709), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(G77), .B2(new_n723), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n705), .A2(KEYINPUT32), .A3(new_n372), .ZN(new_n734));
  OAI21_X1  g0534(.A(KEYINPUT32), .B1(new_n705), .B2(new_n372), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n718), .A2(G97), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n730), .A2(new_n733), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n698), .B1(new_n728), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n490), .A2(new_n206), .ZN(new_n740));
  INV_X1    g0540(.A(G355), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n740), .A2(new_n741), .B1(G116), .B2(new_n206), .ZN(new_n742));
  INV_X1    g0542(.A(G45), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n237), .A2(new_n743), .ZN(new_n744));
  AOI211_X1 g0544(.A(new_n490), .B(new_n649), .C1(new_n743), .C2(new_n210), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(KEYINPUT93), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n697), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n748), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n693), .B(new_n739), .C1(new_n747), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n751), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n637), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n696), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(G396));
  NOR2_X1   g0559(.A1(new_n314), .A2(new_n633), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n313), .A2(new_n633), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n317), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(new_n762), .B2(new_n314), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n623), .A2(new_n639), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT97), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n623), .A2(new_n766), .A3(new_n639), .A4(new_n763), .ZN(new_n767));
  INV_X1    g0567(.A(new_n763), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n765), .A2(new_n767), .B1(new_n664), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(new_n688), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT98), .Z(new_n771));
  OAI21_X1  g0571(.A(new_n693), .B1(new_n769), .B2(new_n688), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G137), .A2(new_n716), .B1(new_n725), .B2(G150), .ZN(new_n774));
  INV_X1    g0574(.A(G143), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n774), .B1(new_n775), .B2(new_n711), .C1(new_n372), .C2(new_n722), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT34), .Z(new_n777));
  INV_X1    g0577(.A(new_n718), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n368), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n490), .B1(new_n701), .B2(new_n283), .ZN(new_n780));
  INV_X1    g0580(.A(new_n709), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G68), .ZN(new_n782));
  INV_X1    g0582(.A(G132), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n783), .B2(new_n705), .ZN(new_n784));
  NOR4_X1   g0584(.A1(new_n777), .A2(new_n779), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G107), .A2(new_n702), .B1(new_n706), .B2(G311), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n490), .B1(new_n781), .B2(G87), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n786), .A2(new_n736), .A3(new_n787), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G116), .A2(new_n723), .B1(new_n716), .B2(G303), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n521), .B2(new_n711), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n788), .B(new_n790), .C1(G283), .C2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n697), .B1(new_n785), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n698), .A2(new_n750), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n694), .B1(G77), .B2(new_n797), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT95), .Z(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n749), .B2(new_n768), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n773), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G384));
  NOR2_X1   g0603(.A1(new_n691), .A2(new_n245), .ZN(new_n804));
  INV_X1    g0604(.A(new_n631), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n600), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n760), .B1(new_n765), .B2(new_n767), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n362), .A2(new_n633), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n363), .A2(new_n366), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n366), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n362), .B(new_n633), .C1(new_n810), .C2(new_n351), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT38), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n384), .A2(G68), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT72), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n387), .A2(new_n376), .A3(new_n382), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n373), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n389), .B(new_n282), .C1(new_n821), .C2(KEYINPUT16), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n412), .B1(new_n822), .B2(new_n399), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n816), .B1(new_n423), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n399), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n385), .A2(new_n388), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n374), .B1(new_n826), .B2(new_n373), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n819), .A2(new_n820), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n287), .B1(new_n828), .B2(new_n375), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n825), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(KEYINPUT99), .B(new_n427), .C1(new_n830), .C2(new_n412), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n631), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n824), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT100), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT37), .ZN(new_n835));
  INV_X1    g0635(.A(new_n832), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n430), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n400), .A2(new_n805), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT37), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n414), .A2(new_n839), .A3(new_n840), .A4(new_n427), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(KEYINPUT100), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(KEYINPUT37), .B2(new_n833), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n815), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n833), .A2(KEYINPUT37), .ZN(new_n845));
  INV_X1    g0645(.A(new_n842), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n847), .A2(KEYINPUT38), .A3(new_n835), .A4(new_n837), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n806), .B1(new_n814), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n414), .A2(new_n839), .A3(new_n427), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n841), .ZN(new_n853));
  INV_X1    g0653(.A(new_n430), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n854), .B2(new_n839), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n815), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT39), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n351), .A2(new_n362), .A3(new_n639), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n844), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n859), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n850), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n665), .A2(new_n431), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n609), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n864), .B(new_n866), .Z(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT102), .B1(new_n685), .B2(KEYINPUT31), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n869), .B(new_n667), .C1(new_n681), .C2(new_n639), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n868), .A2(new_n666), .A3(new_n686), .A4(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n872), .A2(new_n430), .A3(new_n367), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n768), .B1(new_n809), .B2(new_n811), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n849), .A2(new_n876), .ZN(new_n877));
  XOR2_X1   g0677(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n876), .A2(new_n857), .A3(KEYINPUT40), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n873), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(G330), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n873), .A3(new_n880), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n804), .B1(new_n867), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n867), .B2(new_n885), .ZN(new_n887));
  INV_X1    g0687(.A(new_n455), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n888), .A2(KEYINPUT35), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(KEYINPUT35), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n889), .A2(G116), .A3(new_n213), .A4(new_n890), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n891), .B(KEYINPUT36), .ZN(new_n892));
  NOR3_X1   g0692(.A1(new_n369), .A2(new_n209), .A3(new_n202), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n216), .A2(G50), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n626), .B(new_n289), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n887), .A2(new_n892), .A3(new_n895), .ZN(G367));
  OR3_X1    g0696(.A1(new_n639), .A2(new_n614), .A3(new_n613), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n564), .A3(new_n615), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n564), .B2(new_n897), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT43), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT104), .Z(new_n901));
  NAND2_X1  g0701(.A1(new_n484), .A2(new_n633), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n487), .A2(new_n902), .B1(new_n478), .B2(new_n633), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n646), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n528), .B1(new_n483), .B2(new_n486), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n639), .B1(new_n906), .B2(new_n478), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n904), .A2(KEYINPUT42), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT103), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n899), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n899), .A2(new_n911), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n913), .A2(KEYINPUT43), .A3(new_n914), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n910), .B(new_n915), .Z(new_n916));
  INV_X1    g0716(.A(new_n644), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n903), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT105), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n916), .A2(new_n918), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n916), .A2(KEYINPUT105), .A3(new_n918), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n650), .B(KEYINPUT41), .Z(new_n925));
  NAND2_X1  g0725(.A1(new_n643), .A2(new_n640), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n646), .B1(new_n926), .B2(new_n645), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n638), .B(new_n927), .Z(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n689), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n647), .A2(new_n903), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT44), .Z(new_n931));
  NOR2_X1   g0731(.A1(new_n647), .A2(new_n903), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT45), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(KEYINPUT106), .A3(new_n644), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n644), .A2(KEYINPUT106), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(new_n933), .A3(new_n931), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n929), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n925), .B1(new_n938), .B2(new_n689), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n692), .A2(G1), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT107), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n924), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n753), .B1(new_n649), .B2(new_n307), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n649), .A2(new_n490), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n233), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n693), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(G150), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n775), .A2(new_n715), .B1(new_n711), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n949), .B1(G50), .B2(new_n723), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n778), .A2(new_n216), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n706), .A2(G137), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n490), .B1(new_n701), .B2(new_n368), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n709), .A2(new_n202), .ZN(new_n954));
  NOR4_X1   g0754(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n950), .B(new_n955), .C1(new_n372), .C2(new_n793), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n701), .A2(new_n567), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT46), .ZN(new_n958));
  INV_X1    g0758(.A(G311), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n577), .A2(new_n711), .B1(new_n715), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(G317), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n265), .B1(new_n705), .B2(new_n961), .C1(new_n452), .C2(new_n709), .ZN(new_n962));
  NOR3_X1   g0762(.A1(new_n958), .A2(new_n960), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(new_n521), .B2(new_n793), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n722), .A2(new_n708), .B1(new_n778), .B2(new_n457), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT108), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n956), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT47), .Z(new_n968));
  OAI221_X1 g0768(.A(new_n947), .B1(new_n899), .B2(new_n756), .C1(new_n968), .C2(new_n698), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n943), .A2(new_n969), .ZN(G387));
  NAND2_X1  g0770(.A1(new_n928), .A2(new_n941), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT109), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n230), .A2(new_n743), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT110), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n305), .A2(new_n283), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT50), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n652), .B(new_n743), .C1(new_n216), .C2(new_n202), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n945), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n973), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n974), .B2(new_n978), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(G107), .B2(new_n206), .C1(new_n652), .C2(new_n740), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n693), .B1(new_n981), .B2(new_n752), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G77), .A2(new_n702), .B1(new_n706), .B2(G150), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n983), .B(new_n490), .C1(new_n452), .C2(new_n709), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n216), .A2(new_n722), .B1(new_n724), .B2(new_n278), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n283), .A2(new_n711), .B1(new_n715), .B2(new_n372), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n778), .A2(new_n308), .ZN(new_n987));
  NOR4_X1   g0787(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n702), .A2(G294), .B1(new_n718), .B2(G283), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n577), .A2(new_n722), .B1(new_n711), .B2(new_n961), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n716), .A2(G322), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n959), .C2(new_n793), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT48), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n989), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT112), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n994), .B2(new_n993), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n997), .A2(KEYINPUT49), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n490), .B1(new_n706), .B2(G326), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n567), .B2(new_n709), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n997), .B2(KEYINPUT49), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n988), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n982), .B1(new_n926), .B2(new_n756), .C1(new_n1002), .C2(new_n698), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n972), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n650), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n929), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n689), .B2(new_n928), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(G393));
  XNOR2_X1  g0808(.A(new_n934), .B(new_n917), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n938), .B(new_n650), .C1(new_n1009), .C2(new_n929), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n240), .A2(new_n945), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n752), .B1(new_n452), .B2(new_n206), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n701), .A2(new_n708), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n265), .B1(new_n709), .B2(new_n457), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G322), .C2(new_n706), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1015), .B1(new_n567), .B2(new_n778), .C1(new_n521), .C2(new_n722), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(G303), .B2(new_n794), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n959), .A2(new_n711), .B1(new_n715), .B2(new_n961), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT52), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n948), .A2(new_n715), .B1(new_n711), .B2(new_n372), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT51), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n778), .A2(new_n202), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n490), .B1(new_n709), .B2(new_n218), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n701), .A2(new_n216), .B1(new_n705), .B2(new_n775), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n278), .B2(new_n722), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G50), .B2(new_n794), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n1017), .A2(new_n1019), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n694), .B1(new_n1011), .B2(new_n1012), .C1(new_n1028), .C2(new_n698), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n903), .B2(new_n751), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(new_n1009), .B2(new_n941), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1010), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT113), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1010), .A2(KEYINPUT113), .A3(new_n1031), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(G390));
  INV_X1    g0836(.A(KEYINPUT116), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n860), .B1(new_n807), .B2(new_n813), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n844), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n1039));
  AOI21_X1  g0839(.A(KEYINPUT39), .B1(new_n848), .B2(new_n856), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1038), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n762), .A2(new_n314), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n633), .B(new_n1043), .C1(new_n658), .C2(new_n660), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT114), .B1(new_n1044), .B2(new_n760), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT114), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n760), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n662), .C2(new_n1043), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1045), .A2(new_n1048), .A3(new_n812), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n861), .B1(new_n848), .B2(new_n856), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1041), .A2(KEYINPUT115), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n768), .A2(new_n882), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n871), .A2(new_n812), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT115), .B1(new_n1041), .B2(new_n1051), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1037), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n687), .A2(new_n812), .A3(new_n1053), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1041), .A2(new_n1051), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n765), .A2(new_n767), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n1047), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n812), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n860), .A2(new_n1064), .B1(new_n859), .B2(new_n862), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1051), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1067), .A2(KEYINPUT116), .A3(new_n1055), .A4(new_n1052), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1058), .A2(new_n1060), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n431), .A2(G330), .A3(new_n871), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT117), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n873), .A2(KEYINPUT117), .A3(G330), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n866), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n871), .A2(new_n1053), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1059), .B(new_n1075), .C1(new_n812), .C2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n812), .B1(new_n687), .B2(new_n1053), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1063), .B1(new_n1055), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1074), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1069), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1073), .A2(new_n1072), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(new_n609), .A3(new_n865), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1079), .B2(new_n1077), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1058), .A2(new_n1060), .A3(new_n1068), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1082), .A2(new_n650), .A3(new_n1086), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1058), .A2(new_n941), .A3(new_n1068), .A4(new_n1060), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n694), .B1(new_n305), .B2(new_n797), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n794), .A2(G137), .ZN(new_n1090));
  INV_X1    g0890(.A(G125), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n490), .B1(new_n705), .B2(new_n1091), .C1(new_n283), .C2(new_n709), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G159), .B2(new_n718), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n702), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n701), .B2(new_n948), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n716), .A2(G128), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g0897(.A(KEYINPUT54), .B(G143), .Z(new_n1098));
  AOI22_X1  g0898(.A1(G132), .A2(new_n712), .B1(new_n723), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1090), .A2(new_n1093), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n793), .A2(new_n457), .B1(new_n452), .B2(new_n722), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT118), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n706), .A2(G294), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n731), .A2(new_n782), .A3(new_n1103), .A4(new_n265), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n1104), .A2(new_n1022), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n567), .B2(new_n711), .C1(new_n708), .C2(new_n715), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1100), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1089), .B1(new_n1107), .B2(new_n697), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n859), .A2(new_n862), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1108), .B1(new_n1110), .B2(new_n750), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1088), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1087), .A2(new_n1113), .ZN(G378));
  NAND2_X1  g0914(.A1(new_n1086), .A2(new_n1074), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n875), .B1(new_n848), .B2(new_n844), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n878), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n880), .B(G330), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n328), .A2(new_n294), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n805), .A2(new_n293), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1119), .B(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1120), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1119), .B(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1122), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1118), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(new_n879), .A3(G330), .A4(new_n880), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n864), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n864), .A3(new_n1131), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1115), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n650), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT57), .B1(new_n1115), .B2(new_n1136), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(G97), .A2(new_n725), .B1(new_n712), .B2(G107), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1142), .B1(new_n567), .B2(new_n715), .C1(new_n308), .C2(new_n722), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n701), .A2(new_n202), .B1(new_n705), .B2(new_n708), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n709), .A2(new_n368), .ZN(new_n1145));
  INV_X1    g0945(.A(G41), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n265), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1143), .A2(new_n951), .A3(new_n1144), .A4(new_n1148), .ZN(new_n1149));
  OR2_X1    g0949(.A1(new_n1149), .A2(KEYINPUT58), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(KEYINPUT58), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1147), .B(new_n283), .C1(G33), .C2(G41), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G132), .A2(new_n725), .B1(new_n723), .B2(G137), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n702), .A2(new_n1098), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT119), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n712), .A2(G128), .B1(G150), .B2(new_n718), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n716), .A2(G125), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n259), .B(new_n1146), .C1(new_n709), .C2(new_n372), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(G124), .C2(new_n706), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1153), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n694), .B1(G50), .B2(new_n797), .C1(new_n1164), .C2(new_n698), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n1128), .B2(new_n749), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1136), .B2(new_n941), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1141), .A2(new_n1167), .ZN(G375));
  INV_X1    g0968(.A(new_n925), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1084), .A2(new_n1079), .A3(new_n1077), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1081), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT120), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n941), .B(KEYINPUT121), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n813), .A2(new_n749), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n694), .B1(G68), .B2(new_n797), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n794), .A2(new_n1098), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n778), .A2(new_n283), .ZN(new_n1177));
  INV_X1    g0977(.A(G128), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n701), .A2(new_n372), .B1(new_n705), .B2(new_n1178), .ZN(new_n1179));
  NOR4_X1   g0979(.A1(new_n1177), .A2(new_n1179), .A3(new_n265), .A4(new_n1145), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G137), .A2(new_n712), .B1(new_n723), .B2(G150), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n715), .A2(new_n783), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT122), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n1176), .A2(new_n1180), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n457), .A2(new_n722), .B1(new_n711), .B2(new_n708), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G294), .B2(new_n716), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n701), .A2(new_n452), .B1(new_n705), .B2(new_n577), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n987), .A2(new_n1187), .A3(new_n490), .A4(new_n954), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1186), .B(new_n1188), .C1(new_n567), .C2(new_n793), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1175), .B1(new_n1190), .B2(new_n697), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1080), .A2(new_n1173), .B1(new_n1174), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1172), .A2(new_n1192), .ZN(G381));
  INV_X1    g0993(.A(G390), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(G393), .A2(G396), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(new_n1195), .A3(new_n802), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1196), .A2(G387), .A3(G381), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1005), .B1(new_n1069), .B2(new_n1081), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1112), .B1(new_n1198), .B2(new_n1086), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1197), .A2(new_n1199), .A3(new_n1141), .A4(new_n1167), .ZN(G407));
  INV_X1    g1000(.A(G213), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(G343), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1199), .A2(new_n1202), .ZN(new_n1203));
  OAI211_X1 g1003(.A(G407), .B(G213), .C1(G375), .C2(new_n1203), .ZN(G409));
  NAND2_X1  g1004(.A1(G387), .A2(new_n1194), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(G390), .A2(new_n943), .A3(new_n969), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT124), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G387), .B2(new_n1194), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n758), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1195), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1207), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1205), .A2(new_n1208), .A3(new_n1206), .A4(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(G378), .B(new_n1167), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1166), .B1(new_n1136), .B2(new_n1173), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n1129), .A2(new_n864), .A3(new_n1131), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n864), .B1(new_n1131), .B2(new_n1129), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1169), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n1086), .B2(new_n1074), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT123), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(KEYINPUT123), .B(new_n1220), .C1(new_n1086), .C2(new_n1074), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1199), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1202), .B1(new_n1216), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1081), .A2(KEYINPUT60), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(new_n1170), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n650), .B1(new_n1227), .B2(new_n1170), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1192), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1230), .A2(new_n802), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1230), .A2(new_n802), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT62), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT125), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1202), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  AOI211_X1 g1038(.A(KEYINPUT125), .B(new_n1202), .C1(new_n1216), .C2(new_n1225), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1234), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1202), .A2(G2897), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1233), .A2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1215), .B1(new_n1242), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT61), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1213), .A2(new_n1252), .A3(new_n1214), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1226), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT63), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1233), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1251), .A2(new_n1258), .ZN(G405));
  NAND2_X1  g1059(.A1(G375), .A2(new_n1199), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1216), .A2(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(new_n1233), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1263), .A2(new_n1215), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1215), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1260), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1263), .A2(new_n1215), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1260), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1215), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1266), .A2(new_n1270), .ZN(G402));
endmodule


