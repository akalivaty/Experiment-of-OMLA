

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XOR2_X1 U326 ( .A(n345), .B(n420), .Z(n294) );
  XNOR2_X1 U327 ( .A(G106GAT), .B(n311), .ZN(n295) );
  NOR2_X1 U328 ( .A1(n466), .A2(n406), .ZN(n407) );
  XNOR2_X1 U329 ( .A(G43GAT), .B(KEYINPUT68), .ZN(n305) );
  XNOR2_X1 U330 ( .A(KEYINPUT112), .B(KEYINPUT48), .ZN(n415) );
  XNOR2_X1 U331 ( .A(n416), .B(n415), .ZN(n536) );
  XOR2_X1 U332 ( .A(n315), .B(n579), .Z(n494) );
  XNOR2_X1 U333 ( .A(n333), .B(n332), .ZN(n534) );
  XNOR2_X1 U334 ( .A(n458), .B(KEYINPUT62), .ZN(n459) );
  XNOR2_X1 U335 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U336 ( .A(n460), .B(n459), .ZN(G1355GAT) );
  XNOR2_X1 U337 ( .A(n465), .B(n464), .ZN(G1353GAT) );
  XNOR2_X1 U338 ( .A(KEYINPUT36), .B(KEYINPUT102), .ZN(n315) );
  INV_X1 U339 ( .A(KEYINPUT81), .ZN(n314) );
  XOR2_X1 U340 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n297) );
  XNOR2_X1 U341 ( .A(KEYINPUT9), .B(KEYINPUT79), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n298), .B(KEYINPUT10), .Z(n300) );
  XOR2_X1 U344 ( .A(G134GAT), .B(KEYINPUT80), .Z(n441) );
  XNOR2_X1 U345 ( .A(n441), .B(KEYINPUT66), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n345) );
  XNOR2_X1 U348 ( .A(G36GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n301), .B(G218GAT), .ZN(n420) );
  NAND2_X1 U350 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n294), .B(n302), .ZN(n303) );
  XOR2_X1 U352 ( .A(n304), .B(n303), .Z(n313) );
  XNOR2_X1 U353 ( .A(n305), .B(G29GAT), .ZN(n306) );
  XOR2_X1 U354 ( .A(n306), .B(KEYINPUT69), .Z(n308) );
  XNOR2_X1 U355 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n365) );
  XOR2_X1 U357 ( .A(KEYINPUT75), .B(G92GAT), .Z(n310) );
  XNOR2_X1 U358 ( .A(G99GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U360 ( .A(n365), .B(n295), .Z(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n561) );
  XNOR2_X1 U362 ( .A(n314), .B(n561), .ZN(n579) );
  XOR2_X1 U363 ( .A(KEYINPUT0), .B(G176GAT), .Z(n317) );
  XNOR2_X1 U364 ( .A(KEYINPUT65), .B(KEYINPUT86), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n333) );
  XOR2_X1 U366 ( .A(G190GAT), .B(G134GAT), .Z(n319) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G99GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n320), .B(KEYINPUT84), .Z(n322) );
  XOR2_X1 U370 ( .A(G120GAT), .B(G71GAT), .Z(n369) );
  XNOR2_X1 U371 ( .A(G169GAT), .B(n369), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n393) );
  XOR2_X1 U374 ( .A(n393), .B(KEYINPUT20), .Z(n324) );
  NAND2_X1 U375 ( .A1(G227GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U377 ( .A(n326), .B(n325), .Z(n331) );
  XOR2_X1 U378 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n328) );
  XNOR2_X1 U379 ( .A(KEYINPUT85), .B(G183GAT), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U381 ( .A(KEYINPUT17), .B(n329), .Z(n418) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(n418), .ZN(n330) );
  XNOR2_X1 U383 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U384 ( .A(KEYINPUT89), .B(KEYINPUT23), .Z(n335) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U387 ( .A(n336), .B(KEYINPUT24), .Z(n340) );
  XNOR2_X1 U388 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n337), .B(KEYINPUT2), .ZN(n440) );
  XNOR2_X1 U390 ( .A(G78GAT), .B(KEYINPUT74), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n338), .B(G148GAT), .ZN(n380) );
  XNOR2_X1 U392 ( .A(n440), .B(n380), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U394 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n342) );
  XNOR2_X1 U395 ( .A(G218GAT), .B(G106GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U397 ( .A(n344), .B(n343), .Z(n347) );
  XOR2_X1 U398 ( .A(G22GAT), .B(G155GAT), .Z(n392) );
  XNOR2_X1 U399 ( .A(n345), .B(n392), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U401 ( .A(KEYINPUT21), .B(G211GAT), .Z(n349) );
  XNOR2_X1 U402 ( .A(KEYINPUT87), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U404 ( .A(G197GAT), .B(n350), .Z(n417) );
  XOR2_X1 U405 ( .A(n351), .B(n417), .Z(n564) );
  NOR2_X1 U406 ( .A1(n534), .A2(n564), .ZN(n352) );
  XNOR2_X1 U407 ( .A(n352), .B(KEYINPUT26), .ZN(n550) );
  INV_X1 U408 ( .A(KEYINPUT54), .ZN(n431) );
  XOR2_X1 U409 ( .A(G141GAT), .B(G22GAT), .Z(n354) );
  XOR2_X1 U410 ( .A(G113GAT), .B(G1GAT), .Z(n447) );
  XOR2_X1 U411 ( .A(G169GAT), .B(G8GAT), .Z(n424) );
  XNOR2_X1 U412 ( .A(n447), .B(n424), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n355), .B(G36GAT), .Z(n360) );
  XOR2_X1 U415 ( .A(KEYINPUT70), .B(KEYINPUT29), .Z(n357) );
  XNOR2_X1 U416 ( .A(G197GAT), .B(G15GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U418 ( .A(n358), .B(G50GAT), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U420 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n362) );
  NAND2_X1 U421 ( .A1(G229GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U423 ( .A(n364), .B(n363), .Z(n367) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT71), .ZN(n366) );
  XOR2_X1 U425 ( .A(n367), .B(n366), .Z(n506) );
  INV_X1 U426 ( .A(n506), .ZN(n586) );
  XNOR2_X1 U427 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n368), .B(KEYINPUT72), .ZN(n396) );
  XOR2_X1 U429 ( .A(n396), .B(n369), .Z(n371) );
  NAND2_X1 U430 ( .A1(G230GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n371), .B(n370), .ZN(n384) );
  XOR2_X1 U432 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n373) );
  XNOR2_X1 U433 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n373), .B(n372), .ZN(n375) );
  INV_X1 U435 ( .A(KEYINPUT32), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U437 ( .A(G176GAT), .B(G64GAT), .Z(n419) );
  XNOR2_X1 U438 ( .A(G204GAT), .B(n419), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n379) );
  INV_X1 U440 ( .A(KEYINPUT33), .ZN(n378) );
  XNOR2_X1 U441 ( .A(n379), .B(n378), .ZN(n382) );
  XNOR2_X1 U442 ( .A(n380), .B(KEYINPUT78), .ZN(n381) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n385), .B(n295), .ZN(n466) );
  XOR2_X1 U446 ( .A(G64GAT), .B(G8GAT), .Z(n387) );
  XNOR2_X1 U447 ( .A(KEYINPUT70), .B(G1GAT), .ZN(n386) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U449 ( .A(KEYINPUT82), .B(KEYINPUT12), .Z(n389) );
  XNOR2_X1 U450 ( .A(KEYINPUT83), .B(KEYINPUT15), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n404) );
  XOR2_X1 U453 ( .A(n392), .B(G78GAT), .Z(n395) );
  XNOR2_X1 U454 ( .A(n393), .B(G211GAT), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U456 ( .A(KEYINPUT14), .B(n396), .Z(n398) );
  NAND2_X1 U457 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U459 ( .A(n400), .B(n399), .Z(n402) );
  XNOR2_X1 U460 ( .A(G183GAT), .B(G71GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U462 ( .A(n404), .B(n403), .Z(n590) );
  INV_X1 U463 ( .A(n590), .ZN(n493) );
  NOR2_X1 U464 ( .A1(n493), .A2(n494), .ZN(n405) );
  XOR2_X1 U465 ( .A(KEYINPUT45), .B(n405), .Z(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(KEYINPUT111), .ZN(n408) );
  NOR2_X1 U467 ( .A1(n586), .A2(n408), .ZN(n414) );
  XOR2_X1 U468 ( .A(n466), .B(KEYINPUT41), .Z(n574) );
  NAND2_X1 U469 ( .A1(n586), .A2(n574), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n409), .B(KEYINPUT46), .ZN(n411) );
  NOR2_X1 U471 ( .A1(n561), .A2(n590), .ZN(n410) );
  AND2_X1 U472 ( .A1(n411), .A2(n410), .ZN(n412) );
  XOR2_X1 U473 ( .A(n412), .B(KEYINPUT47), .Z(n413) );
  NOR2_X1 U474 ( .A1(n414), .A2(n413), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n428) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n422) );
  NAND2_X1 U477 ( .A1(G226GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U479 ( .A(n423), .B(KEYINPUT95), .Z(n426) );
  XNOR2_X1 U480 ( .A(n424), .B(G92GAT), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U482 ( .A(n428), .B(n427), .Z(n526) );
  INV_X1 U483 ( .A(n526), .ZN(n429) );
  NOR2_X1 U484 ( .A1(n536), .A2(n429), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n456) );
  XOR2_X1 U486 ( .A(G57GAT), .B(KEYINPUT92), .Z(n433) );
  XNOR2_X1 U487 ( .A(KEYINPUT90), .B(KEYINPUT1), .ZN(n432) );
  XNOR2_X1 U488 ( .A(n433), .B(n432), .ZN(n455) );
  XOR2_X1 U489 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n435) );
  XNOR2_X1 U490 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U492 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n436) );
  XNOR2_X1 U494 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U495 ( .A(n439), .B(n438), .Z(n453) );
  XOR2_X1 U496 ( .A(n441), .B(n440), .Z(n443) );
  NAND2_X1 U497 ( .A1(G225GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U498 ( .A(n443), .B(n442), .ZN(n451) );
  XOR2_X1 U499 ( .A(G155GAT), .B(G162GAT), .Z(n445) );
  XNOR2_X1 U500 ( .A(G127GAT), .B(G148GAT), .ZN(n444) );
  XNOR2_X1 U501 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U502 ( .A(n446), .B(G85GAT), .Z(n449) );
  XNOR2_X1 U503 ( .A(G29GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n476) );
  INV_X1 U508 ( .A(n476), .ZN(n523) );
  NOR2_X1 U509 ( .A1(n456), .A2(n523), .ZN(n565) );
  NAND2_X1 U510 ( .A1(n550), .A2(n565), .ZN(n457) );
  XOR2_X1 U511 ( .A(n457), .B(KEYINPUT125), .Z(n461) );
  NOR2_X1 U512 ( .A1(n494), .A2(n461), .ZN(n460) );
  INV_X1 U513 ( .A(G218GAT), .ZN(n458) );
  INV_X1 U514 ( .A(n461), .ZN(n589) );
  NAND2_X1 U515 ( .A1(n589), .A2(n466), .ZN(n465) );
  XOR2_X1 U516 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n463) );
  INV_X1 U517 ( .A(G204GAT), .ZN(n462) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n482) );
  OR2_X1 U519 ( .A1(n506), .A2(n466), .ZN(n497) );
  NOR2_X1 U520 ( .A1(n579), .A2(n493), .ZN(n467) );
  XNOR2_X1 U521 ( .A(n467), .B(KEYINPUT16), .ZN(n480) );
  XNOR2_X1 U522 ( .A(n526), .B(KEYINPUT96), .ZN(n468) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n468), .ZN(n471) );
  NAND2_X1 U524 ( .A1(n471), .A2(n523), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT97), .B(n469), .Z(n535) );
  NOR2_X1 U526 ( .A1(n534), .A2(n535), .ZN(n470) );
  XOR2_X1 U527 ( .A(n564), .B(KEYINPUT28), .Z(n530) );
  INV_X1 U528 ( .A(n530), .ZN(n537) );
  NAND2_X1 U529 ( .A1(n470), .A2(n537), .ZN(n479) );
  NAND2_X1 U530 ( .A1(n471), .A2(n550), .ZN(n475) );
  NAND2_X1 U531 ( .A1(n534), .A2(n526), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n564), .A2(n472), .ZN(n473) );
  XOR2_X1 U533 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n477) );
  NAND2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U536 ( .A1(n479), .A2(n478), .ZN(n492) );
  NAND2_X1 U537 ( .A1(n480), .A2(n492), .ZN(n508) );
  NOR2_X1 U538 ( .A1(n497), .A2(n508), .ZN(n489) );
  NAND2_X1 U539 ( .A1(n489), .A2(n523), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n483), .Z(G1324GAT) );
  XOR2_X1 U542 ( .A(G8GAT), .B(KEYINPUT99), .Z(n485) );
  NAND2_X1 U543 ( .A1(n489), .A2(n526), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U546 ( .A1(n489), .A2(n534), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U548 ( .A(G15GAT), .B(n488), .ZN(G1326GAT) );
  XOR2_X1 U549 ( .A(G22GAT), .B(KEYINPUT101), .Z(n491) );
  NAND2_X1 U550 ( .A1(n489), .A2(n530), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(G1327GAT) );
  XOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .Z(n500) );
  NAND2_X1 U553 ( .A1(n493), .A2(n492), .ZN(n495) );
  NOR2_X1 U554 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n496), .B(KEYINPUT37), .ZN(n522) );
  NOR2_X1 U556 ( .A1(n497), .A2(n522), .ZN(n498) );
  XNOR2_X1 U557 ( .A(n498), .B(KEYINPUT38), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n523), .A2(n504), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n504), .A2(n526), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n504), .A2(n534), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  NAND2_X1 U565 ( .A1(n530), .A2(n504), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n505), .ZN(G1331GAT) );
  NAND2_X1 U567 ( .A1(n574), .A2(n506), .ZN(n507) );
  XOR2_X1 U568 ( .A(KEYINPUT103), .B(n507), .Z(n521) );
  NOR2_X1 U569 ( .A1(n508), .A2(n521), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n509), .B(KEYINPUT104), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n517), .A2(n523), .ZN(n513) );
  XOR2_X1 U572 ( .A(KEYINPUT105), .B(KEYINPUT42), .Z(n511) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT106), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U576 ( .A(G64GAT), .B(KEYINPUT107), .Z(n515) );
  NAND2_X1 U577 ( .A1(n517), .A2(n526), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n515), .B(n514), .ZN(G1333GAT) );
  NAND2_X1 U579 ( .A1(n517), .A2(n534), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n530), .A2(n517), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  XOR2_X1 U585 ( .A(G85GAT), .B(KEYINPUT109), .Z(n525) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n531) );
  NAND2_X1 U587 ( .A1(n531), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n531), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U591 ( .A1(n534), .A2(n531), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n528), .B(KEYINPUT110), .ZN(n529) );
  XNOR2_X1 U593 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(KEYINPUT44), .ZN(n533) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  INV_X1 U597 ( .A(n534), .ZN(n569) );
  NOR2_X1 U598 ( .A1(n536), .A2(n535), .ZN(n551) );
  NAND2_X1 U599 ( .A1(n551), .A2(n537), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n569), .A2(n538), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n547), .A2(n586), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(n539), .Z(n540) );
  XNOR2_X1 U603 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n542) );
  NAND2_X1 U605 ( .A1(n547), .A2(n574), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n545) );
  NAND2_X1 U609 ( .A1(n547), .A2(n590), .ZN(n544) );
  XNOR2_X1 U610 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n549) );
  NAND2_X1 U613 ( .A1(n547), .A2(n579), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(G1343GAT) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U616 ( .A(KEYINPUT116), .B(n552), .Z(n560) );
  NAND2_X1 U617 ( .A1(n560), .A2(n586), .ZN(n553) );
  XNOR2_X1 U618 ( .A(n553), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n555) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT117), .B(n556), .Z(n558) );
  NAND2_X1 U623 ( .A1(n560), .A2(n574), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n560), .A2(n590), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .Z(n563) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1347GAT) );
  XNOR2_X1 U630 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n567) );
  AND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n586), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n572) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(n573), .Z(n576) );
  NAND2_X1 U640 ( .A1(n578), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1349GAT) );
  NAND2_X1 U642 ( .A1(n590), .A2(n578), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n583) );
  XNOR2_X1 U645 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT123), .ZN(n581) );
  XNOR2_X1 U647 ( .A(KEYINPUT124), .B(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1351GAT) );
  XNOR2_X1 U649 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n584), .B(KEYINPUT60), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(n585), .Z(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1352GAT) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(G211GAT), .ZN(G1354GAT) );
endmodule

