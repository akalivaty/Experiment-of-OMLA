//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT64), .A2(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT64), .A2(G146), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G143), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n191), .A2(G146), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G146), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n195), .B1(new_n196), .B2(new_n191), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT72), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT67), .B1(new_n201), .B2(G134), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n204), .A3(G137), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(new_n201), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT66), .A2(G137), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT11), .A2(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(G134), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n206), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G131), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT68), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n217), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n206), .A2(new_n211), .A3(new_n214), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT72), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n194), .B(new_n222), .C1(new_n197), .C2(new_n198), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n200), .A2(new_n221), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n190), .A2(new_n225), .A3(G128), .A4(new_n192), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n226), .B1(new_n228), .B2(new_n197), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n206), .A2(new_n211), .A3(new_n216), .A4(new_n214), .ZN(new_n230));
  AOI21_X1  g044(.A(G134), .B1(new_n208), .B2(new_n209), .ZN(new_n231));
  INV_X1    g045(.A(new_n212), .ZN(new_n232));
  OAI21_X1  g046(.A(G131), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT30), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  XOR2_X1   g057(.A(new_n242), .B(new_n243), .Z(new_n244));
  NOR2_X1   g058(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT71), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n233), .A2(new_n230), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n233), .A2(new_n230), .A3(KEYINPUT69), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(new_n229), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  OR2_X1    g066(.A1(new_n199), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n252), .A2(new_n199), .B1(new_n218), .B2(new_n220), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n251), .A2(KEYINPUT70), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n249), .A2(new_n256), .A3(new_n250), .A4(new_n229), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n246), .B(KEYINPUT30), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n251), .A2(KEYINPUT70), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n253), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n259), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT71), .B1(new_n261), .B2(new_n236), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n245), .B1(new_n258), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n224), .A2(new_n244), .A3(new_n234), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT27), .Z(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G101), .ZN(new_n270));
  XOR2_X1   g084(.A(new_n269), .B(new_n270), .Z(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n263), .A2(new_n264), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n265), .B(KEYINPUT28), .ZN(new_n275));
  INV_X1    g089(.A(new_n244), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n261), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n272), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n264), .B1(new_n263), .B2(new_n273), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n187), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT32), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n263), .A2(new_n265), .A3(new_n272), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n271), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT29), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT28), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n244), .B1(new_n224), .B2(new_n234), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT73), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n289), .B1(new_n290), .B2(new_n265), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n266), .A2(KEYINPUT73), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n288), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n266), .A2(KEYINPUT28), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n296));
  AOI21_X1  g110(.A(G902), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G472), .B1(new_n287), .B2(new_n298), .ZN(new_n299));
  OAI211_X1 g113(.A(KEYINPUT32), .B(new_n187), .C1(new_n280), .C2(new_n281), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n284), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  INV_X1    g116(.A(G953), .ZN(new_n303));
  AND4_X1   g117(.A1(G143), .A2(new_n302), .A3(new_n303), .A4(G214), .ZN(new_n304));
  AOI21_X1  g118(.A(G143), .B1(new_n267), .B2(G214), .ZN(new_n305));
  OAI21_X1  g119(.A(G131), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT17), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n302), .A2(new_n303), .A3(G214), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n191), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n267), .A2(G143), .A3(G214), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n216), .A3(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT16), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n313), .A3(G125), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(G146), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n319), .ZN(new_n321));
  INV_X1    g135(.A(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT17), .B(G131), .C1(new_n304), .C2(new_n305), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n312), .A2(new_n320), .A3(new_n323), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT18), .A2(G131), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n309), .A2(new_n310), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n309), .B2(new_n310), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n315), .A2(G140), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n313), .A2(G125), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n196), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT78), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n314), .A2(new_n316), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G146), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n329), .A2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(G113), .B(G122), .ZN(new_n341));
  INV_X1    g155(.A(G104), .ZN(new_n342));
  XNOR2_X1  g156(.A(new_n341), .B(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n325), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT89), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT89), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n325), .A2(new_n340), .A3(new_n346), .A4(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n306), .A2(new_n311), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n320), .A2(KEYINPUT77), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n317), .A2(new_n351), .A3(G146), .A4(new_n319), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT19), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n333), .A2(new_n354), .A3(new_n335), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n337), .A2(KEYINPUT19), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n355), .A2(new_n334), .A3(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n340), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n343), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(KEYINPUT88), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT88), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n362), .A3(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n348), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT90), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n348), .A2(new_n361), .A3(KEYINPUT90), .A4(new_n363), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT20), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT91), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT91), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n372), .A3(KEYINPUT20), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n367), .A2(KEYINPUT92), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n367), .A2(KEYINPUT92), .ZN(new_n375));
  NOR3_X1   g189(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT20), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n371), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n343), .B1(new_n325), .B2(new_n340), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n381), .B1(new_n345), .B2(new_n347), .ZN(new_n382));
  OAI21_X1  g196(.A(G475), .B1(new_n382), .B2(G902), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n303), .A2(G952), .ZN(new_n385));
  INV_X1    g199(.A(G234), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(new_n302), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G902), .ZN(new_n389));
  AOI211_X1 g203(.A(new_n389), .B(new_n303), .C1(G234), .C2(G237), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT21), .B(G898), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n388), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n191), .A2(G128), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n227), .A2(G143), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n393), .A2(new_n394), .A3(new_n204), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n191), .A2(KEYINPUT13), .A3(G128), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n394), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n399), .A2(G134), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n240), .A2(G122), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n240), .A2(G122), .ZN(new_n403));
  OAI21_X1  g217(.A(G107), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n403), .A2(new_n402), .A3(G107), .ZN(new_n405));
  AOI211_X1 g219(.A(new_n395), .B(new_n400), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n204), .B1(new_n393), .B2(new_n394), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n405), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n401), .A2(KEYINPUT14), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n401), .B1(new_n403), .B2(KEYINPUT14), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n409), .B1(new_n410), .B2(KEYINPUT94), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(KEYINPUT94), .B2(new_n410), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n412), .B2(G107), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n406), .A2(new_n413), .A3(KEYINPUT95), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(KEYINPUT9), .B(G234), .Z(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT81), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G217), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n418), .A2(new_n419), .A3(G953), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT95), .B1(new_n406), .B2(new_n413), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n415), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n420), .B1(new_n415), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n389), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G478), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(KEYINPUT15), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  OAI221_X1 g242(.A(new_n389), .B1(KEYINPUT15), .B2(new_n426), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n384), .A2(new_n392), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n419), .B1(G234), .B2(new_n389), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n350), .A2(new_n352), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n227), .A2(G119), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n238), .A2(G128), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT24), .B(G110), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT76), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT76), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT23), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n238), .B2(G128), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n436), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n440), .B(new_n442), .C1(G110), .C2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n434), .A2(new_n447), .A3(new_n336), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT79), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n434), .A2(new_n450), .A3(new_n447), .A4(new_n336), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n323), .A2(new_n320), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT74), .A4(new_n436), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(G110), .A3(new_n456), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n437), .A2(new_n438), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n453), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT75), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n459), .B(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n303), .A2(G221), .A3(G234), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT80), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G137), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n452), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n465), .B1(new_n452), .B2(new_n461), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n389), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT25), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n452), .A2(new_n461), .ZN(new_n471));
  INV_X1    g285(.A(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n452), .A2(new_n461), .A3(new_n465), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT25), .A3(new_n389), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n433), .B1(new_n470), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n432), .A2(G902), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G221), .B1(new_n418), .B2(G902), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n303), .A2(G227), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n482), .B(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(G107), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT82), .A3(G104), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT3), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n485), .A2(G104), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G101), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n491), .A2(new_n485), .A3(KEYINPUT82), .A4(G104), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n489), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n342), .A2(G107), .ZN(new_n494));
  OAI21_X1  g308(.A(G101), .B1(new_n494), .B2(new_n488), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n229), .A3(KEYINPUT10), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n499));
  AOI22_X1  g313(.A1(new_n190), .A2(new_n192), .B1(G128), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n496), .B1(new_n226), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n498), .B1(new_n502), .B2(KEYINPUT10), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n487), .A2(new_n492), .A3(new_n489), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n490), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n487), .A2(new_n489), .A3(KEYINPUT83), .A4(new_n492), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT84), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(KEYINPUT84), .A3(new_n507), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n200), .A2(new_n223), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n506), .B2(new_n508), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n503), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n221), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n484), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n513), .A2(new_n517), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n221), .B1(new_n521), .B2(new_n503), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n497), .A2(new_n229), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n221), .B1(new_n524), .B2(new_n502), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT85), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n226), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n493), .B(new_n495), .C1(new_n528), .C2(new_n500), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n496), .B(new_n226), .C1(new_n197), .C2(new_n228), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n519), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT85), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT12), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT86), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n531), .B2(KEYINPUT12), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n525), .A2(KEYINPUT86), .A3(new_n526), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n534), .A2(new_n538), .B1(new_n519), .B2(new_n518), .ZN(new_n539));
  INV_X1    g353(.A(new_n484), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n523), .B(G469), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(G469), .A2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(G469), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n534), .A2(new_n538), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n546), .A2(new_n520), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n518), .A2(new_n519), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n540), .B1(new_n522), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n545), .B(new_n389), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n481), .B1(new_n544), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G214), .B1(G237), .B2(G902), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n516), .A2(new_n244), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n242), .A2(new_n243), .ZN(new_n555));
  INV_X1    g369(.A(new_n242), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT5), .ZN(new_n557));
  OAI21_X1  g371(.A(G113), .B1(new_n239), .B2(KEYINPUT5), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n513), .A2(new_n554), .B1(new_n497), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(G110), .B(G122), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n561), .B2(new_n562), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OR2_X1    g380(.A1(new_n229), .A2(G125), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n199), .A2(G125), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n303), .A2(G224), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(new_n570), .Z(new_n571));
  OR3_X1    g385(.A1(new_n561), .A2(KEYINPUT6), .A3(new_n562), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n566), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n569), .A2(G224), .A3(new_n303), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n567), .A2(KEYINPUT7), .A3(new_n570), .A4(new_n568), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT7), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n560), .A2(new_n496), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n562), .B(KEYINPUT8), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n557), .A2(KEYINPUT87), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n558), .B1(new_n557), .B2(KEYINPUT87), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n555), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n578), .B(new_n579), .C1(new_n582), .C2(new_n496), .ZN(new_n583));
  AND4_X1   g397(.A1(new_n574), .A2(new_n575), .A3(new_n577), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n561), .A2(new_n562), .ZN(new_n585));
  AOI21_X1  g399(.A(G902), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n573), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(G210), .B1(G237), .B2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n573), .A2(new_n588), .A3(new_n586), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n553), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n551), .A2(new_n592), .ZN(new_n593));
  AND4_X1   g407(.A1(new_n301), .A2(new_n431), .A3(new_n479), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(new_n490), .ZN(G3));
  OAI21_X1  g409(.A(new_n389), .B1(new_n280), .B2(new_n281), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT96), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n598), .B(new_n389), .C1(new_n280), .C2(new_n281), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(G472), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n282), .A2(KEYINPUT97), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n604), .B1(new_n596), .B2(KEYINPUT96), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n605), .A2(new_n606), .A3(new_n599), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT33), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n609), .B1(new_n423), .B2(new_n424), .ZN(new_n610));
  INV_X1    g424(.A(new_n420), .ZN(new_n611));
  INV_X1    g425(.A(new_n421), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n611), .B1(new_n612), .B2(new_n414), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n422), .A3(KEYINPUT33), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n426), .A2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n610), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n425), .A2(new_n426), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n380), .B2(new_n383), .ZN(new_n619));
  INV_X1    g433(.A(new_n392), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n573), .A2(new_n588), .A3(new_n586), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n588), .B1(new_n573), .B2(new_n586), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n552), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AND2_X1   g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n479), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n522), .A2(new_n548), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n627), .A2(new_n484), .B1(new_n546), .B2(new_n520), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n628), .A2(G469), .A3(G902), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n480), .B1(new_n629), .B2(new_n543), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n608), .A2(new_n625), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n342), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT98), .B(KEYINPUT34), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n631), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n603), .B2(new_n607), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n371), .B(new_n373), .C1(KEYINPUT20), .C2(new_n369), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n383), .A3(new_n430), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n623), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT99), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR2_X1   g458(.A1(new_n468), .A2(new_n469), .ZN(new_n645));
  AOI21_X1  g459(.A(KEYINPUT25), .B1(new_n475), .B2(new_n389), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n432), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT101), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT100), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n452), .A2(new_n461), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n649), .B1(new_n452), .B2(new_n461), .ZN(new_n652));
  OAI22_X1  g466(.A1(new_n651), .A2(new_n652), .B1(KEYINPUT36), .B2(new_n465), .ZN(new_n653));
  INV_X1    g467(.A(new_n652), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n465), .A2(KEYINPUT36), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n650), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n653), .A2(new_n656), .A3(new_n478), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n647), .A2(new_n648), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n653), .A2(new_n656), .A3(new_n478), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n477), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n607), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n601), .B1(new_n605), .B2(new_n599), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT102), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n431), .A2(new_n592), .A3(new_n551), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n661), .B1(new_n603), .B2(new_n607), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n666), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT37), .B(G110), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G12));
  NAND4_X1  g487(.A1(new_n551), .A2(new_n592), .A3(new_n660), .A4(new_n658), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n285), .A2(new_n286), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n297), .B1(new_n675), .B2(KEYINPUT29), .ZN(new_n676));
  AOI22_X1  g490(.A1(new_n676), .A2(G472), .B1(new_n282), .B2(new_n283), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n674), .B1(new_n677), .B2(new_n300), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT103), .B(G900), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n390), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n387), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n639), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT104), .B(G128), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G30));
  NAND2_X1  g500(.A1(new_n590), .A2(new_n591), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT38), .Z(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n553), .B1(new_n429), .B2(new_n428), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n384), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n647), .A2(new_n657), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n691), .A2(KEYINPUT105), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n263), .A2(new_n265), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n271), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n291), .A2(new_n272), .A3(new_n292), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n697), .A2(new_n389), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n604), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n282), .B2(new_n283), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n300), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n689), .A2(new_n694), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT105), .B1(new_n691), .B2(new_n693), .ZN(new_n703));
  OR2_X1    g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n681), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n551), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT40), .Z(new_n710));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n616), .A2(new_n617), .ZN(new_n714));
  AND3_X1   g528(.A1(new_n369), .A2(new_n372), .A3(KEYINPUT20), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n372), .B1(new_n369), .B2(KEYINPUT20), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n377), .B(KEYINPUT93), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n383), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n714), .B(new_n681), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n619), .A2(KEYINPUT107), .A3(new_n681), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n678), .A2(new_n713), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n593), .A2(new_n301), .A3(new_n662), .ZN(new_n726));
  OAI21_X1  g540(.A(KEYINPUT108), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G146), .ZN(G48));
  OAI21_X1  g543(.A(G469), .B1(new_n628), .B2(G902), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n550), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n481), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n625), .A2(new_n301), .A3(new_n479), .A4(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT41), .B(G113), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G15));
  NAND4_X1  g549(.A1(new_n640), .A2(new_n732), .A3(new_n301), .A4(new_n479), .ZN(new_n736));
  XNOR2_X1  g550(.A(KEYINPUT109), .B(G116), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G18));
  AND2_X1   g552(.A1(new_n732), .A2(new_n592), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n431), .A2(new_n739), .A3(new_n301), .A4(new_n662), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G119), .ZN(G21));
  AND4_X1   g555(.A1(new_n480), .A2(new_n730), .A3(new_n550), .A4(new_n620), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n687), .A2(new_n742), .A3(new_n384), .A4(new_n690), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n272), .B1(new_n293), .B2(new_n294), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n274), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n187), .B1(new_n745), .B2(new_n281), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n596), .A2(G472), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT110), .B(new_n187), .C1(new_n745), .C2(new_n281), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n479), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n743), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G122), .ZN(G24));
  AND2_X1   g567(.A1(new_n722), .A2(new_n723), .ZN(new_n754));
  AND4_X1   g568(.A1(new_n692), .A2(new_n748), .A3(new_n749), .A4(new_n750), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(KEYINPUT111), .A3(new_n739), .A4(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n722), .A3(new_n723), .A4(new_n739), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  OR2_X1    g575(.A1(new_n300), .A2(KEYINPUT113), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n300), .A2(KEYINPUT113), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n677), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n479), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n630), .A2(new_n687), .A3(new_n553), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT42), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n765), .A2(new_n725), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n301), .A2(new_n766), .A3(new_n479), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n725), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT112), .B(new_n769), .C1(new_n725), .C2(new_n770), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n768), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n216), .ZN(G33));
  INV_X1    g590(.A(new_n770), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n683), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  INV_X1    g593(.A(new_n687), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n552), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n523), .B1(new_n539), .B2(new_n540), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT45), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n545), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n785), .B2(new_n542), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n629), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n785), .A2(KEYINPUT46), .A3(new_n542), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n481), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n708), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n718), .A2(new_n719), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n714), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n603), .A3(new_n607), .A4(new_n692), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n781), .B(new_n790), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  XOR2_X1   g613(.A(new_n789), .B(KEYINPUT47), .Z(new_n800));
  NOR3_X1   g614(.A1(new_n301), .A2(new_n781), .A3(new_n479), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n754), .A2(new_n801), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n794), .A2(new_n388), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n781), .A2(new_n731), .A3(new_n481), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(new_n755), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n701), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n479), .A3(new_n388), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n791), .A2(new_n618), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n806), .A2(new_n751), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n688), .A2(new_n553), .A3(new_n732), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(KEYINPUT50), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n806), .A2(new_n751), .A3(new_n814), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n812), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT116), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n800), .B1(new_n480), .B2(new_n731), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n552), .A3(new_n780), .A4(new_n813), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n819), .B2(KEYINPUT116), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n805), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n824), .B(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n768), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n626), .B1(new_n677), .B2(new_n300), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n722), .A3(new_n723), .A4(new_n766), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT112), .B1(new_n829), .B2(new_n769), .ZN(new_n830));
  INV_X1    g644(.A(new_n774), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n827), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n733), .A2(new_n752), .A3(new_n736), .A4(new_n740), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n755), .A2(new_n722), .A3(new_n723), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n661), .A2(new_n430), .A3(new_n682), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n301), .A3(new_n383), .A4(new_n638), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n833), .B1(new_n766), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n832), .A2(new_n778), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n841));
  AOI211_X1 g655(.A(KEYINPUT102), .B(new_n661), .C1(new_n603), .C2(new_n607), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n667), .A2(new_n828), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n608), .A2(new_n631), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n380), .A2(new_n383), .A3(new_n430), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT114), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n624), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n844), .B(new_n632), .C1(new_n845), .C2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n840), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n594), .B1(new_n625), .B2(new_n637), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n637), .A2(new_n624), .A3(new_n847), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n671), .A2(new_n851), .A3(KEYINPUT115), .A4(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n839), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n756), .A2(new_n759), .B1(new_n683), .B2(new_n678), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n691), .A2(new_n687), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n630), .A2(new_n692), .A3(new_n682), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n701), .A3(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n856), .A3(new_n728), .A4(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n760), .A2(new_n684), .A3(new_n728), .A4(new_n859), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n855), .A2(new_n856), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n854), .A2(new_n860), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n850), .A2(new_n853), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n733), .A2(new_n752), .A3(new_n736), .A4(new_n740), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n837), .A2(new_n766), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n778), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n775), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(new_n873), .A3(new_n860), .A4(new_n862), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n864), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n866), .A2(new_n867), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n863), .A2(KEYINPUT53), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n854), .A2(new_n860), .A3(new_n862), .A4(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n867), .B1(new_n879), .B2(new_n875), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n819), .A2(KEYINPUT51), .A3(new_n822), .ZN(new_n882));
  INV_X1    g696(.A(new_n619), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n385), .B1(new_n810), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n765), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n806), .A2(new_n885), .A3(new_n807), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT48), .Z(new_n887));
  AOI211_X1 g701(.A(new_n884), .B(new_n887), .C1(new_n739), .C2(new_n813), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n826), .A2(new_n881), .A3(new_n882), .A4(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(G952), .B2(G953), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n626), .A2(new_n553), .A3(new_n481), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n731), .A2(KEYINPUT49), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n731), .A2(KEYINPUT49), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  OR4_X1    g708(.A1(new_n689), .A2(new_n894), .A3(new_n701), .A4(new_n792), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n890), .A2(new_n895), .ZN(G75));
  AOI21_X1  g710(.A(new_n389), .B1(new_n866), .B2(new_n875), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(KEYINPUT56), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n566), .A2(new_n572), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT118), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n571), .B(KEYINPUT55), .Z(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n303), .A2(G952), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n906), .B1(new_n898), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n904), .A2(new_n909), .ZN(G51));
  NAND2_X1  g724(.A1(new_n866), .A2(new_n875), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n866), .A2(new_n867), .A3(new_n875), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n542), .B(KEYINPUT57), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(new_n549), .B2(new_n547), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n897), .B(new_n784), .C1(new_n783), .C2(new_n782), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n905), .B1(new_n917), .B2(new_n918), .ZN(G54));
  NAND3_X1  g733(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n366), .A2(new_n368), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n920), .A2(new_n922), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n905), .ZN(G60));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT59), .Z(new_n928));
  AND2_X1   g742(.A1(new_n874), .A2(new_n864), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n874), .A2(new_n877), .ZN(new_n930));
  OAI21_X1  g744(.A(KEYINPUT54), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n928), .B1(new_n931), .B2(new_n913), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n610), .A2(new_n614), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n926), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n928), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n876), .B2(new_n880), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n937), .A2(KEYINPUT120), .A3(new_n933), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n933), .A2(new_n928), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n905), .B1(new_n914), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n935), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT121), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n935), .A2(new_n938), .A3(new_n940), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT60), .Z(new_n947));
  NAND4_X1  g761(.A1(new_n911), .A2(new_n656), .A3(new_n653), .A4(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n911), .A2(new_n947), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n948), .B(new_n906), .C1(new_n475), .C2(new_n949), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT61), .Z(G66));
  INV_X1    g765(.A(new_n391), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n303), .B1(new_n952), .B2(G224), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n868), .A2(new_n869), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n303), .ZN(new_n955));
  INV_X1    g769(.A(G898), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n901), .B1(new_n956), .B2(G953), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  OAI22_X1  g772(.A1(new_n258), .A2(new_n262), .B1(new_n236), .B2(new_n235), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n355), .A2(new_n356), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n798), .A2(new_n803), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n775), .A2(new_n872), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n855), .A2(new_n728), .ZN(new_n966));
  AND4_X1   g780(.A1(new_n708), .A2(new_n885), .A3(new_n857), .A4(new_n789), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT122), .ZN(new_n968));
  NOR4_X1   g782(.A1(new_n963), .A2(new_n965), .A3(new_n966), .A4(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n303), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n303), .A2(G900), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n962), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(G953), .B1(new_n969), .B2(new_n970), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n976), .A2(KEYINPUT124), .A3(new_n973), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n961), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G227), .A2(G900), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(G953), .ZN(new_n980));
  INV_X1    g794(.A(new_n961), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n711), .A2(new_n728), .A3(new_n855), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(KEYINPUT62), .ZN(new_n984));
  OAI211_X1 g798(.A(new_n777), .B(new_n708), .C1(new_n619), .C2(new_n847), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n798), .A2(new_n803), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n981), .B1(new_n988), .B2(G953), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n978), .A2(new_n980), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n972), .A2(new_n962), .A3(new_n974), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT124), .B1(new_n976), .B2(new_n973), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(G953), .B(new_n979), .C1(new_n993), .C2(new_n981), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n990), .A2(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(new_n879), .A2(new_n875), .ZN(new_n996));
  NAND2_X1  g810(.A1(G472), .A2(G902), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT126), .Z(new_n998));
  XOR2_X1   g812(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n996), .A2(new_n285), .A3(new_n696), .A4(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT127), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n987), .B2(new_n954), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n271), .A3(new_n695), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1000), .B1(new_n971), .B2(new_n954), .ZN(new_n1005));
  INV_X1    g819(.A(new_n285), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n905), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(G57));
endmodule


