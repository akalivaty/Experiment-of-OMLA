//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT79), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G155gat), .ZN(new_n207));
  INV_X1    g006(.A(G162gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT79), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n209), .A2(new_n210), .A3(new_n203), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT78), .A2(G148gat), .ZN(new_n213));
  OAI21_X1  g012(.A(G141gat), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n206), .A2(new_n211), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT80), .ZN(new_n218));
  AND3_X1   g017(.A1(new_n203), .A2(new_n218), .A3(KEYINPUT2), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n218), .B1(new_n203), .B2(KEYINPUT2), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G141gat), .B(G148gat), .Z(new_n222));
  NAND2_X1  g021(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n205), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n203), .B(KEYINPUT77), .ZN(new_n225));
  AOI22_X1  g024(.A1(new_n217), .A2(new_n221), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(G127gat), .B(G134gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n228));
  INV_X1    g027(.A(G127gat), .ZN(new_n229));
  OR3_X1    g028(.A1(new_n229), .A2(KEYINPUT68), .A3(G134gat), .ZN(new_n230));
  INV_X1    g029(.A(G113gat), .ZN(new_n231));
  INV_X1    g030(.A(G120gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g033(.A1(G113gat), .A2(G120gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n228), .A2(new_n230), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  NOR2_X1   g038(.A1(G113gat), .A2(G120gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n233), .A2(KEYINPUT69), .A3(new_n235), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n234), .A4(new_n227), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n206), .A2(new_n211), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n214), .A2(new_n216), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n248), .A2(new_n221), .A3(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n223), .ZN(new_n251));
  XNOR2_X1  g050(.A(G141gat), .B(G148gat), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n225), .B(new_n209), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n250), .A2(new_n253), .A3(new_n237), .A4(new_n243), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT4), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n250), .A2(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n250), .A2(new_n259), .A3(new_n253), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n258), .A2(new_n244), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n202), .B1(new_n256), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT39), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n244), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n254), .ZN(new_n265));
  INV_X1    g064(.A(new_n202), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n262), .A2(new_n263), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  AOI211_X1 g068(.A(KEYINPUT39), .B(new_n202), .C1(new_n256), .C2(new_n261), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT0), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G57gat), .ZN(new_n273));
  INV_X1    g072(.A(G85gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n270), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n279));
  AOI21_X1  g078(.A(KEYINPUT84), .B1(new_n279), .B2(new_n275), .ZN(new_n280));
  OAI211_X1 g079(.A(KEYINPUT40), .B(new_n269), .C1(new_n278), .C2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n282), .B1(new_n265), .B2(new_n266), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT81), .B1(new_n254), .B2(KEYINPUT4), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n246), .B1(new_n226), .B2(new_n245), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n202), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n254), .A2(new_n287), .A3(KEYINPUT4), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n261), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n283), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n256), .A2(new_n282), .A3(new_n261), .A4(new_n202), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT86), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT86), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n294), .A3(new_n291), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n276), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  INV_X1    g096(.A(G64gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(G92gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT66), .A2(KEYINPUT25), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n304));
  NOR2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n307), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  OR2_X1    g112(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT65), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n319), .A2(G169gat), .A3(G176gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT66), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n305), .A2(KEYINPUT23), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n316), .A2(new_n321), .A3(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n303), .B1(new_n310), .B2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n321), .A2(new_n324), .ZN(new_n327));
  INV_X1    g126(.A(new_n303), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n316), .A4(new_n309), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT67), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n305), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT26), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n305), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n321), .A3(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT27), .B(G183gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n339), .A2(KEYINPUT28), .A3(new_n312), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT28), .B1(new_n339), .B2(new_n312), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n332), .B(new_n338), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n330), .A2(new_n331), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n330), .A2(new_n343), .B1(new_n346), .B2(new_n331), .ZN(new_n347));
  AND2_X1   g146(.A1(G197gat), .A2(G204gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(G197gat), .A2(G204gat), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(G218gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G211gat), .ZN(new_n352));
  INV_X1    g151(.A(G211gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(G218gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(G211gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n357), .A2(new_n359), .A3(G218gat), .ZN(new_n360));
  AOI211_X1 g159(.A(new_n350), .B(new_n355), .C1(new_n356), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n355), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n356), .ZN(new_n363));
  INV_X1    g162(.A(new_n350), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n345), .A2(new_n347), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n361), .B2(new_n365), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT73), .B(G211gat), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT22), .B1(new_n371), .B2(G218gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n355), .B1(new_n372), .B2(new_n350), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n363), .A2(new_n364), .A3(new_n362), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(KEYINPUT74), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n330), .A2(new_n343), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n331), .A2(new_n346), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n376), .B1(new_n379), .B2(new_n344), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n302), .B1(new_n368), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT76), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n376), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n345), .B2(new_n347), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n366), .A3(new_n344), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n301), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT30), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(KEYINPUT30), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n385), .A2(new_n386), .A3(new_n301), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n281), .B(new_n296), .C1(new_n389), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT87), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n269), .B1(new_n278), .B2(new_n280), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT85), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT40), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n277), .B1(new_n270), .B2(new_n276), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n279), .A2(KEYINPUT84), .A3(new_n275), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n268), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT85), .B1(new_n402), .B2(KEYINPUT40), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n394), .A2(new_n395), .A3(new_n399), .A4(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n367), .B1(new_n345), .B2(new_n347), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n379), .A2(new_n376), .A3(new_n344), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT37), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT37), .B1(new_n385), .B2(new_n386), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n408), .B2(KEYINPUT88), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT38), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT88), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n405), .A2(new_n406), .A3(new_n411), .A4(KEYINPUT37), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n409), .A2(new_n410), .A3(new_n301), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n383), .A2(new_n388), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT37), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n301), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT38), .B1(new_n416), .B2(new_n408), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n290), .A2(new_n275), .A3(new_n291), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT6), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n275), .B1(new_n290), .B2(new_n291), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n296), .A2(new_n422), .B1(KEYINPUT6), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G228gat), .ZN(new_n425));
  INV_X1    g224(.A(G233gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n346), .B1(new_n361), .B2(new_n365), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n259), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n257), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n260), .A2(new_n346), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n366), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n427), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n375), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT74), .B1(new_n373), .B2(new_n374), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT82), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n430), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n370), .A2(new_n375), .B1(new_n260), .B2(new_n346), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n427), .B1(new_n440), .B2(KEYINPUT82), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n439), .A2(new_n441), .A3(KEYINPUT83), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  INV_X1    g242(.A(new_n427), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n444), .B1(new_n437), .B2(new_n438), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n440), .A2(KEYINPUT82), .B1(new_n257), .B2(new_n429), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n434), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G22gat), .B(G78gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(KEYINPUT31), .B(G50gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G106gat), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT83), .B1(new_n439), .B2(new_n441), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n445), .A2(new_n446), .A3(new_n443), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(new_n449), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(new_n456), .A3(new_n434), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n452), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n455), .B2(new_n434), .ZN(new_n460));
  AOI211_X1 g259(.A(new_n449), .B(new_n433), .C1(new_n453), .C2(new_n454), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n418), .A2(new_n424), .B1(new_n458), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n399), .A2(new_n403), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT87), .B1(new_n464), .B2(new_n393), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n404), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n392), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n421), .A2(new_n423), .ZN(new_n469));
  AOI211_X1 g268(.A(new_n420), .B(new_n275), .C1(new_n290), .C2(new_n291), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT30), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n473));
  AOI211_X1 g272(.A(new_n382), .B(new_n301), .C1(new_n385), .C2(new_n386), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n467), .B2(new_n392), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n458), .B(new_n462), .C1(new_n471), .C2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n377), .A2(new_n245), .ZN(new_n479));
  INV_X1    g278(.A(G227gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n426), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n330), .A2(new_n244), .A3(new_n343), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(KEYINPUT71), .B(G71gat), .ZN(new_n487));
  INV_X1    g286(.A(G99gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G15gat), .B(G43gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n330), .A2(new_n244), .A3(new_n343), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n244), .B1(new_n330), .B2(new_n343), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT34), .B1(new_n495), .B2(new_n481), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n482), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT34), .ZN(new_n498));
  INV_X1    g297(.A(new_n481), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n483), .A2(KEYINPUT32), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n501), .B1(new_n496), .B2(new_n500), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n492), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n483), .A2(KEYINPUT32), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n506));
  AOI211_X1 g305(.A(KEYINPUT34), .B(new_n481), .C1(new_n479), .C2(new_n482), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n492), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n496), .A2(new_n500), .A3(new_n501), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n478), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  NOR3_X1   g311(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT72), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT36), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n504), .A2(new_n511), .ZN(new_n515));
  OR2_X1    g314(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n477), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n466), .A2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT72), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n513), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n460), .A2(new_n461), .A3(new_n459), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n452), .B1(new_n450), .B2(new_n457), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n521), .B(new_n522), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n392), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n389), .B1(KEYINPUT75), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n421), .B(new_n423), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(new_n468), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT35), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n515), .B1(new_n462), .B2(new_n458), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n526), .A2(new_n475), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n424), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT94), .ZN(new_n538));
  XNOR2_X1  g337(.A(G43gat), .B(G50gat), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n539), .A2(KEYINPUT89), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(KEYINPUT89), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(KEYINPUT15), .A3(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(KEYINPUT90), .B(G36gat), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(G29gat), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT14), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  OR3_X1    g345(.A1(new_n545), .A2(G29gat), .A3(G36gat), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n544), .A2(KEYINPUT91), .A3(new_n546), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n542), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n551));
  NOR3_X1   g350(.A1(new_n551), .A2(KEYINPUT15), .A3(new_n539), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G8gat), .ZN(new_n555));
  XOR2_X1   g354(.A(G15gat), .B(G22gat), .Z(new_n556));
  INV_X1    g355(.A(G1gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n555), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n557), .A2(KEYINPUT16), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n558), .B1(new_n556), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n560), .B(new_n562), .Z(new_n563));
  OR2_X1    g362(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  OR3_X1    g363(.A1(new_n549), .A2(KEYINPUT17), .A3(new_n552), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT17), .B1(new_n549), .B2(new_n552), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n563), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT18), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n554), .B(new_n563), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n568), .B(KEYINPUT93), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT13), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n564), .A2(new_n567), .A3(KEYINPUT18), .A4(new_n568), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G113gat), .B(G141gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(G197gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT11), .ZN(new_n580));
  INV_X1    g379(.A(G169gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT12), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n577), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n571), .A2(new_n583), .A3(new_n575), .A4(new_n576), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n537), .A2(new_n538), .A3(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n466), .A2(new_n517), .B1(new_n530), .B2(new_n535), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT94), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT9), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595));
  NAND2_X1  g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n594), .A2(new_n595), .A3(new_n596), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n298), .A2(G57gat), .ZN(new_n600));
  XOR2_X1   g399(.A(KEYINPUT96), .B(G57gat), .Z(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(new_n298), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n596), .B1(new_n598), .B2(new_n593), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n596), .B1(new_n592), .B2(new_n593), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT95), .B1(new_n605), .B2(new_n597), .ZN(new_n606));
  AND3_X1   g405(.A1(new_n599), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n563), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT98), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT99), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(new_n229), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n613), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT97), .B(G155gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G183gat), .B(G211gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n618), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT7), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  NAND2_X1  g425(.A1(G99gat), .A2(G106gat), .ZN(new_n627));
  AOI22_X1  g426(.A1(KEYINPUT8), .A2(new_n627), .B1(new_n274), .B2(new_n300), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n626), .B1(new_n625), .B2(new_n628), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT101), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n565), .A2(new_n566), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT102), .ZN(new_n636));
  NAND2_X1  g435(.A1(G232gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT100), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n635), .A2(new_n636), .B1(KEYINPUT41), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n554), .A2(new_n634), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT102), .A4(new_n634), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n640), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G190gat), .B(G218gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(KEYINPUT103), .B(G134gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n639), .A2(KEYINPUT41), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(new_n208), .ZN(new_n649));
  INV_X1    g448(.A(new_n646), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n640), .A2(new_n650), .A3(new_n641), .A4(new_n642), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n649), .B1(new_n647), .B2(new_n651), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n623), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n629), .A2(new_n630), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n607), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n599), .A2(new_n604), .A3(new_n606), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n632), .B2(new_n633), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT104), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n659), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  INV_X1    g465(.A(G176gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(G204gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n663), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT10), .B1(new_n659), .B2(new_n661), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n634), .A2(new_n673), .A3(new_n660), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n671), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT105), .B(new_n671), .C1(new_n672), .C2(new_n674), .ZN(new_n678));
  AOI211_X1 g477(.A(new_n665), .B(new_n670), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n675), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n670), .B1(new_n681), .B2(new_n665), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n588), .A2(new_n591), .A3(new_n656), .A4(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n528), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT106), .B(G1gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1324gat));
  NOR2_X1   g486(.A1(new_n389), .A2(new_n392), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT16), .B(G8gat), .Z(new_n690));
  AOI21_X1  g489(.A(KEYINPUT107), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT42), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n555), .B2(new_n689), .ZN(G1325gat));
  INV_X1    g492(.A(G15gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n514), .A2(new_n516), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n684), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n684), .A2(new_n515), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n694), .B2(new_n698), .ZN(G1326gat));
  INV_X1    g498(.A(G22gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n462), .A2(new_n458), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n684), .A2(KEYINPUT108), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT108), .B1(new_n684), .B2(new_n701), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n700), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n709), .A2(G22gat), .A3(new_n705), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n708), .A2(new_n710), .ZN(G1327gat));
  NAND3_X1  g510(.A1(new_n588), .A2(new_n591), .A3(new_n683), .ZN(new_n712));
  INV_X1    g511(.A(new_n655), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n712), .A2(new_n622), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n528), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717));
  INV_X1    g516(.A(G29gat), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n717), .B1(new_n716), .B2(new_n718), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n471), .A2(new_n476), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n513), .B1(new_n515), .B2(KEYINPUT72), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n701), .ZN(new_n723));
  AOI221_X4 g522(.A(KEYINPUT111), .B1(new_n531), .B2(new_n534), .C1(new_n723), .C2(KEYINPUT35), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT111), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n530), .B2(new_n535), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n518), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n728), .A3(new_n655), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n713), .B1(new_n518), .B2(new_n536), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT110), .B1(new_n730), .B2(new_n728), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n732), .B(KEYINPUT44), .C1(new_n589), .C2(new_n713), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n729), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n622), .B(KEYINPUT109), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n590), .ZN(new_n736));
  AND4_X1   g535(.A1(new_n715), .A2(new_n734), .A3(new_n683), .A4(new_n736), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n719), .A2(new_n720), .B1(new_n718), .B2(new_n737), .ZN(G1328gat));
  INV_X1    g537(.A(new_n543), .ZN(new_n739));
  INV_X1    g538(.A(new_n688), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n714), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(KEYINPUT46), .ZN(new_n743));
  AND4_X1   g542(.A1(new_n683), .A2(new_n734), .A3(new_n740), .A4(new_n736), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(new_n743), .C1(new_n739), .C2(new_n744), .ZN(G1329gat));
  INV_X1    g544(.A(G43gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n515), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n714), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  AND4_X1   g547(.A1(new_n683), .A2(new_n734), .A3(new_n695), .A4(new_n736), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n746), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1330gat));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n753));
  INV_X1    g552(.A(new_n701), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n734), .A2(new_n683), .A3(new_n754), .A4(new_n736), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  INV_X1    g555(.A(G50gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n714), .A2(new_n757), .A3(new_n754), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n753), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1331gat));
  AND3_X1   g560(.A1(new_n727), .A2(new_n656), .A3(new_n590), .ZN(new_n762));
  INV_X1    g561(.A(new_n683), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR3_X1    g563(.A1(new_n764), .A2(KEYINPUT113), .A3(new_n528), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT113), .B1(new_n764), .B2(new_n528), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n601), .ZN(G1332gat));
  NOR2_X1   g567(.A1(new_n764), .A2(new_n688), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n764), .B2(new_n515), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n762), .A2(G71gat), .A3(new_n763), .A4(new_n695), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n776), .B2(new_n778), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n774), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n781), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n783), .A2(KEYINPUT50), .A3(new_n779), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1334gat));
  NOR2_X1   g584(.A1(new_n764), .A2(new_n701), .ZN(new_n786));
  XOR2_X1   g585(.A(new_n786), .B(G78gat), .Z(G1335gat));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n622), .A2(new_n683), .A3(new_n587), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n734), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n788), .B1(new_n734), .B2(new_n789), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n715), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g593(.A(KEYINPUT116), .B(new_n715), .C1(new_n790), .C2(new_n791), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(G85gat), .A3(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n727), .A2(new_n623), .A3(new_n655), .A4(new_n590), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT51), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n799), .A2(new_n274), .A3(new_n715), .A4(new_n763), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n796), .A2(new_n800), .ZN(G1336gat));
  NAND2_X1  g600(.A1(new_n734), .A2(new_n789), .ZN(new_n802));
  OAI21_X1  g601(.A(G92gat), .B1(new_n802), .B2(new_n688), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n683), .A2(G92gat), .A3(new_n688), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n803), .B(new_n804), .C1(new_n798), .C2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n740), .B1(new_n790), .B2(new_n791), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT51), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n797), .B(new_n810), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n808), .A2(G92gat), .B1(new_n811), .B2(new_n805), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n807), .B1(new_n812), .B2(new_n804), .ZN(G1337gat));
  NOR2_X1   g612(.A1(new_n790), .A2(new_n791), .ZN(new_n814));
  OAI21_X1  g613(.A(G99gat), .B1(new_n814), .B2(new_n696), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n488), .A3(new_n747), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n815), .B1(new_n683), .B2(new_n816), .ZN(G1338gat));
  OAI21_X1  g616(.A(G106gat), .B1(new_n802), .B2(new_n701), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n683), .A2(new_n701), .A3(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n818), .B(new_n819), .C1(new_n798), .C2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n754), .B1(new_n790), .B2(new_n791), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n823), .A2(G106gat), .B1(new_n811), .B2(new_n820), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n824), .B2(new_n819), .ZN(G1339gat));
  NOR2_X1   g624(.A1(new_n572), .A2(new_n574), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n568), .B1(new_n564), .B2(new_n567), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n582), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n586), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n653), .A2(new_n654), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n672), .A2(new_n674), .A3(new_n671), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n831), .B(new_n832), .C1(new_n677), .C2(new_n678), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n670), .B1(new_n675), .B2(KEYINPUT54), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT55), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n832), .B1(new_n677), .B2(new_n678), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  INV_X1    g636(.A(new_n834), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n835), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT118), .B1(new_n841), .B2(new_n680), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(new_n679), .C1(new_n835), .C2(new_n840), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n830), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n833), .A2(KEYINPUT55), .A3(new_n834), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n839), .B1(new_n837), .B2(new_n838), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n680), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(new_n843), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n841), .A2(KEYINPUT118), .A3(new_n680), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n852), .A2(new_n853), .A3(new_n830), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n587), .B1(new_n842), .B2(new_n844), .ZN(new_n856));
  INV_X1    g655(.A(new_n829), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n763), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n713), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n735), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n623), .A2(new_n655), .A3(new_n763), .A4(new_n587), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR3_X1   g662(.A1(new_n863), .A2(new_n528), .A3(new_n740), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n531), .ZN(new_n865));
  OAI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n590), .ZN(new_n866));
  INV_X1    g665(.A(new_n525), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n587), .A2(new_n231), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n865), .B2(new_n683), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n763), .A2(new_n232), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n871), .B1(new_n868), .B2(new_n872), .ZN(G1341gat));
  INV_X1    g672(.A(new_n735), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n865), .A2(new_n229), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n864), .A2(new_n622), .A3(new_n867), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n229), .B2(new_n876), .ZN(G1342gat));
  NAND2_X1  g676(.A1(new_n655), .A2(new_n688), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT120), .Z(new_n879));
  OR3_X1    g678(.A1(new_n863), .A2(new_n528), .A3(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(G134gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n867), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n884));
  OAI21_X1  g683(.A(G134gat), .B1(new_n865), .B2(new_n713), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n881), .A2(new_n886), .A3(new_n882), .A4(new_n867), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(G1343gat));
  OAI21_X1  g687(.A(new_n858), .B1(new_n849), .B2(new_n590), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n713), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n845), .A2(KEYINPUT119), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n853), .B1(new_n852), .B2(new_n830), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n862), .B1(new_n893), .B2(new_n623), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n701), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n695), .A2(new_n528), .A3(new_n740), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n897), .B(new_n754), .C1(new_n861), .C2(new_n862), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n895), .A2(new_n587), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n863), .A2(new_n701), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n901), .A2(new_n215), .A3(new_n587), .A4(new_n896), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT58), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT58), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n900), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1344gat));
  NOR2_X1   g706(.A1(new_n212), .A2(new_n213), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n683), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n901), .A2(new_n896), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT57), .B1(new_n863), .B2(new_n701), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n830), .A2(new_n680), .A3(new_n841), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n622), .B1(new_n890), .B2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n897), .B(new_n754), .C1(new_n862), .C2(new_n914), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n896), .B(KEYINPUT121), .Z(new_n916));
  NAND4_X1  g715(.A1(new_n912), .A2(new_n763), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n911), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n895), .A2(new_n763), .A3(new_n896), .A4(new_n898), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n919), .A2(new_n911), .A3(new_n908), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n910), .B1(new_n918), .B2(new_n920), .ZN(G1345gat));
  NAND3_X1  g720(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n207), .A3(new_n874), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n901), .A2(new_n622), .A3(new_n896), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT122), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT122), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n901), .A2(new_n926), .A3(new_n622), .A4(new_n896), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n923), .B1(new_n928), .B2(new_n207), .ZN(G1346gat));
  OAI21_X1  g728(.A(G162gat), .B1(new_n922), .B2(new_n713), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT123), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n880), .A2(G162gat), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n695), .A2(new_n701), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n933), .ZN(new_n935));
  NOR4_X1   g734(.A1(new_n880), .A2(KEYINPUT123), .A3(G162gat), .A4(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n930), .B1(new_n934), .B2(new_n936), .ZN(G1347gat));
  NOR2_X1   g736(.A1(new_n715), .A2(new_n688), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n531), .B(new_n938), .C1(new_n861), .C2(new_n862), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n590), .ZN(new_n940));
  INV_X1    g739(.A(new_n938), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n855), .A2(new_n860), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n874), .ZN(new_n943));
  INV_X1    g742(.A(new_n862), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(new_n867), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n587), .A2(new_n581), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(G1348gat));
  NOR3_X1   g747(.A1(new_n939), .A2(new_n667), .A3(new_n683), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n763), .A3(new_n867), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n667), .B2(new_n950), .ZN(G1349gat));
  NAND4_X1  g750(.A1(new_n945), .A2(KEYINPUT124), .A3(new_n531), .A4(new_n735), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT124), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n953), .B1(new_n939), .B2(new_n874), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(new_n954), .A3(G183gat), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n945), .A2(new_n622), .A3(new_n339), .A4(new_n867), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(KEYINPUT60), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT60), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n959), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n939), .B2(new_n713), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT125), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n965), .B(G190gat), .C1(new_n939), .C2(new_n713), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n963), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n964), .B1(new_n963), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n655), .A2(new_n312), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n946), .B2(new_n969), .ZN(G1351gat));
  AND2_X1   g769(.A1(new_n912), .A2(new_n915), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n696), .A2(new_n938), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n971), .A2(new_n587), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n975), .A2(G197gat), .ZN(new_n976));
  OAI211_X1 g775(.A(new_n933), .B(new_n938), .C1(new_n861), .C2(new_n862), .ZN(new_n977));
  OR3_X1    g776(.A1(new_n977), .A2(G197gat), .A3(new_n590), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n976), .A2(new_n978), .ZN(G1352gat));
  NAND4_X1  g778(.A1(new_n912), .A2(new_n763), .A3(new_n915), .A4(new_n974), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G204gat), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n943), .A2(new_n944), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n982), .A2(new_n669), .A3(new_n933), .A4(new_n938), .ZN(new_n983));
  OAI21_X1  g782(.A(KEYINPUT127), .B1(new_n983), .B2(new_n683), .ZN(new_n984));
  INV_X1    g783(.A(new_n977), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  NAND4_X1  g785(.A1(new_n985), .A2(new_n986), .A3(new_n669), .A4(new_n763), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n984), .B2(new_n987), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n981), .B1(new_n989), .B2(new_n990), .ZN(G1353gat));
  OR3_X1    g790(.A1(new_n977), .A2(new_n623), .A3(new_n371), .ZN(new_n992));
  NAND4_X1  g791(.A1(new_n912), .A2(new_n622), .A3(new_n915), .A4(new_n974), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  AOI21_X1  g795(.A(G218gat), .B1(new_n985), .B2(new_n655), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n971), .A2(new_n974), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n713), .A2(new_n351), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(G1355gat));
endmodule


