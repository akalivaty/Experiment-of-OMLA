//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  OAI211_X1 g006(.A(new_n187), .B(new_n192), .C1(new_n188), .C2(G137), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G137), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n190), .A2(new_n191), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT67), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n188), .B2(G137), .ZN(new_n197));
  INV_X1    g011(.A(G137), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n198), .A2(KEYINPUT67), .A3(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n197), .A2(new_n194), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G131), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(KEYINPUT65), .A2(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(G143), .A3(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n204), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(KEYINPUT1), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n207), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n207), .B2(KEYINPUT1), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n214), .A2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n205), .A2(new_n206), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(new_n214), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n212), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n202), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(KEYINPUT65), .A2(G146), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT65), .A2(G146), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n215), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g038(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n220), .A2(new_n221), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n208), .B1(new_n230), .B2(G143), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n195), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n198), .A2(G134), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n189), .B2(KEYINPUT11), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n191), .B1(new_n237), .B2(new_n193), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n229), .B(new_n234), .C1(new_n235), .C2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G119), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(G116), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G119), .ZN(new_n247));
  INV_X1    g061(.A(G113), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT2), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT2), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G113), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n245), .A2(new_n247), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n245), .B2(new_n247), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n240), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n245), .A2(new_n247), .ZN(new_n256));
  INV_X1    g070(.A(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n245), .A2(new_n247), .A3(new_n252), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n219), .A2(new_n239), .A3(new_n255), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT73), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n261), .A2(new_n265), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT29), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  INV_X1    g083(.A(G237), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(KEYINPUT71), .A2(G237), .ZN(new_n272));
  AOI21_X1  g086(.A(G953), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G210), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT27), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT26), .B(G101), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n267), .A2(new_n268), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(KEYINPUT66), .B1(new_n198), .B2(G134), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n194), .B1(new_n280), .B2(new_n192), .ZN(new_n281));
  INV_X1    g095(.A(new_n193), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n195), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n231), .A2(new_n233), .B1(new_n224), .B2(new_n228), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n284), .B2(new_n285), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n219), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n255), .A2(new_n260), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n255), .A2(new_n260), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n292), .B(new_n219), .C1(new_n287), .C2(new_n288), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n289), .A2(new_n295), .A3(new_n290), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n294), .A2(KEYINPUT28), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n279), .B2(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n284), .A2(new_n285), .B1(new_n202), .B2(new_n218), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT72), .B1(new_n299), .B2(new_n292), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n219), .A2(new_n239), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n290), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n293), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT28), .ZN(new_n305));
  AOI211_X1 g119(.A(KEYINPUT73), .B(KEYINPUT28), .C1(new_n299), .C2(new_n292), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n265), .B1(new_n261), .B2(new_n262), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n305), .A2(new_n277), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT74), .ZN(new_n310));
  OAI211_X1 g124(.A(KEYINPUT30), .B(new_n219), .C1(new_n287), .C2(new_n288), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT30), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n292), .B1(new_n301), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n219), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n239), .A2(KEYINPUT70), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n311), .A2(new_n313), .B1(new_n317), .B2(new_n292), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n310), .B1(new_n318), .B2(new_n277), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n293), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n278), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n309), .A2(new_n319), .A3(new_n322), .A4(new_n268), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n298), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G472), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n277), .B1(new_n305), .B2(new_n308), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT31), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n327), .B1(new_n318), .B2(new_n277), .ZN(new_n328));
  AND4_X1   g142(.A1(new_n327), .A2(new_n320), .A3(new_n277), .A4(new_n293), .ZN(new_n329));
  NOR3_X1   g143(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G472), .A2(G902), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n330), .A2(KEYINPUT32), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT32), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n318), .A2(new_n277), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT31), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n318), .A2(new_n327), .A3(new_n277), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n267), .B1(KEYINPUT28), .B2(new_n304), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n277), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n339), .B2(new_n331), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n325), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G140), .ZN(new_n342));
  INV_X1    g156(.A(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G227), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n342), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(new_n284), .ZN(new_n346));
  INV_X1    g160(.A(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G107), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT81), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n347), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n347), .A3(G107), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n353));
  INV_X1    g167(.A(G107), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(G104), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n349), .A2(new_n350), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G101), .ZN(new_n357));
  NOR2_X1   g171(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n354), .A2(G104), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G101), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n347), .A2(G107), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n358), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n363), .A2(new_n364), .A3(new_n348), .A4(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n357), .A2(new_n367), .A3(KEYINPUT10), .ZN(new_n368));
  INV_X1    g182(.A(new_n212), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n207), .A2(new_n209), .B1(G128), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n357), .B(new_n367), .C1(new_n369), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n218), .A2(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n348), .B1(new_n359), .B2(new_n362), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n358), .B1(new_n365), .B2(new_n360), .ZN(new_n376));
  OAI21_X1  g190(.A(G101), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n367), .A3(KEYINPUT4), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT4), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G101), .C1(new_n375), .C2(new_n376), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n285), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n346), .B1(new_n374), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n368), .A2(new_n218), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n372), .A2(new_n373), .ZN(new_n384));
  AND4_X1   g198(.A1(new_n346), .A2(new_n383), .A3(new_n384), .A4(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n345), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n345), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n383), .A2(new_n384), .A3(new_n381), .A4(new_n346), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n357), .A2(new_n367), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n372), .B1(new_n389), .B2(new_n218), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n390), .A2(KEYINPUT12), .A3(new_n284), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT12), .B1(new_n390), .B2(new_n284), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n387), .B(new_n388), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n386), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G469), .ZN(new_n395));
  INV_X1    g209(.A(G902), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n388), .A2(new_n387), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT82), .ZN(new_n399));
  INV_X1    g213(.A(new_n382), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n388), .A2(new_n401), .A3(new_n387), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n345), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n405), .A3(G469), .ZN(new_n406));
  NAND2_X1  g220(.A1(G469), .A2(G902), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT9), .B(G234), .ZN(new_n409));
  OAI21_X1  g223(.A(G221), .B1(new_n409), .B2(G902), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n408), .A2(KEYINPUT83), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(KEYINPUT83), .B1(new_n408), .B2(new_n410), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  INV_X1    g229(.A(G122), .ZN(new_n416));
  NOR3_X1   g230(.A1(new_n416), .A2(KEYINPUT14), .A3(G116), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT93), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n354), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT14), .B1(new_n416), .B2(G116), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(new_n246), .A3(G122), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n416), .A2(G116), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT93), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n246), .A2(G122), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(new_n423), .A3(new_n354), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n214), .A2(G128), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n210), .A2(G143), .ZN(new_n429));
  OAI21_X1  g243(.A(G134), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n210), .A2(G143), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n214), .A2(G128), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n188), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n425), .A2(new_n427), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n214), .A2(KEYINPUT13), .A3(G128), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT91), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT13), .B1(new_n214), .B2(G128), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n437), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT91), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n440), .A3(new_n432), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G134), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n433), .A2(KEYINPUT92), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n431), .A2(new_n432), .A3(new_n445), .A4(new_n188), .ZN(new_n446));
  INV_X1    g260(.A(new_n427), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n354), .B1(new_n426), .B2(new_n423), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n444), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n435), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT76), .B(G217), .Z(new_n451));
  NOR3_X1   g265(.A1(new_n451), .A2(G953), .A3(new_n409), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n429), .B1(KEYINPUT13), .B2(new_n431), .ZN(new_n455));
  OAI211_X1 g269(.A(G134), .B(new_n441), .C1(new_n455), .C2(new_n437), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n426), .A2(new_n423), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G107), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n427), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n456), .A2(new_n446), .A3(new_n459), .A4(new_n444), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n452), .B1(new_n460), .B2(new_n435), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n396), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT94), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n450), .A2(new_n453), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n460), .A2(new_n435), .A3(new_n452), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n415), .B1(new_n463), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(KEYINPUT94), .B(G902), .C1(new_n464), .C2(new_n465), .ZN(new_n470));
  INV_X1    g284(.A(new_n415), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n469), .A2(KEYINPUT95), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT95), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n464), .A2(new_n465), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n467), .B1(new_n475), .B2(new_n396), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n471), .B1(new_n476), .B2(new_n470), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n415), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g294(.A1(G475), .A2(G902), .ZN(new_n481));
  XNOR2_X1  g295(.A(G113), .B(G122), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(new_n347), .ZN(new_n483));
  AOI21_X1  g297(.A(G143), .B1(new_n273), .B2(G214), .ZN(new_n484));
  AND2_X1   g298(.A1(G143), .A2(G214), .ZN(new_n485));
  AND2_X1   g299(.A1(KEYINPUT71), .A2(G237), .ZN(new_n486));
  NOR2_X1   g300(.A1(KEYINPUT71), .A2(G237), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n343), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n191), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n484), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n343), .B1(new_n486), .B2(new_n487), .ZN(new_n494));
  INV_X1    g308(.A(G214), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n214), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(KEYINPUT88), .A3(new_n191), .A4(new_n488), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n490), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT89), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n490), .A2(new_n493), .A3(KEYINPUT89), .A4(new_n497), .ZN(new_n501));
  INV_X1    g315(.A(G140), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(G125), .ZN(new_n503));
  INV_X1    g317(.A(G125), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G140), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT87), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT87), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n509), .A3(KEYINPUT19), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(KEYINPUT77), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT19), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n503), .A2(new_n505), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n510), .A2(new_n515), .A3(new_n230), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n502), .A3(G125), .ZN(new_n518));
  OAI211_X1 g332(.A(G146), .B(new_n518), .C1(new_n506), .C2(new_n517), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n500), .A2(new_n501), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n496), .A2(new_n488), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT18), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n523), .B1(new_n524), .B2(new_n191), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n496), .A2(KEYINPUT18), .A3(G131), .A4(new_n488), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n507), .A2(G146), .A3(new_n509), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n511), .A2(new_n230), .A3(new_n514), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n483), .B1(new_n522), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n518), .B1(new_n506), .B2(new_n517), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n204), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n519), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT17), .B(G131), .C1(new_n484), .C2(new_n489), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT90), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n490), .A2(new_n493), .A3(new_n539), .A4(new_n497), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n523), .A2(KEYINPUT90), .A3(KEYINPUT17), .A4(G131), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n542), .A2(new_n483), .A3(new_n531), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n481), .B1(new_n532), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT20), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(new_n481), .C1(new_n532), .C2(new_n543), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n483), .B1(new_n542), .B2(new_n531), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n396), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n545), .A2(new_n547), .B1(G475), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g364(.A1(new_n343), .A2(G952), .ZN(new_n551));
  NAND2_X1  g365(.A1(G234), .A2(G237), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n552), .A2(G902), .A3(G953), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT21), .B(G898), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n554), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n480), .A2(new_n550), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G214), .B1(G237), .B2(G902), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT84), .ZN(new_n562));
  OAI21_X1  g376(.A(G210), .B1(G237), .B2(G902), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n504), .B(new_n212), .C1(new_n213), .C2(new_n217), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n285), .B2(new_n504), .ZN(new_n566));
  INV_X1    g380(.A(G224), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  XOR2_X1   g382(.A(new_n566), .B(new_n568), .Z(new_n569));
  OAI21_X1  g383(.A(KEYINPUT85), .B1(new_n245), .B2(KEYINPUT5), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n245), .A2(KEYINPUT5), .A3(new_n247), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT68), .B(G119), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT85), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT5), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(G116), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n570), .A2(new_n571), .A3(G113), .A4(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n389), .A2(new_n259), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(G110), .B(G122), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n378), .A2(new_n380), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n577), .B(new_n578), .C1(new_n292), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT6), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n577), .B1(new_n292), .B2(new_n579), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n578), .A2(KEYINPUT86), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n583), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n569), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n578), .B(KEYINPUT8), .ZN(new_n588));
  INV_X1    g402(.A(new_n577), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n389), .B1(new_n259), .B2(new_n576), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT7), .ZN(new_n592));
  OR3_X1    g406(.A1(new_n566), .A2(new_n592), .A3(new_n568), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n566), .B1(new_n592), .B2(new_n568), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n591), .A2(new_n593), .A3(new_n580), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n396), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n564), .B1(new_n587), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n569), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n580), .A2(KEYINPUT6), .B1(new_n582), .B2(new_n583), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n582), .A2(KEYINPUT6), .A3(new_n583), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(new_n396), .A3(new_n563), .A4(new_n595), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n562), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n560), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n451), .B1(G234), .B2(new_n396), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT23), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n572), .B2(G128), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n241), .A2(new_n210), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n572), .B2(new_n210), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n609), .B1(new_n611), .B2(new_n608), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT24), .B(G110), .Z(new_n613));
  OAI22_X1  g427(.A1(new_n612), .A2(G110), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n519), .A3(new_n529), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(G110), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n613), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n616), .A2(new_n617), .A3(new_n535), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT22), .B(G137), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n343), .A2(G221), .A3(G234), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT78), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n615), .A2(new_n618), .A3(new_n622), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n624), .A2(new_n625), .A3(new_n396), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT25), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n624), .A2(new_n625), .A3(KEYINPUT25), .A4(new_n396), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n607), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n625), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n606), .A2(G902), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n341), .A2(new_n413), .A3(new_n605), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  INV_X1    g450(.A(G472), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(new_n339), .B2(new_n396), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n330), .A2(new_n332), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n413), .A2(new_n640), .A3(new_n634), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n561), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n597), .B2(new_n602), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n559), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n549), .A2(G475), .ZN(new_n646));
  INV_X1    g460(.A(new_n547), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n542), .A2(new_n483), .A3(new_n531), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n525), .A2(new_n526), .B1(new_n529), .B2(new_n528), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n520), .B1(new_n498), .B2(new_n499), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n501), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n648), .B1(new_n651), .B2(new_n483), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n546), .B1(new_n652), .B2(new_n481), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n646), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT33), .B1(new_n461), .B2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(new_n475), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G478), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n414), .A2(new_n396), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n466), .B2(new_n414), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n645), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n642), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT34), .B(G104), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G6));
  INV_X1    g481(.A(KEYINPUT97), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n647), .B2(new_n653), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n545), .A2(KEYINPUT97), .A3(new_n547), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT95), .B1(new_n469), .B2(new_n472), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n477), .A2(new_n474), .A3(new_n478), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n672), .A2(new_n673), .B1(G475), .B2(new_n549), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n559), .A2(new_n671), .A3(new_n644), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n642), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT35), .B(G107), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  NOR2_X1   g492(.A1(new_n623), .A2(KEYINPUT36), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n619), .B(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n633), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n630), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT98), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT98), .B1(new_n630), .B2(new_n682), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n413), .A2(new_n605), .A3(new_n688), .A4(new_n640), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G12));
  OAI21_X1  g505(.A(KEYINPUT32), .B1(new_n330), .B2(new_n332), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n339), .A2(new_n334), .A3(new_n331), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n687), .B1(new_n694), .B2(new_n325), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n646), .B1(new_n473), .B2(new_n479), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n670), .B2(new_n669), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT99), .B(G900), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n554), .B1(new_n556), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n697), .A2(new_n698), .A3(new_n644), .A4(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n671), .A2(new_n644), .A3(new_n674), .A4(new_n701), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n695), .A2(new_n702), .A3(new_n413), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  NAND2_X1  g520(.A1(new_n597), .A2(new_n602), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n707), .B(new_n708), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n672), .A2(new_n673), .ZN(new_n710));
  INV_X1    g524(.A(new_n683), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n643), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n709), .A2(new_n654), .A3(new_n710), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g527(.A(new_n700), .B(KEYINPUT39), .Z(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n411), .A2(new_n412), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n713), .B1(new_n717), .B2(KEYINPUT40), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(KEYINPUT40), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n321), .A2(new_n277), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n396), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n277), .B1(new_n294), .B2(new_n296), .ZN(new_n722));
  OAI21_X1  g536(.A(G472), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n333), .B2(new_n340), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT102), .Z(new_n725));
  NOR2_X1   g539(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n214), .ZN(G45));
  INV_X1    g541(.A(new_n644), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n654), .A2(new_n662), .A3(new_n701), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n341), .A2(new_n413), .A3(new_n730), .A4(new_n688), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G146), .ZN(G48));
  AOI21_X1  g546(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n733));
  AOI211_X1 g547(.A(G469), .B(G902), .C1(new_n386), .C2(new_n393), .ZN(new_n734));
  INV_X1    g548(.A(new_n410), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n341), .A2(new_n664), .A3(new_n634), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT41), .B(G113), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G15));
  NAND4_X1  g553(.A1(new_n675), .A2(new_n341), .A3(new_n634), .A4(new_n736), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G116), .ZN(G18));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n644), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n560), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n695), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(KEYINPUT103), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT103), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n695), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G119), .ZN(G21));
  INV_X1    g563(.A(new_n736), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n480), .B2(new_n550), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n654), .A2(KEYINPUT105), .A3(new_n710), .ZN(new_n753));
  AOI211_X1 g567(.A(new_n750), .B(new_n645), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n297), .A2(new_n308), .ZN(new_n755));
  OAI211_X1 g569(.A(KEYINPUT104), .B(new_n336), .C1(new_n755), .C2(new_n277), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n277), .B1(new_n297), .B2(new_n308), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n757), .B1(new_n758), .B2(new_n328), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n337), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n638), .B1(new_n760), .B2(new_n331), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n754), .A2(new_n634), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR2_X1   g577(.A1(new_n742), .A2(new_n729), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n711), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G125), .ZN(G27));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n341), .A2(new_n634), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n408), .A2(new_n410), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n597), .A2(new_n602), .A3(new_n561), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n729), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n767), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n341), .A2(new_n771), .A3(KEYINPUT42), .A4(new_n634), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NOR2_X1   g590(.A1(new_n769), .A2(new_n770), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n697), .A3(new_n701), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n768), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(new_n188), .ZN(G36));
  AOI21_X1  g594(.A(KEYINPUT45), .B1(new_n403), .B2(new_n405), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n395), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT45), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n407), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n734), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(new_n786), .B2(new_n785), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n788), .A2(new_n410), .A3(new_n714), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT106), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT43), .B1(new_n550), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n550), .A2(new_n662), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n640), .A2(new_n683), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT44), .ZN(new_n797));
  INV_X1    g611(.A(new_n770), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(KEYINPUT44), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT108), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT108), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n790), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(new_n198), .ZN(G39));
  NAND2_X1  g618(.A1(new_n788), .A2(new_n410), .ZN(new_n805));
  XNOR2_X1  g619(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  OR3_X1    g621(.A1(new_n729), .A2(new_n634), .A3(new_n770), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n341), .A3(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(new_n502), .ZN(G42));
  INV_X1    g624(.A(new_n709), .ZN(new_n811));
  INV_X1    g625(.A(new_n562), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n634), .A2(new_n811), .A3(new_n812), .A4(new_n410), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n733), .A2(new_n734), .ZN(new_n814));
  XOR2_X1   g628(.A(new_n814), .B(KEYINPUT110), .Z(new_n815));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n815), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n793), .B1(new_n818), .B2(KEYINPUT49), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n813), .A2(new_n725), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n728), .B1(new_n752), .B2(new_n753), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n769), .A2(new_n711), .A3(new_n700), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n724), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n705), .A2(new_n731), .A3(new_n765), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n731), .A2(new_n823), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(KEYINPUT52), .A3(new_n705), .A4(new_n765), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT53), .B1(new_n829), .B2(KEYINPUT113), .ZN(new_n830));
  INV_X1    g644(.A(new_n747), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n746), .B1(new_n695), .B2(new_n743), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n762), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n635), .A2(new_n737), .A3(new_n689), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT111), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n707), .A2(new_n812), .A3(new_n559), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n835), .B1(new_n836), .B2(new_n663), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n477), .A2(new_n478), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n603), .A2(new_n550), .A3(new_n838), .A4(new_n559), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n550), .A2(new_n661), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n840), .A2(KEYINPUT111), .A3(new_n603), .A4(new_n559), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n837), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n740), .B1(new_n842), .B2(new_n641), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n833), .A2(new_n834), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n838), .A2(new_n700), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n671), .A2(new_n646), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT112), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n798), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n695), .A2(new_n413), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n761), .A2(new_n711), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n849), .A2(new_n850), .B1(new_n851), .B2(new_n771), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n779), .B1(new_n773), .B2(new_n774), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n844), .A2(new_n829), .A3(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n830), .B(new_n855), .Z(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n826), .A2(new_n828), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n843), .A2(new_n834), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n761), .A2(new_n634), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n745), .A2(new_n747), .B1(new_n864), .B2(new_n754), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n865), .A3(new_n853), .A4(new_n852), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n861), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n859), .A2(KEYINPUT53), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n861), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n844), .A2(new_n829), .A3(new_n854), .A4(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT54), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  OR2_X1    g685(.A1(new_n858), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n750), .A2(new_n770), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n725), .A2(new_n634), .A3(new_n554), .A4(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n654), .A3(new_n662), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n864), .A2(new_n554), .A3(new_n794), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n643), .A3(new_n811), .A4(new_n736), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  OR2_X1    g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n815), .A2(new_n735), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT115), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n807), .A2(new_n883), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n876), .A2(new_n798), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n794), .A2(new_n554), .A3(new_n873), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT116), .Z(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n851), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n889), .B2(new_n851), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n881), .B(new_n886), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT51), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n807), .A2(new_n882), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n894), .B1(new_n896), .B2(new_n885), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n881), .B(new_n897), .C1(new_n891), .C2(new_n892), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n876), .A2(new_n644), .A3(new_n736), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n551), .C1(new_n663), .C2(new_n874), .ZN(new_n900));
  INV_X1    g714(.A(new_n768), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n889), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n902), .A2(KEYINPUT48), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(KEYINPUT48), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n895), .A2(new_n898), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n872), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n820), .B1(new_n907), .B2(new_n908), .ZN(G75));
  NOR2_X1   g723(.A1(new_n343), .A2(G952), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n599), .A2(new_n600), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(new_n598), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT55), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n867), .ZN(new_n915));
  INV_X1    g729(.A(new_n870), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(new_n396), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(G210), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n910), .B(new_n920), .C1(new_n918), .C2(new_n922), .ZN(G51));
  XOR2_X1   g737(.A(new_n407), .B(KEYINPUT57), .Z(new_n924));
  NOR3_X1   g738(.A1(new_n915), .A2(new_n916), .A3(new_n857), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n925), .B2(new_n871), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n928), .A2(new_n394), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n917), .A2(new_n783), .A3(new_n782), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n910), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n917), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  INV_X1    g747(.A(new_n652), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n910), .ZN(G60));
  XOR2_X1   g751(.A(new_n657), .B(KEYINPUT120), .Z(new_n938));
  XNOR2_X1  g752(.A(new_n659), .B(KEYINPUT59), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n872), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n910), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n925), .A2(new_n871), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n940), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n945), .ZN(G63));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT121), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT60), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n867), .A2(new_n870), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(KEYINPUT122), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n867), .A2(new_n870), .A3(new_n952), .A4(new_n949), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n631), .A3(new_n953), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n954), .A2(new_n942), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n951), .A2(new_n953), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n680), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(KEYINPUT61), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT124), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  INV_X1    g774(.A(new_n680), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n951), .B2(new_n953), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n942), .B(new_n954), .C1(new_n962), .C2(KEYINPUT123), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n962), .A2(KEYINPUT123), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n959), .B(new_n960), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n957), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n962), .A2(KEYINPUT123), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n955), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n959), .B1(new_n970), .B2(new_n960), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n958), .B1(new_n966), .B2(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n557), .B2(new_n567), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT125), .Z(new_n974));
  INV_X1    g788(.A(new_n844), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n343), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n911), .B1(G898), .B2(new_n343), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n976), .B(new_n977), .Z(G69));
  OAI21_X1  g792(.A(new_n311), .B1(KEYINPUT30), .B2(new_n299), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n510), .A2(new_n515), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n982), .B1(G900), .B2(G953), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n705), .A2(new_n765), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n731), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n901), .A2(new_n821), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n853), .B(new_n987), .C1(new_n790), .C2(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n803), .A2(new_n989), .A3(new_n809), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n984), .B1(new_n990), .B2(new_n343), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT127), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n550), .A2(new_n838), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n770), .B1(new_n994), .B2(new_n663), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n901), .A2(new_n716), .A3(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n803), .A2(new_n809), .A3(new_n997), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n726), .A2(new_n986), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT62), .ZN(new_n1000));
  AOI21_X1  g814(.A(G953), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n981), .B(KEYINPUT126), .Z(new_n1002));
  OAI211_X1 g816(.A(new_n992), .B(new_n993), .C1(new_n1001), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n803), .A2(new_n809), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n1004), .A2(new_n1000), .A3(new_n996), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n1005), .B2(new_n343), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT127), .B1(new_n1006), .B2(new_n991), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n343), .B1(G227), .B2(G900), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n1003), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(G72));
  OR2_X1    g825(.A1(new_n1005), .A2(new_n720), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n990), .A2(new_n278), .A3(new_n318), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n975), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n319), .A2(new_n322), .ZN(new_n1018));
  AOI211_X1 g832(.A(new_n1017), .B(new_n856), .C1(new_n335), .C2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n335), .A2(new_n1017), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n318), .A2(new_n277), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n942), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1014), .A2(new_n1019), .A3(new_n1022), .ZN(G57));
endmodule


