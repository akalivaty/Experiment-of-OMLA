//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1286, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G97), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n212), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n215), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(new_n208), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G33), .A2(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G77), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n249), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  MUX2_X1   g0056(.A(G222), .B(G223), .S(G1698), .Z(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  AND2_X1   g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(new_n208), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n248), .A2(KEYINPUT67), .A3(G1), .A4(G13), .ZN(new_n262));
  AND2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G226), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT66), .A2(G41), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT66), .A2(G41), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n264), .B1(new_n271), .B2(G45), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n261), .A2(G274), .A3(new_n262), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G169), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n208), .B1(new_n212), .B2(new_n253), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT69), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n279), .B(G58), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n253), .A2(G20), .ZN(new_n283));
  OR2_X1    g0083(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n223), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT8), .ZN(new_n287));
  OAI21_X1  g0087(.A(KEYINPUT69), .B1(new_n287), .B2(G58), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n282), .B(new_n283), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g0091(.A(KEYINPUT70), .B(new_n278), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(KEYINPUT71), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT71), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(new_n264), .A3(G13), .A4(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n202), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n277), .B1(new_n295), .B2(new_n297), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n209), .A2(G1), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n300), .B1(new_n304), .B2(new_n202), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n278), .B1(new_n289), .B2(new_n291), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n305), .B1(new_n307), .B2(KEYINPUT70), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n276), .B1(new_n293), .B2(new_n308), .ZN(new_n309));
  OR2_X1    g0109(.A1(new_n309), .A2(KEYINPUT72), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n275), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(KEYINPUT72), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n308), .B2(new_n293), .ZN(new_n317));
  AOI211_X1 g0117(.A(new_n302), .B(new_n277), .C1(new_n295), .C2(new_n297), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G50), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n319), .B(new_n300), .C1(new_n306), .C2(new_n320), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n321), .A2(KEYINPUT74), .A3(new_n292), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT9), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n308), .A2(new_n316), .A3(new_n293), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT74), .B1(new_n321), .B2(new_n292), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n275), .A2(G190), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n329), .B1(new_n330), .B2(new_n275), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n315), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  AOI211_X1 g0133(.A(KEYINPUT10), .B(new_n331), .C1(new_n323), .C2(new_n327), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n314), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n267), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n224), .A2(G1698), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n252), .A2(new_n339), .A3(new_n254), .A4(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT75), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(new_n249), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n261), .A2(G238), .A3(new_n262), .A4(new_n265), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n272), .B2(new_n273), .ZN(new_n347));
  NOR3_X1   g0147(.A1(new_n345), .A2(KEYINPUT13), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT13), .ZN(new_n349));
  INV_X1    g0149(.A(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n341), .A2(new_n342), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n249), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n341), .A2(KEYINPUT75), .A3(new_n342), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n349), .B1(new_n350), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n337), .B(G169), .C1(new_n348), .C2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(G169), .B1(new_n348), .B2(new_n357), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT13), .B1(new_n345), .B2(new_n347), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n350), .A2(new_n356), .A3(new_n349), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n365), .A2(KEYINPUT77), .A3(new_n337), .A4(G169), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n348), .A2(new_n357), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(G179), .ZN(new_n368));
  NAND4_X1  g0168(.A1(new_n360), .A2(new_n362), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n304), .A2(new_n217), .ZN(new_n370));
  XNOR2_X1  g0170(.A(new_n370), .B(KEYINPUT76), .ZN(new_n371));
  INV_X1    g0171(.A(new_n290), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n372), .A2(new_n202), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n209), .A2(G33), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n374), .A2(new_n250), .B1(new_n209), .B2(G68), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n277), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(KEYINPUT11), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(KEYINPUT11), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT12), .B1(new_n298), .B2(G68), .ZN(new_n379));
  OR3_X1    g0179(.A1(new_n298), .A2(KEYINPUT12), .A3(G68), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n377), .A2(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n371), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n369), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n367), .A2(G190), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n365), .A2(G200), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT3), .B(G33), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G232), .A2(G1698), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n338), .A2(G238), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n391), .B(new_n354), .C1(G107), .C2(new_n388), .ZN(new_n392));
  INV_X1    g0192(.A(G244), .ZN(new_n393));
  OAI221_X1 g0193(.A(new_n392), .B1(new_n273), .B2(new_n272), .C1(new_n266), .C2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(G179), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G20), .A2(G77), .ZN(new_n396));
  XNOR2_X1  g0196(.A(KEYINPUT15), .B(G87), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT8), .B(G58), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n396), .B1(new_n397), .B2(new_n374), .C1(new_n372), .C2(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n399), .A2(new_n277), .B1(new_n250), .B2(new_n299), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(new_n250), .B2(new_n304), .ZN(new_n401));
  INV_X1    g0201(.A(G169), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n395), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G190), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n394), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT73), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n401), .B1(G200), .B2(new_n394), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND4_X1   g0209(.A1(new_n383), .A2(new_n387), .A3(new_n404), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT16), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n253), .B2(KEYINPUT3), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n251), .A2(KEYINPUT78), .A3(G33), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n254), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT7), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(G20), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n388), .B2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n217), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n223), .A2(new_n217), .ZN(new_n421));
  OAI21_X1  g0221(.A(G20), .B1(new_n421), .B2(new_n201), .ZN(new_n422));
  INV_X1    g0222(.A(G159), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n423), .B2(new_n372), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n411), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT79), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT79), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n411), .C1(new_n420), .C2(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n255), .A2(new_n417), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n419), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n424), .B1(new_n430), .B2(G68), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n278), .B1(new_n431), .B2(KEYINPUT16), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n426), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n282), .B1(new_n286), .B2(new_n288), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n298), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n318), .B2(new_n434), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n261), .A2(G232), .A3(new_n262), .A4(new_n265), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT80), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n272), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n261), .A2(G274), .A3(new_n262), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n267), .A2(G1698), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G223), .B2(G1698), .ZN(new_n444));
  OAI22_X1  g0244(.A1(new_n444), .A2(new_n255), .B1(new_n253), .B2(new_n219), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n441), .A2(new_n442), .B1(new_n445), .B2(new_n354), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G169), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(G179), .A3(new_n446), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n437), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(KEYINPUT18), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n433), .A2(new_n436), .B1(new_n448), .B2(new_n449), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT18), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n440), .A2(new_n405), .A3(new_n446), .ZN(new_n456));
  NOR2_X1   g0256(.A1(G223), .A2(G1698), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n457), .B1(new_n267), .B2(G1698), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n388), .B1(G33), .B2(G87), .ZN(new_n459));
  OAI22_X1  g0259(.A1(new_n459), .A2(new_n249), .B1(new_n272), .B2(new_n273), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n438), .A2(new_n439), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n438), .A2(new_n439), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n456), .B1(new_n463), .B2(G200), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(new_n433), .A3(new_n436), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT17), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n464), .A2(new_n433), .A3(KEYINPUT17), .A4(new_n436), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n452), .A2(new_n455), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AND3_X1   g0270(.A1(new_n336), .A2(new_n410), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n298), .A2(G97), .ZN(new_n473));
  XNOR2_X1  g0273(.A(G97), .B(G107), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT6), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NOR3_X1   g0276(.A1(new_n475), .A2(new_n225), .A3(G107), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n479), .A2(G20), .B1(G77), .B2(new_n290), .ZN(new_n480));
  INV_X1    g0280(.A(G107), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n255), .A2(new_n209), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n473), .B1(new_n484), .B2(new_n277), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n393), .A2(G1698), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n388), .A2(KEYINPUT4), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT4), .B1(new_n388), .B2(new_n486), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n388), .A2(G250), .A3(G1698), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n249), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT5), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n264), .B(G45), .C1(new_n495), .C2(G41), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n496), .B1(new_n271), .B2(new_n495), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n442), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT5), .B1(new_n269), .B2(new_n270), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n261), .B(new_n262), .C1(new_n499), .C2(new_n496), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n226), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(G200), .B1(new_n494), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n264), .A2(G33), .ZN(new_n503));
  XNOR2_X1  g0303(.A(new_n503), .B(KEYINPUT81), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n301), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT82), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT82), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n301), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(G97), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n388), .A2(new_n486), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n512), .A2(new_n492), .A3(new_n491), .A4(new_n487), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n354), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n261), .A2(new_n262), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n497), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G257), .B1(new_n497), .B2(new_n442), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n517), .A3(G190), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n485), .A2(new_n502), .A3(new_n509), .A4(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n393), .A2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n388), .B(new_n520), .C1(G238), .C2(G1698), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n521), .B1(new_n253), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n354), .ZN(new_n524));
  INV_X1    g0324(.A(G45), .ZN(new_n525));
  OR3_X1    g0325(.A1(new_n525), .A2(G1), .A3(G274), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n220), .B1(new_n525), .B2(G1), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n261), .A2(new_n526), .A3(new_n262), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n402), .ZN(new_n530));
  AND2_X1   g0330(.A1(new_n526), .A2(new_n527), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n523), .A2(new_n354), .B1(new_n263), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n311), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n388), .A2(new_n209), .A3(G68), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT19), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n535), .B1(new_n374), .B2(new_n225), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n209), .B1(new_n342), .B2(new_n535), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n219), .A2(new_n225), .A3(new_n481), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT83), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(KEYINPUT83), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n537), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(new_n397), .ZN(new_n545));
  OAI22_X1  g0345(.A1(new_n544), .A2(new_n278), .B1(new_n298), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n301), .A2(new_n507), .A3(new_n504), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n507), .B1(new_n301), .B2(new_n504), .ZN(new_n548));
  NOR3_X1   g0348(.A1(new_n547), .A2(new_n548), .A3(new_n397), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n530), .B(new_n533), .C1(new_n546), .C2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n477), .B1(new_n475), .B2(new_n474), .ZN(new_n551));
  OAI22_X1  g0351(.A1(new_n551), .A2(new_n209), .B1(new_n250), .B2(new_n372), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n481), .B1(new_n418), .B2(new_n419), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n277), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n473), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n509), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n402), .B1(new_n494), .B2(new_n501), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n514), .A2(new_n517), .A3(new_n311), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n529), .A2(G200), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n547), .A2(new_n548), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n543), .A2(new_n541), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n534), .A3(new_n536), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n277), .B1(new_n299), .B2(new_n397), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n532), .A2(G190), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n560), .A2(new_n562), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n519), .A2(new_n550), .A3(new_n559), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n295), .A2(new_n522), .A3(new_n297), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT85), .ZN(new_n570));
  XNOR2_X1  g0370(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n301), .A2(new_n504), .A3(G116), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n492), .B(new_n209), .C1(G33), .C2(new_n225), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n522), .A2(G20), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n573), .A2(new_n277), .A3(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n571), .A2(new_n572), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n388), .A2(G264), .A3(G1698), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n388), .A2(G257), .A3(new_n338), .ZN(new_n581));
  XNOR2_X1  g0381(.A(KEYINPUT84), .B(G303), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n255), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n354), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n263), .B(G270), .C1(new_n499), .C2(new_n496), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(new_n498), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n579), .B(new_n588), .C1(new_n405), .C2(new_n587), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n578), .A2(G169), .A3(new_n587), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(G179), .A2(new_n585), .A3(new_n586), .A4(new_n498), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n578), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n578), .A2(KEYINPUT21), .A3(new_n587), .A4(G169), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n589), .A2(new_n592), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n568), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n220), .A2(G1698), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(new_n252), .A3(new_n254), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT86), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n388), .A2(G257), .A3(G1698), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT86), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n388), .A2(new_n603), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G294), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n354), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n516), .A2(G264), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n607), .A2(new_n608), .A3(new_n498), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(new_n311), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n606), .A2(new_n354), .B1(new_n516), .B2(G264), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n402), .B1(new_n611), .B2(new_n498), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n598), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n609), .A2(G169), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n614), .B(KEYINPUT87), .C1(new_n311), .C2(new_n609), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n298), .A2(G107), .ZN(new_n616));
  OR2_X1    g0416(.A1(new_n616), .A2(KEYINPUT25), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(KEYINPUT25), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n561), .A2(G107), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n252), .A2(new_n254), .A3(new_n209), .A4(G87), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT22), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT22), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n388), .A2(new_n622), .A3(new_n209), .A4(G87), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT24), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT23), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n209), .B2(G107), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n481), .A2(KEYINPUT23), .A3(G20), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n627), .A2(new_n628), .B1(new_n283), .B2(G116), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n625), .B1(new_n624), .B2(new_n629), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n277), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n619), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n613), .A2(new_n615), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT88), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT88), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n613), .A2(new_n615), .A3(new_n636), .A4(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n609), .A2(G200), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n611), .A2(G190), .A3(new_n498), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n619), .A2(new_n638), .A3(new_n639), .A4(new_n632), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n597), .A2(new_n635), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n472), .A2(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n467), .A2(new_n468), .ZN(new_n643));
  INV_X1    g0443(.A(new_n404), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n387), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n643), .B1(new_n383), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n453), .B(KEYINPUT18), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI22_X1  g0448(.A1(new_n646), .A2(new_n648), .B1(new_n333), .B2(new_n334), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n314), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT91), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n640), .A2(new_n519), .A3(new_n559), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n633), .B1(new_n612), .B2(new_n610), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n594), .A2(new_n595), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(new_n656), .A3(new_n592), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n547), .A2(new_n548), .A3(new_n219), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT90), .B1(new_n546), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT90), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n562), .A2(new_n565), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n528), .B(KEYINPUT89), .Z(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n524), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n664), .A2(G200), .B1(G190), .B2(new_n532), .ZN(new_n665));
  INV_X1    g0465(.A(new_n549), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n666), .A2(new_n565), .B1(new_n311), .B2(new_n532), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n664), .A2(new_n402), .ZN(new_n668));
  AOI22_X1  g0468(.A1(new_n662), .A2(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n654), .A2(new_n657), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n667), .A2(new_n668), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n662), .A2(new_n665), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n671), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND4_X1   g0477(.A1(KEYINPUT26), .A2(new_n674), .A3(new_n550), .A4(new_n567), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n672), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n471), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n652), .A2(new_n682), .ZN(G369));
  NAND3_X1  g0483(.A1(new_n264), .A2(new_n209), .A3(G13), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(KEYINPUT27), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G213), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(G343), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n579), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n596), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n656), .A2(new_n592), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n691), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(KEYINPUT92), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(G330), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n633), .A2(new_n689), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n635), .A2(new_n637), .A3(new_n640), .A4(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n634), .A2(new_n690), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT93), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n705), .A2(KEYINPUT93), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n693), .A2(new_n690), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n707), .B2(new_n708), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n655), .A2(new_n689), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n710), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n271), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n213), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n539), .A2(G116), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(G1), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n206), .B2(new_n719), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n689), .B1(new_n672), .B2(new_n680), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n635), .A2(new_n637), .A3(new_n592), .A4(new_n656), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n726), .A2(new_n669), .A3(new_n654), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n674), .A2(new_n550), .A3(new_n567), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n671), .B1(new_n728), .B2(KEYINPUT26), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(KEYINPUT26), .B2(new_n675), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n689), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT94), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n611), .A2(new_n532), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n494), .A2(new_n501), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT30), .A4(new_n593), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT30), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n611), .A2(new_n532), .A3(new_n514), .A4(new_n517), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n585), .A2(new_n586), .A3(G179), .A4(new_n498), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(G179), .B1(new_n514), .B2(new_n517), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n742), .A2(new_n664), .A3(new_n609), .A4(new_n587), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n737), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n745));
  AOI21_X1  g0545(.A(KEYINPUT31), .B1(new_n744), .B2(new_n689), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n734), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n744), .A2(new_n689), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(KEYINPUT31), .A3(new_n689), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(KEYINPUT94), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n641), .A2(new_n689), .ZN(new_n754));
  OAI21_X1  g0554(.A(G330), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n733), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT95), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n733), .A2(KEYINPUT95), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n723), .B1(new_n760), .B2(G1), .ZN(G364));
  NAND2_X1  g0561(.A1(new_n698), .A2(new_n699), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT96), .ZN(new_n763));
  INV_X1    g0563(.A(G13), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n264), .B1(new_n765), .B2(G45), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n719), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n763), .A2(new_n701), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n767), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n388), .A2(new_n213), .ZN(new_n770));
  INV_X1    g0570(.A(G355), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n770), .A2(new_n771), .B1(G116), .B2(new_n213), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n242), .A2(new_n525), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n255), .A2(new_n213), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n207), .B2(new_n525), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G13), .A2(G33), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G20), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n208), .B1(G20), .B2(new_n402), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n769), .B1(new_n776), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n209), .A2(new_n405), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n311), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(KEYINPUT97), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n786), .A2(KEYINPUT97), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G322), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n330), .A2(G179), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n209), .A2(G190), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(G283), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n255), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n405), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(G326), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G179), .A2(G200), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n209), .B1(new_n801), .B2(G190), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n798), .A2(G190), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(G294), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n784), .A2(new_n793), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n794), .A2(new_n785), .ZN(new_n809));
  INV_X1    g0609(.A(G311), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n807), .A2(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n794), .A2(new_n801), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n811), .B1(G329), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g0614(.A1(new_n792), .A2(new_n800), .A3(new_n806), .A4(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n790), .A2(new_n223), .B1(new_n250), .B2(new_n809), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT98), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n388), .B1(new_n807), .B2(new_n219), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n812), .A2(new_n423), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT32), .ZN(new_n821));
  INV_X1    g0621(.A(new_n799), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n820), .A2(new_n821), .B1(new_n202), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n795), .ZN(new_n824));
  AOI211_X1 g0624(.A(new_n819), .B(new_n823), .C1(G107), .C2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n802), .A2(new_n225), .ZN(new_n826));
  INV_X1    g0626(.A(new_n804), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n217), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(new_n821), .C2(new_n820), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n818), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n816), .A2(new_n817), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n815), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n783), .B1(new_n832), .B2(new_n780), .ZN(new_n833));
  INV_X1    g0633(.A(new_n779), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n695), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n768), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  NOR2_X1   g0637(.A1(new_n404), .A2(new_n689), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n407), .A2(new_n408), .B1(new_n401), .B2(new_n689), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n840), .B2(new_n644), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n724), .B(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(new_n755), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT100), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n769), .B1(new_n843), .B2(new_n755), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n809), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G159), .B1(G137), .B2(new_n799), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n827), .C1(new_n790), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT34), .Z(new_n853));
  NOR2_X1   g0653(.A1(new_n802), .A2(new_n223), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n388), .B1(new_n807), .B2(new_n202), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n795), .A2(new_n217), .B1(new_n812), .B2(new_n856), .ZN(new_n857));
  NOR4_X1   g0657(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n857), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n255), .B1(new_n809), .B2(new_n522), .C1(new_n481), .C2(new_n807), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n791), .B2(G294), .ZN(new_n860));
  OAI22_X1  g0660(.A1(new_n795), .A2(new_n219), .B1(new_n812), .B2(new_n810), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT99), .Z(new_n862));
  NOR2_X1   g0662(.A1(new_n822), .A2(new_n808), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n826), .B(new_n863), .C1(G283), .C2(new_n804), .ZN(new_n864));
  AND3_X1   g0664(.A1(new_n860), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n780), .B1(new_n858), .B2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n780), .A2(new_n777), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n767), .B1(new_n250), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n401), .A2(new_n689), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n409), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n838), .B1(new_n870), .B2(new_n404), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n866), .B(new_n868), .C1(new_n871), .C2(new_n778), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n847), .A2(new_n872), .ZN(G384));
  NOR2_X1   g0673(.A1(new_n765), .A2(new_n264), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n670), .A2(new_n671), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n678), .B1(new_n675), .B2(new_n676), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n871), .B(new_n690), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n839), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n382), .A2(new_n689), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n383), .A2(new_n387), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n387), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n382), .B(new_n689), .C1(new_n881), .C2(new_n369), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n431), .A2(KEYINPUT16), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n277), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n431), .A2(KEYINPUT16), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n436), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n687), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g0691(.A1(new_n467), .A2(new_n468), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n891), .B1(new_n647), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT37), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n889), .B1(new_n450), .B2(new_n890), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n895), .B2(new_n465), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n437), .A2(new_n890), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT101), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT101), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n437), .A2(new_n899), .A3(new_n890), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g0701(.A(KEYINPUT102), .B(KEYINPUT37), .Z(new_n902));
  AND3_X1   g0702(.A1(new_n451), .A2(new_n465), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n896), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n885), .B1(new_n893), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n891), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n469), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n895), .A2(new_n465), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n899), .B1(new_n437), .B2(new_n890), .ZN(new_n910));
  AOI211_X1 g0710(.A(KEYINPUT101), .B(new_n687), .C1(new_n433), .C2(new_n436), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n451), .A2(new_n465), .A3(new_n902), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n909), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n914), .A3(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n905), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n884), .A2(new_n917), .B1(new_n647), .B2(new_n890), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n383), .A2(new_n689), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT103), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n907), .A2(KEYINPUT38), .A3(new_n914), .ZN(new_n922));
  AOI21_X1  g0722(.A(KEYINPUT38), .B1(new_n907), .B2(new_n914), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n921), .B(KEYINPUT39), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n451), .A2(new_n465), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n902), .B1(new_n901), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n469), .A2(new_n912), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n901), .A2(new_n903), .ZN(new_n930));
  XNOR2_X1  g0730(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n915), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n924), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n921), .B1(new_n916), .B2(KEYINPUT39), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n920), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n725), .A2(new_n471), .A3(new_n732), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n652), .A2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n745), .A2(new_n746), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n943), .B1(new_n641), .B2(new_n689), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n841), .B1(new_n880), .B2(new_n882), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n931), .B1(new_n912), .B2(new_n913), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n927), .B2(new_n928), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n944), .B(new_n945), .C1(new_n922), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT40), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT40), .B1(new_n905), .B2(new_n915), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n944), .A2(new_n883), .A3(new_n871), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n471), .A3(new_n944), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n948), .A2(KEYINPUT40), .B1(new_n950), .B2(new_n951), .ZN(new_n955));
  INV_X1    g0755(.A(new_n944), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n472), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n954), .A2(G330), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n874), .B1(new_n942), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n942), .B2(new_n958), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n479), .A2(KEYINPUT35), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n961), .A2(G116), .A3(new_n210), .A4(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT36), .ZN(new_n964));
  NOR3_X1   g0764(.A1(new_n421), .A2(new_n206), .A3(new_n250), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n217), .A2(G50), .ZN(new_n966));
  OAI211_X1 g0766(.A(G1), .B(new_n764), .C1(new_n965), .C2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n960), .A2(new_n964), .A3(new_n967), .ZN(G367));
  OAI221_X1 g0768(.A(new_n781), .B1(new_n213), .B2(new_n397), .C1(new_n238), .C2(new_n774), .ZN(new_n969));
  AND2_X1   g0769(.A1(new_n969), .A2(new_n769), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n659), .A2(new_n661), .A3(new_n689), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n669), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n671), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n582), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n790), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n388), .B1(new_n848), .B2(G283), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n824), .A2(G97), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n978), .C1(new_n979), .C2(new_n812), .ZN(new_n980));
  INV_X1    g0780(.A(new_n807), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n807), .B2(new_n522), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(new_n822), .C2(new_n810), .ZN(new_n985));
  INV_X1    g0785(.A(G294), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n827), .A2(new_n986), .B1(new_n802), .B2(new_n481), .ZN(new_n987));
  NOR4_X1   g0787(.A1(new_n976), .A2(new_n980), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n803), .A2(G68), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n851), .B2(new_n822), .C1(new_n790), .C2(new_n850), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT109), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n807), .A2(new_n223), .B1(new_n795), .B2(new_n250), .ZN(new_n992));
  INV_X1    g0792(.A(G137), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n388), .B1(new_n812), .B2(new_n993), .C1(new_n827), .C2(new_n423), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n992), .B(new_n994), .C1(G50), .C2(new_n848), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n988), .B1(new_n991), .B2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT47), .ZN(new_n997));
  INV_X1    g0797(.A(new_n780), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n970), .B1(new_n974), .B2(new_n834), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n766), .B(KEYINPUT108), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n556), .A2(new_n689), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n519), .A2(new_n559), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n674), .A2(new_n689), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT107), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT44), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n716), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n716), .B(new_n1008), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n713), .A2(new_n715), .A3(new_n1005), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT45), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n710), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1014), .B(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n710), .ZN(new_n1019));
  NAND4_X1  g0819(.A1(new_n1018), .A2(new_n1019), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n708), .A2(new_n707), .A3(new_n712), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n700), .A3(new_n713), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n708), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n711), .B1(new_n1024), .B2(new_n706), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n701), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n758), .B2(new_n759), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1016), .A2(new_n1020), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n760), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n719), .B(KEYINPUT41), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1001), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n712), .B(new_n1005), .C1(new_n707), .C2(new_n708), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT42), .ZN(new_n1035));
  AND2_X1   g0835(.A1(new_n635), .A2(new_n637), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n559), .B1(new_n1036), .B2(new_n1003), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n690), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(KEYINPUT105), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT106), .ZN(new_n1040));
  OR3_X1    g0840(.A1(new_n1034), .A2(new_n1040), .A3(KEYINPUT42), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1040), .B1(new_n1034), .B2(KEYINPUT42), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT43), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n974), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT105), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g0849(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1046), .A2(new_n1045), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1049), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1051), .B(new_n1052), .C1(new_n1053), .C2(new_n1043), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n710), .A2(new_n1005), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1050), .A2(new_n1054), .A3(new_n710), .A4(new_n1005), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n999), .B1(new_n1033), .B2(new_n1059), .ZN(G387));
  NOR2_X1   g0860(.A1(new_n1028), .A2(new_n719), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1027), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1061), .B1(new_n760), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n770), .A2(new_n720), .B1(G107), .B2(new_n213), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n235), .A2(new_n525), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n720), .ZN(new_n1066));
  AOI211_X1 g0866(.A(G45), .B(new_n1066), .C1(G68), .C2(G77), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n398), .A2(G50), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT50), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n774), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1064), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n848), .A2(new_n582), .B1(G311), .B2(new_n804), .ZN(new_n1072));
  INV_X1    g0872(.A(G322), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n822), .C1(new_n790), .C2(new_n979), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n981), .A2(G294), .B1(new_n803), .B2(G283), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n388), .B1(new_n813), .B2(G326), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n522), .B2(new_n795), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n434), .A2(new_n827), .B1(new_n217), .B2(new_n809), .ZN(new_n1086));
  XNOR2_X1  g0886(.A(new_n1086), .B(KEYINPUT110), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n803), .A2(new_n545), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n822), .B2(new_n423), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n981), .A2(G77), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n813), .A2(G150), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1090), .A2(new_n978), .A3(new_n1091), .A4(new_n388), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1089), .B(new_n1092), .C1(new_n791), .C2(G50), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1084), .A2(new_n1085), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n769), .B1(new_n782), .B2(new_n1071), .C1(new_n1094), .C2(new_n998), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n709), .B2(new_n779), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n1062), .B2(new_n1001), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1063), .A2(new_n1097), .ZN(G393));
  INV_X1    g0898(.A(new_n1016), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1020), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1003), .A2(new_n1004), .A3(new_n779), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n781), .B1(new_n225), .B2(new_n213), .C1(new_n245), .C2(new_n774), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n769), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT111), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n255), .B1(new_n795), .B2(new_n481), .C1(new_n975), .C2(new_n827), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G283), .A2(new_n981), .B1(new_n848), .B2(G294), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n1073), .B2(new_n812), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(G116), .C2(new_n803), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n791), .A2(G311), .B1(G317), .B2(new_n799), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT52), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1109), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n790), .A2(new_n423), .B1(new_n850), .B2(new_n822), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT51), .Z(new_n1117));
  AOI22_X1  g0917(.A1(G68), .A2(new_n981), .B1(new_n813), .B2(G143), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n388), .C1(new_n219), .C2(new_n795), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT112), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n802), .A2(new_n250), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n398), .B2(new_n809), .C1(new_n827), .C2(new_n202), .ZN(new_n1123));
  OR3_X1    g0923(.A1(new_n1117), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1114), .A2(KEYINPUT113), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1115), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1105), .B1(new_n1126), .B2(new_n780), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1101), .A2(new_n1001), .B1(new_n1102), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1028), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n719), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1029), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1128), .A2(new_n1132), .ZN(G390));
  AOI21_X1  g0933(.A(new_n767), .B1(new_n434), .B2(new_n867), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT115), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n791), .A2(G132), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n807), .A2(new_n850), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT53), .ZN(new_n1138));
  INV_X1    g0938(.A(G128), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1137), .A2(new_n1138), .B1(new_n1139), .B2(new_n822), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n1138), .B2(new_n1137), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT54), .B(G143), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n809), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n388), .B1(new_n795), .B2(new_n202), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(G125), .C2(new_n813), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n803), .A2(G159), .B1(G137), .B2(new_n804), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1136), .A2(new_n1141), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n791), .A2(G116), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n388), .B(new_n1121), .C1(G87), .C2(new_n981), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G107), .A2(new_n804), .B1(new_n799), .B2(G283), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n217), .A2(new_n795), .B1(new_n809), .B2(new_n225), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(G294), .B2(new_n813), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1147), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT39), .B1(new_n922), .B2(new_n923), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(KEYINPUT103), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n935), .A3(new_n924), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1135), .B1(new_n998), .B2(new_n1154), .C1(new_n1157), .C2(new_n778), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n944), .A2(G330), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n945), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n920), .B1(new_n878), .B2(new_n883), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n936), .A2(new_n937), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(new_n920), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n933), .A2(new_n915), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n870), .A2(new_n404), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n838), .B1(new_n731), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n883), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1164), .B(new_n1165), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1161), .B1(new_n1163), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n884), .A2(new_n1164), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1172), .A2(new_n1156), .A3(new_n935), .A4(new_n924), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G330), .B(new_n871), .C1(new_n753), .C2(new_n754), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1174), .A2(new_n1168), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1158), .B1(new_n1177), .B2(new_n1000), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1159), .A2(new_n871), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1168), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1180), .A2(new_n1175), .A3(new_n1167), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1174), .A2(new_n1168), .B1(new_n1159), .B2(new_n945), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n878), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT114), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1174), .A2(new_n1168), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1160), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT114), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(new_n1188), .A3(new_n878), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1185), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1182), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n471), .A2(new_n1159), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n652), .A2(new_n940), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n719), .B1(new_n1195), .B2(new_n1177), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1173), .A2(new_n1169), .A3(new_n1175), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1160), .B1(new_n1173), .B2(new_n1169), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1194), .A3(new_n1191), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1178), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G378));
  INV_X1    g1002(.A(KEYINPUT57), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1193), .B1(new_n1199), .B2(new_n1191), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n890), .B1(new_n317), .B2(new_n322), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT55), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n335), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1206), .B(new_n314), .C1(new_n333), .C2(new_n334), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1209), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n953), .B2(G330), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n955), .A2(new_n699), .A3(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n939), .B1(new_n1214), .B2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n918), .B1(new_n1157), .B2(new_n920), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n953), .A2(G330), .A3(new_n1213), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(new_n955), .B2(new_n699), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1217), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1203), .B1(new_n1204), .B2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1181), .B1(new_n1189), .B2(new_n1185), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1194), .B1(new_n1177), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT118), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT118), .B1(new_n1228), .B2(new_n939), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1225), .B(KEYINPUT57), .C1(new_n1227), .C2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1223), .A2(new_n1230), .A3(new_n1131), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1222), .A2(new_n1000), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1215), .A2(new_n777), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n271), .A2(new_n388), .ZN(new_n1234));
  INV_X1    g1034(.A(G41), .ZN(new_n1235));
  AOI211_X1 g1035(.A(G50), .B(new_n1234), .C1(new_n253), .C2(new_n1235), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(G58), .A2(new_n824), .B1(new_n813), .B2(G283), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(new_n397), .B2(new_n809), .C1(new_n790), .C2(new_n481), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1090), .A2(new_n989), .A3(new_n1234), .ZN(new_n1239));
  OAI22_X1  g1039(.A1(new_n827), .A2(new_n225), .B1(new_n822), .B2(new_n522), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1238), .A2(new_n1239), .A3(new_n1240), .ZN(new_n1241));
  XOR2_X1   g1041(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n1242));
  AOI21_X1  g1042(.A(new_n1236), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n807), .A2(new_n1142), .B1(new_n809), .B2(new_n993), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G132), .B2(new_n804), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n803), .A2(G150), .B1(G125), .B2(new_n799), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1245), .B(new_n1246), .C1(new_n1139), .C2(new_n790), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(KEYINPUT59), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n253), .B(new_n1235), .C1(new_n795), .C2(new_n423), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G124), .B2(new_n813), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n1243), .B1(new_n1248), .B2(new_n1252), .C1(new_n1242), .C2(new_n1241), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1253), .A2(new_n780), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n767), .B(new_n1254), .C1(new_n202), .C2(new_n867), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1232), .B1(new_n1233), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1231), .A2(new_n1256), .ZN(G375));
  NAND2_X1  g1057(.A1(new_n1168), .A2(new_n777), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n809), .A2(new_n850), .B1(new_n812), .B2(new_n1139), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n388), .B1(new_n802), .B2(new_n202), .C1(new_n223), .C2(new_n795), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1259), .B(new_n1260), .C1(G159), .C2(new_n981), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT120), .Z(new_n1262));
  OAI22_X1  g1062(.A1(new_n856), .A2(new_n822), .B1(new_n827), .B2(new_n1142), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(new_n791), .B2(G137), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n807), .A2(new_n225), .B1(new_n812), .B2(new_n808), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1266), .B(KEYINPUT119), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n790), .A2(new_n796), .ZN(new_n1268));
  OAI221_X1 g1068(.A(new_n1088), .B1(new_n822), .B2(new_n986), .C1(new_n522), .C2(new_n827), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n255), .B1(new_n795), .B2(new_n250), .C1(new_n481), .C2(new_n809), .ZN(new_n1270));
  OR4_X1    g1070(.A1(new_n1267), .A2(new_n1268), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n998), .B1(new_n1265), .B2(new_n1271), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n767), .B(new_n1272), .C1(new_n217), .C2(new_n867), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1191), .A2(new_n1001), .B1(new_n1258), .B2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1195), .A2(new_n1032), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1224), .A2(new_n1193), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1275), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(G381));
  AND2_X1   g1080(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .A4(new_n1279), .ZN(new_n1284));
  OR4_X1    g1084(.A1(G387), .A2(new_n1284), .A3(G375), .A4(G378), .ZN(G407));
  NAND2_X1  g1085(.A1(new_n688), .A2(G213), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1286), .B(KEYINPUT121), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1201), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G375), .C2(new_n1288), .ZN(G409));
  OAI21_X1  g1089(.A(new_n1001), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1233), .A2(new_n1255), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1031), .B1(new_n1217), .B2(new_n1221), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1225), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1201), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT122), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1231), .A2(new_n1256), .A3(G378), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1294), .A2(KEYINPUT122), .A3(new_n1201), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1297), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1287), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1224), .A2(KEYINPUT60), .A3(new_n1193), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(new_n1131), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1195), .A2(KEYINPUT60), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1278), .B2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1283), .B1(new_n1305), .B2(new_n1275), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1304), .A2(new_n1278), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G384), .B(new_n1274), .C1(new_n1307), .C2(new_n1303), .ZN(new_n1308));
  AND2_X1   g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1300), .A2(new_n1301), .A3(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  NOR2_X1   g1111(.A1(new_n1311), .A2(KEYINPUT125), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1287), .A2(G2897), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1306), .A2(new_n1308), .A3(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1315), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1314), .A2(new_n1318), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1300), .A2(new_n1301), .A3(new_n1309), .A4(new_n1320), .ZN(new_n1321));
  XNOR2_X1  g1121(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1313), .A2(new_n1319), .A3(new_n1321), .A4(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT123), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(G387), .B2(new_n1281), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n836), .B1(new_n1063), .B2(new_n1097), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1282), .A2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1031), .B1(new_n1029), .B2(new_n760), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1058), .B(new_n1057), .C1(new_n1328), .C2(new_n1001), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(G390), .A2(new_n1329), .A3(new_n999), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(G390), .B1(new_n1329), .B2(new_n999), .ZN(new_n1332));
  OAI22_X1  g1132(.A1(new_n1325), .A2(new_n1327), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1327), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(new_n1281), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1334), .A2(new_n1335), .A3(new_n1324), .A4(new_n1330), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1333), .A2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1323), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1310), .A2(KEYINPUT63), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1300), .A2(new_n1341), .A3(new_n1301), .A4(new_n1309), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT61), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1319), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1339), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(KEYINPUT126), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT126), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1339), .A2(new_n1348), .A3(new_n1345), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1349), .ZN(G405));
  XNOR2_X1  g1150(.A(G375), .B(G378), .ZN(new_n1351));
  XNOR2_X1  g1151(.A(new_n1351), .B(new_n1309), .ZN(new_n1352));
  AND3_X1   g1152(.A1(new_n1352), .A2(new_n1338), .A3(KEYINPUT127), .ZN(new_n1353));
  AOI21_X1  g1153(.A(KEYINPUT127), .B1(new_n1352), .B2(new_n1338), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1352), .A2(new_n1338), .ZN(new_n1355));
  NOR3_X1   g1155(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .ZN(G402));
endmodule


