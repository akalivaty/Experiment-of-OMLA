//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084, new_n1085;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT73), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  OR2_X1    g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n191), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G110), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT70), .B1(new_n195), .B2(G119), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT70), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n199), .A3(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(new_n196), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n203), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT71), .A2(G125), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(KEYINPUT71), .A2(G125), .ZN(new_n214));
  OAI21_X1  g028(.A(G140), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(G125), .A2(G140), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n211), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT71), .A2(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n212), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT16), .A2(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n210), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G140), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n219), .B2(new_n212), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT16), .B1(new_n226), .B2(new_n216), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(G146), .A3(new_n222), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n209), .B1(new_n224), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n204), .ZN(new_n230));
  INV_X1    g044(.A(G110), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n198), .A2(new_n201), .A3(new_n231), .A4(new_n200), .ZN(new_n232));
  AND2_X1   g046(.A1(G125), .A2(G140), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n210), .B1(new_n233), .B2(new_n216), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G125), .B(G140), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(KEYINPUT72), .A3(new_n210), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n230), .A2(new_n232), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n228), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n194), .B1(new_n229), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n208), .A2(new_n204), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(G110), .B2(new_n202), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n218), .A2(new_n223), .A3(new_n210), .ZN(new_n245));
  AOI21_X1  g059(.A(G146), .B1(new_n227), .B2(new_n222), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n244), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n194), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n240), .ZN(new_n249));
  INV_X1    g063(.A(G902), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n242), .A2(new_n249), .A3(KEYINPUT25), .A4(new_n250), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(KEYINPUT74), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G217), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n256), .B1(G234), .B2(new_n250), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT74), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(new_n258), .A3(new_n252), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n242), .A2(new_n249), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n257), .A2(G902), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n260), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT27), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT69), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n210), .A2(G143), .ZN(new_n273));
  INV_X1    g087(.A(G143), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  OR2_X1    g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G143), .B(G146), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT0), .A3(G128), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT11), .ZN(new_n283));
  INV_X1    g097(.A(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(G137), .ZN(new_n285));
  INV_X1    g099(.A(G137), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(KEYINPUT11), .A3(G134), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(G137), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G131), .ZN(new_n290));
  AOI21_X1  g104(.A(G131), .B1(new_n284), .B2(G137), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n285), .A2(new_n291), .A3(new_n287), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n284), .A2(G137), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n286), .A2(G134), .ZN(new_n295));
  OAI21_X1  g109(.A(G131), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(new_n292), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT1), .B1(new_n274), .B2(G146), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n276), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n280), .A2(new_n302), .A3(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n282), .A2(new_n293), .B1(new_n298), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n199), .A2(G116), .ZN(new_n306));
  INV_X1    g120(.A(G116), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G119), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G113), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT2), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G113), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n313), .ZN(new_n315));
  XNOR2_X1  g129(.A(G116), .B(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n317), .A3(KEYINPUT66), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n317), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT66), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n305), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT28), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n272), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n285), .A2(new_n291), .A3(new_n287), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n286), .A2(G134), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(new_n288), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT64), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT64), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n296), .A2(new_n292), .A3(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n329), .A2(KEYINPUT65), .A3(new_n331), .A4(new_n304), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n282), .A2(new_n293), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n297), .A2(KEYINPUT64), .B1(new_n301), .B2(new_n303), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT65), .B1(new_n335), .B2(new_n331), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n319), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(new_n322), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n324), .B1(new_n338), .B2(KEYINPUT28), .ZN(new_n339));
  AOI211_X1 g153(.A(new_n272), .B(new_n323), .C1(new_n337), .C2(new_n322), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n271), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AND4_X1   g155(.A1(new_n302), .A2(new_n273), .A3(new_n275), .A4(G128), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n299), .A2(G128), .B1(new_n273), .B2(new_n275), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n292), .B(new_n296), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n333), .A2(KEYINPUT30), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n319), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n329), .A2(new_n331), .A3(new_n304), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT65), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n333), .A3(new_n332), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT30), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n325), .B1(G131), .B2(new_n289), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n279), .A2(new_n281), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n344), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n321), .A2(new_n318), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n270), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n352), .A2(KEYINPUT31), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n341), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT67), .B1(new_n352), .B2(new_n357), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n351), .B1(new_n334), .B2(new_n336), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n305), .A2(KEYINPUT30), .B1(new_n314), .B2(new_n317), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT67), .ZN(new_n365));
  INV_X1    g179(.A(new_n357), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(KEYINPUT31), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT68), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n361), .A2(new_n370), .A3(new_n367), .A4(KEYINPUT31), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n360), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(G472), .A2(G902), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n265), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G472), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n338), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n323), .B1(new_n337), .B2(new_n322), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n377), .B(new_n270), .C1(new_n378), .C2(new_n324), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n364), .A2(new_n322), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n380), .B2(new_n271), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n355), .A2(new_n356), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n323), .B1(new_n322), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n384), .B1(new_n323), .B2(new_n322), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n270), .A2(KEYINPUT29), .ZN(new_n386));
  AOI21_X1  g200(.A(G902), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n376), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n377), .B1(new_n378), .B2(new_n324), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n358), .B1(new_n389), .B2(new_n271), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n365), .B1(new_n364), .B2(new_n366), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT67), .B(new_n357), .C1(new_n362), .C2(new_n363), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n370), .B1(new_n393), .B2(KEYINPUT31), .ZN(new_n394));
  INV_X1    g208(.A(new_n371), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n374), .A2(new_n265), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n388), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n264), .B1(new_n375), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G478), .B1(KEYINPUT85), .B2(KEYINPUT15), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n400), .B1(KEYINPUT85), .B2(KEYINPUT15), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n274), .A2(G128), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n195), .A2(G143), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G134), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n284), .ZN(new_n407));
  INV_X1    g221(.A(G107), .ZN(new_n408));
  XNOR2_X1  g222(.A(G116), .B(G122), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G122), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G116), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n412), .B2(KEYINPUT14), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT84), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(G116), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n307), .A2(G122), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT14), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n413), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n414), .B1(new_n413), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n410), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n409), .B(new_n408), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT13), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n403), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n404), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n403), .A2(new_n423), .ZN(new_n426));
  OAI21_X1  g240(.A(G134), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n427), .A3(new_n407), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT9), .B(G234), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n429), .A2(new_n256), .A3(G953), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n421), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n421), .B2(new_n428), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n250), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT86), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n421), .A2(new_n428), .ZN(new_n436));
  INV_X1    g250(.A(new_n430), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n431), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n250), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n402), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n401), .B1(new_n434), .B2(KEYINPUT86), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n266), .A2(G143), .A3(G214), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G143), .B1(new_n266), .B2(G214), .ZN(new_n448));
  OAI21_X1  g262(.A(G131), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  INV_X1    g264(.A(G237), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n187), .A3(G214), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n274), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n326), .A3(new_n446), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n449), .A2(new_n450), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n326), .B1(new_n453), .B2(new_n446), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT17), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n224), .A2(new_n455), .A3(new_n228), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n236), .A2(new_n238), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n215), .A2(new_n217), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n459), .B1(new_n210), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(KEYINPUT18), .A2(G131), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n453), .A2(new_n446), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT18), .B(G131), .C1(new_n447), .C2(new_n448), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n461), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(G113), .B(G122), .ZN(new_n466));
  INV_X1    g280(.A(G104), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n458), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT83), .ZN(new_n470));
  INV_X1    g284(.A(new_n454), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n456), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT19), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n237), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n210), .B(new_n474), .C1(new_n460), .C2(new_n473), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n449), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n472), .A2(new_n475), .A3(new_n228), .A4(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n468), .B1(new_n477), .B2(new_n465), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n445), .B1(new_n469), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT20), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n445), .C1(new_n469), .C2(new_n478), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n468), .B1(new_n458), .B2(new_n465), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n250), .B1(new_n469), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n480), .A2(new_n482), .B1(G475), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G952), .ZN(new_n486));
  AOI211_X1 g300(.A(G953), .B(new_n486), .C1(G234), .C2(G237), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT21), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n488), .A2(G898), .ZN(new_n489));
  OAI21_X1  g303(.A(G953), .B1(new_n488), .B2(G898), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n250), .B1(G234), .B2(G237), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n487), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n444), .A2(new_n485), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT87), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n444), .A2(new_n485), .A3(KEYINPUT87), .A4(new_n494), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G214), .B1(G237), .B2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n279), .A2(new_n281), .A3(new_n220), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n220), .B1(new_n301), .B2(new_n303), .ZN(new_n506));
  OAI211_X1 g320(.A(G224), .B(new_n187), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n187), .A2(G224), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n504), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n307), .A2(G119), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT5), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n310), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n306), .A2(new_n308), .A3(KEYINPUT5), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n514), .A2(new_n515), .B1(new_n316), .B2(new_n315), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT3), .B1(new_n467), .B2(G107), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT3), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n408), .A3(G104), .ZN(new_n519));
  INV_X1    g333(.A(G101), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n467), .A2(G107), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n517), .A2(new_n519), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n467), .A2(G107), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n408), .A2(G104), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT77), .B(G101), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G101), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT77), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g342(.A1(new_n516), .A2(new_n522), .A3(new_n525), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(G110), .B(G122), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n517), .A2(new_n519), .A3(new_n521), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G101), .ZN(new_n532));
  AND3_X1   g346(.A1(new_n532), .A2(KEYINPUT4), .A3(new_n522), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT4), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n534), .A3(G101), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n319), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n529), .B(new_n530), .C1(new_n533), .C2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT6), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n529), .B1(new_n533), .B2(new_n536), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n530), .B1(new_n539), .B2(KEYINPUT80), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT80), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n529), .B(new_n541), .C1(new_n533), .C2(new_n536), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(KEYINPUT80), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n545));
  INV_X1    g359(.A(new_n530), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n544), .A2(new_n545), .A3(new_n542), .A4(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT81), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n540), .A2(KEYINPUT81), .A3(new_n545), .A4(new_n542), .ZN(new_n550));
  AOI211_X1 g364(.A(new_n511), .B(new_n543), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n509), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n507), .A2(new_n510), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n528), .A2(new_n522), .A3(new_n525), .ZN(new_n555));
  INV_X1    g369(.A(new_n516), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n529), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n530), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n508), .A2(new_n552), .A3(new_n509), .A4(new_n504), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT82), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n554), .A2(new_n560), .A3(KEYINPUT82), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n537), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n250), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n503), .B1(new_n551), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n565), .A2(new_n537), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n562), .A2(new_n563), .ZN(new_n570));
  AOI21_X1  g384(.A(G902), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n549), .A2(new_n550), .ZN(new_n572));
  INV_X1    g386(.A(new_n511), .ZN(new_n573));
  INV_X1    g387(.A(new_n543), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n571), .A2(new_n575), .A3(new_n502), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n501), .B1(new_n568), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G221), .B1(new_n429), .B2(G902), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT75), .ZN(new_n579));
  INV_X1    g393(.A(G469), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n250), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT79), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n342), .A2(new_n343), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n555), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n555), .B2(new_n583), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT78), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n299), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n273), .A2(KEYINPUT78), .A3(KEYINPUT1), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(G128), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n342), .B1(new_n589), .B2(new_n276), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n555), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n584), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT12), .B1(new_n592), .B2(new_n353), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n282), .A2(new_n535), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n595));
  OAI22_X1  g409(.A1(new_n594), .A2(new_n533), .B1(new_n595), .B2(new_n555), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n590), .A2(new_n555), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n600), .A3(new_n353), .ZN(new_n601));
  INV_X1    g415(.A(new_n585), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n555), .A2(new_n582), .A3(new_n583), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n602), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT12), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n293), .ZN(new_n606));
  XNOR2_X1  g420(.A(G110), .B(G140), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT76), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n187), .A2(G227), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND4_X1  g424(.A1(new_n593), .A2(new_n601), .A3(new_n606), .A4(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n591), .A2(KEYINPUT10), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n293), .B1(new_n612), .B2(new_n596), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n601), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n581), .B1(new_n617), .B2(new_n580), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n585), .A2(new_n591), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n353), .B1(new_n619), .B2(new_n603), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n601), .B1(new_n620), .B2(new_n605), .ZN(new_n621));
  INV_X1    g435(.A(new_n606), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n615), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n601), .A2(new_n613), .A3(new_n610), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n623), .A2(G469), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n579), .B1(new_n618), .B2(new_n625), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n499), .A2(new_n577), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n399), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NAND2_X1  g443(.A1(new_n396), .A2(new_n250), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT88), .A3(G472), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT88), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n369), .A2(new_n371), .ZN(new_n633));
  AOI21_X1  g447(.A(G902), .B1(new_n633), .B2(new_n390), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n632), .B1(new_n634), .B2(new_n376), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n396), .A2(new_n373), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n611), .A2(new_n616), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n580), .A3(new_n250), .ZN(new_n638));
  INV_X1    g452(.A(new_n581), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n639), .A3(new_n625), .ZN(new_n640));
  INV_X1    g454(.A(new_n579), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n264), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n631), .A2(new_n635), .A3(new_n636), .A4(new_n643), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n644), .B(KEYINPUT89), .Z(new_n645));
  OR2_X1    g459(.A1(new_n439), .A2(KEYINPUT33), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n439), .A2(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n647), .A3(G478), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n434), .A2(G478), .ZN(new_n649));
  AND2_X1   g463(.A1(G478), .A2(G902), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n485), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n577), .A2(new_n494), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n645), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT90), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT34), .B(G104), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  NOR3_X1   g473(.A1(new_n551), .A2(new_n567), .A3(new_n503), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n502), .B1(new_n571), .B2(new_n575), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n494), .B(new_n500), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n480), .A2(new_n482), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n484), .A2(G475), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n444), .ZN(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n645), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G107), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G9));
  OR2_X1    g486(.A1(new_n194), .A2(KEYINPUT36), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT92), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(new_n229), .B2(new_n241), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n673), .A2(KEYINPUT92), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(KEYINPUT92), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n676), .A2(new_n247), .A3(new_n240), .A4(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n675), .A2(new_n262), .A3(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n260), .A2(new_n679), .A3(KEYINPUT93), .ZN(new_n680));
  AOI21_X1  g494(.A(KEYINPUT93), .B1(new_n260), .B2(new_n679), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AND4_X1   g496(.A1(new_n499), .A2(new_n682), .A3(new_n577), .A4(new_n626), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n376), .B1(new_n396), .B2(new_n250), .ZN(new_n684));
  AOI22_X1  g498(.A1(new_n684), .A2(KEYINPUT88), .B1(new_n373), .B2(new_n396), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n683), .A2(new_n685), .A3(new_n635), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT37), .B(G110), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  INV_X1    g503(.A(KEYINPUT96), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n187), .A2(G900), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n492), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n693));
  INV_X1    g507(.A(new_n487), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n692), .A2(KEYINPUT95), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n666), .A2(new_n690), .A3(new_n696), .ZN(new_n697));
  OR2_X1    g511(.A1(new_n442), .A2(new_n443), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n485), .A3(new_n696), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n500), .B1(new_n660), .B2(new_n661), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n702), .A3(new_n642), .ZN(new_n703));
  INV_X1    g517(.A(new_n681), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n260), .A2(new_n679), .A3(KEYINPUT93), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n375), .B2(new_n398), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  NAND2_X1  g523(.A1(new_n568), .A2(new_n576), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT38), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT38), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n260), .A2(new_n679), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n322), .A2(new_n383), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n376), .B1(new_n717), .B2(new_n271), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n361), .A2(new_n367), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(G472), .A2(G902), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(KEYINPUT97), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT97), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n719), .A2(new_n723), .A3(new_n720), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n396), .A2(new_n397), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n716), .B1(new_n725), .B2(new_n375), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n500), .B1(new_n442), .B2(new_n443), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n727), .A2(new_n485), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n715), .A2(new_n726), .A3(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT98), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n696), .B(KEYINPUT39), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n626), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n733), .A2(KEYINPUT99), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(KEYINPUT99), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT40), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(KEYINPUT40), .A3(new_n735), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n729), .A2(new_n730), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n731), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT100), .B(G143), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G45));
  INV_X1    g558(.A(new_n388), .ZN(new_n745));
  INV_X1    g559(.A(new_n397), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n372), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT32), .B1(new_n396), .B2(new_n373), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n626), .B(new_n682), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n696), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n485), .A2(new_n652), .A3(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT101), .B1(new_n702), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT101), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n577), .A2(new_n754), .A3(new_n751), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n749), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n210), .ZN(G48));
  NOR2_X1   g572(.A1(new_n617), .A2(new_n580), .ZN(new_n759));
  AOI211_X1 g573(.A(G469), .B(G902), .C1(new_n611), .C2(new_n616), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT102), .B1(new_n761), .B2(new_n641), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n759), .A2(new_n760), .A3(new_n763), .A4(new_n579), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n399), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n655), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT41), .B(G113), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G15));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n668), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G116), .ZN(G18));
  INV_X1    g585(.A(KEYINPUT103), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n637), .A2(new_n250), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(G469), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n641), .A3(new_n638), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n772), .B1(new_n702), .B2(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n759), .A2(new_n760), .A3(new_n579), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(new_n577), .A3(KEYINPUT103), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n779), .A2(new_n707), .A3(new_n499), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT104), .B(G119), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G21));
  OAI211_X1 g596(.A(new_n368), .B(new_n359), .C1(new_n270), .C2(new_n385), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n373), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n786), .B1(new_n634), .B2(new_n376), .ZN(new_n787));
  OAI211_X1 g601(.A(KEYINPUT105), .B(G472), .C1(new_n372), .C2(G902), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n264), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n494), .B(new_n728), .C1(new_n660), .C2(new_n661), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n762), .A2(new_n764), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G122), .ZN(G24));
  INV_X1    g608(.A(new_n716), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n795), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n752), .B1(new_n776), .B2(new_n778), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G125), .ZN(G27));
  INV_X1    g613(.A(KEYINPUT108), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n372), .B2(new_n746), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n396), .A2(KEYINPUT108), .A3(new_n397), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n375), .A3(new_n745), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n624), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n601), .A2(new_n613), .A3(KEYINPUT106), .A4(new_n610), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n623), .A2(G469), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n638), .A2(new_n807), .A3(new_n639), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n641), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n568), .A2(new_n500), .A3(new_n576), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n810), .A3(new_n752), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n803), .A2(KEYINPUT42), .A3(new_n790), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n375), .A2(new_n398), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(new_n811), .A3(KEYINPUT107), .A4(new_n790), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT42), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT107), .B1(new_n399), .B2(new_n811), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G131), .ZN(G33));
  INV_X1    g633(.A(new_n701), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n809), .A2(new_n810), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n813), .A2(new_n790), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G134), .ZN(G36));
  NAND2_X1  g637(.A1(new_n685), .A2(new_n635), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n665), .A2(new_n652), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT43), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT43), .B1(new_n665), .B2(new_n652), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n827), .A2(new_n716), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT44), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n810), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(KEYINPUT44), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT110), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n623), .A2(KEYINPUT45), .A3(new_n805), .A4(new_n806), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n623), .A2(new_n624), .ZN(new_n837));
  OAI211_X1 g651(.A(G469), .B(new_n836), .C1(new_n837), .C2(KEYINPUT45), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT46), .B1(new_n838), .B2(new_n639), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n760), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(KEYINPUT46), .A3(new_n639), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n579), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT109), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n732), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n843), .B1(new_n842), .B2(new_n732), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT110), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n832), .A2(new_n847), .A3(new_n833), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n835), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G137), .ZN(G39));
  INV_X1    g664(.A(KEYINPUT47), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n840), .A2(new_n841), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n579), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n842), .A2(KEYINPUT47), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR4_X1   g669(.A1(new_n813), .A2(new_n790), .A3(new_n752), .A4(new_n810), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(G140), .ZN(G42));
  INV_X1    g672(.A(KEYINPUT51), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n761), .A2(new_n579), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n854), .A3(new_n860), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n789), .A2(new_n790), .ZN(new_n862));
  INV_X1    g676(.A(new_n810), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n827), .A2(new_n487), .A3(new_n828), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n859), .B1(new_n861), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n725), .A2(new_n375), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n775), .A2(new_n810), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n264), .A2(new_n694), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n868), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n485), .A2(new_n652), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT105), .B1(new_n630), .B2(G472), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n634), .A2(new_n786), .A3(new_n376), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n716), .B(new_n784), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n865), .A2(new_n869), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n876), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n500), .B(new_n775), .C1(new_n712), .C2(new_n714), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n862), .A2(new_n865), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT50), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n862), .A2(KEYINPUT50), .A3(new_n865), .A4(new_n882), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n881), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI211_X1 g703(.A(KEYINPUT120), .B(new_n881), .C1(new_n885), .C2(new_n886), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n867), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n862), .A2(new_n779), .A3(new_n865), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n873), .A2(new_n653), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(G952), .A3(new_n187), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n803), .A2(new_n790), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(new_n880), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT48), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(KEYINPUT121), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI211_X1 g714(.A(new_n894), .B(new_n900), .C1(new_n898), .C2(new_n896), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n891), .A2(new_n892), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n885), .A2(new_n886), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT118), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n885), .A2(new_n906), .A3(new_n886), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n881), .B1(new_n861), .B2(new_n866), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n909), .B2(new_n859), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n902), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n399), .B(new_n765), .C1(new_n655), .C2(new_n668), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n912), .A2(new_n793), .A3(new_n780), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n818), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n810), .A2(new_n665), .A3(new_n698), .A4(new_n750), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n707), .A2(new_n626), .A3(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(new_n822), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n631), .A2(new_n636), .A3(new_n635), .ZN(new_n918));
  AOI22_X1  g732(.A1(new_n918), .A2(new_n683), .B1(new_n399), .B2(new_n627), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT113), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n662), .B2(new_n667), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n577), .A2(KEYINPUT113), .A3(new_n494), .A4(new_n666), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n654), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n918), .A2(new_n643), .A3(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n789), .A2(new_n716), .A3(new_n811), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n917), .A2(new_n919), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT114), .B1(new_n914), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT52), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n796), .A2(new_n797), .B1(new_n707), .B2(new_n703), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n696), .B(new_n728), .C1(new_n660), .C2(new_n661), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(new_n809), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n722), .A2(new_n724), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n372), .B2(new_n746), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n931), .B(new_n795), .C1(new_n748), .C2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n749), .B2(new_n756), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT115), .B1(new_n929), .B2(new_n936), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n702), .A2(new_n775), .A3(new_n772), .ZN(new_n938));
  AOI21_X1  g752(.A(KEYINPUT103), .B1(new_n777), .B2(new_n577), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n751), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n708), .B1(new_n879), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT115), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n935), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n928), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n923), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n686), .B(new_n628), .C1(new_n945), .C2(new_n644), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n925), .A2(new_n822), .A3(new_n916), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT114), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n949), .A3(new_n818), .A4(new_n913), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n929), .A2(new_n936), .A3(KEYINPUT115), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n942), .B1(new_n941), .B2(new_n935), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT52), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n927), .A2(new_n944), .A3(new_n950), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT53), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n928), .B1(new_n929), .B2(new_n936), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n951), .A2(new_n952), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n928), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT53), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(new_n959), .A3(new_n950), .A4(new_n927), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n955), .A2(new_n960), .A3(KEYINPUT54), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n954), .A2(new_n959), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT54), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT117), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n914), .B(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT116), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n948), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n926), .A2(KEYINPUT116), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n959), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n958), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n962), .A2(new_n963), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n909), .A2(new_n903), .A3(new_n859), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n911), .A2(new_n961), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(G952), .B2(G953), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n790), .A2(new_n500), .A3(new_n641), .A4(new_n825), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT111), .Z(new_n976));
  XOR2_X1   g790(.A(new_n761), .B(KEYINPUT49), .Z(new_n977));
  NOR4_X1   g791(.A1(new_n976), .A2(new_n868), .A3(new_n715), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(new_n979), .ZN(G75));
  NAND2_X1  g794(.A1(new_n572), .A2(new_n574), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n511), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n575), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(KEYINPUT55), .ZN(new_n984));
  INV_X1    g798(.A(G210), .ZN(new_n985));
  AOI211_X1 g799(.A(new_n985), .B(new_n250), .C1(new_n962), .C2(new_n970), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(KEYINPUT56), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n187), .A2(G952), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n986), .A2(KEYINPUT56), .A3(new_n984), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n990), .A2(new_n991), .ZN(G51));
  XNOR2_X1  g806(.A(new_n581), .B(KEYINPUT57), .ZN(new_n993));
  INV_X1    g807(.A(new_n971), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n963), .B1(new_n962), .B2(new_n970), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n993), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n637), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n250), .B1(new_n962), .B2(new_n970), .ZN(new_n998));
  INV_X1    g812(.A(new_n838), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n988), .B1(new_n997), .B2(new_n1000), .ZN(G54));
  NOR2_X1   g815(.A1(new_n469), .A2(new_n478), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AND2_X1   g817(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(new_n989), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n998), .B2(new_n1004), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT122), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n998), .A2(new_n1004), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n1002), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT122), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1011), .A2(new_n1012), .A3(new_n989), .A4(new_n1006), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1009), .A2(new_n1013), .ZN(G60));
  XNOR2_X1  g828(.A(new_n650), .B(KEYINPUT59), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n961), .B2(new_n971), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n646), .A2(new_n647), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n989), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1015), .B1(new_n646), .B2(new_n647), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n994), .B2(new_n995), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(KEYINPUT123), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT123), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1022), .B(new_n1019), .C1(new_n994), .C2(new_n995), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1018), .B1(new_n1021), .B2(new_n1023), .ZN(G63));
  INV_X1    g838(.A(KEYINPUT61), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G217), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT124), .Z(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT60), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n962), .B2(new_n970), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n678), .A3(new_n675), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(new_n261), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n989), .B1(new_n1029), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1025), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g848(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1035), .A2(KEYINPUT61), .A3(new_n989), .A4(new_n1030), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1034), .A2(new_n1036), .ZN(G66));
  OAI22_X1  g851(.A1(new_n489), .A2(new_n490), .B1(G224), .B2(new_n187), .ZN(new_n1038));
  XOR2_X1   g852(.A(new_n1038), .B(KEYINPUT126), .Z(new_n1039));
  NAND3_X1  g853(.A1(new_n913), .A2(new_n924), .A3(new_n919), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT125), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g857(.A(new_n1039), .B1(new_n1043), .B2(G953), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n981), .B1(G898), .B2(new_n187), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n1044), .B(new_n1045), .ZN(G69));
  NAND2_X1  g860(.A1(new_n362), .A2(new_n345), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n474), .B1(new_n460), .B2(new_n473), .ZN(new_n1048));
  XNOR2_X1  g862(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  NOR4_X1   g863(.A1(new_n895), .A2(new_n485), .A3(new_n711), .A4(new_n727), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1050), .B1(new_n844), .B2(new_n845), .ZN(new_n1051));
  AND4_X1   g865(.A1(new_n818), .A2(new_n857), .A3(new_n822), .A4(new_n1051), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n941), .A2(new_n757), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1052), .A2(new_n849), .A3(new_n1053), .ZN(new_n1054));
  AND2_X1   g868(.A1(new_n1054), .A2(new_n187), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1049), .B1(new_n1055), .B2(new_n691), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n742), .A2(new_n1053), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1057), .B(KEYINPUT62), .ZN(new_n1058));
  OAI211_X1 g872(.A(new_n399), .B(new_n863), .C1(new_n653), .C2(new_n666), .ZN(new_n1059));
  OR2_X1    g873(.A1(new_n1059), .A2(new_n736), .ZN(new_n1060));
  NAND3_X1  g874(.A1(new_n849), .A2(new_n857), .A3(new_n1060), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n187), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1049), .ZN(new_n1063));
  NAND2_X1  g877(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1056), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g879(.A1(G227), .A2(G900), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1065), .A2(G953), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g881(.A1(new_n1066), .A2(G953), .ZN(new_n1068));
  NAND3_X1  g882(.A1(new_n1056), .A2(new_n1068), .A3(new_n1064), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1067), .A2(new_n1069), .ZN(G72));
  INV_X1    g884(.A(new_n380), .ZN(new_n1071));
  NOR2_X1   g885(.A1(new_n1071), .A2(new_n271), .ZN(new_n1072));
  NOR3_X1   g886(.A1(new_n1058), .A2(new_n1061), .A3(new_n1042), .ZN(new_n1073));
  XNOR2_X1  g887(.A(new_n720), .B(KEYINPUT63), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g889(.A(new_n1074), .ZN(new_n1076));
  OAI21_X1  g890(.A(new_n1076), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1077));
  NOR2_X1   g891(.A1(new_n380), .A2(new_n270), .ZN(new_n1078));
  AOI21_X1  g892(.A(new_n988), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n393), .B1(new_n270), .B2(new_n1071), .ZN(new_n1080));
  NAND4_X1  g894(.A1(new_n955), .A2(new_n960), .A3(new_n1076), .A4(new_n1080), .ZN(new_n1081));
  NAND3_X1  g895(.A1(new_n1075), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g896(.A(KEYINPUT127), .ZN(new_n1083));
  NAND2_X1  g897(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g898(.A1(new_n1075), .A2(new_n1079), .A3(KEYINPUT127), .A4(new_n1081), .ZN(new_n1085));
  NAND2_X1  g899(.A1(new_n1084), .A2(new_n1085), .ZN(G57));
endmodule


