//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:00 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  OR2_X1    g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT67), .ZN(G160));
  NAND2_X1  g048(.A1(new_n462), .A2(G136), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n476));
  INV_X1    g051(.A(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n468), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n474), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G162));
  INV_X1    g055(.A(G138), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n482), .B(new_n487), .C1(new_n484), .C2(new_n483), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n464), .B2(G114), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n498));
  AOI211_X1 g073(.A(new_n498), .B(new_n491), .C1(new_n493), .C2(new_n495), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n489), .B(new_n490), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  AND2_X1   g076(.A1(KEYINPUT5), .A2(G543), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n504), .B(KEYINPUT70), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n506), .A2(new_n505), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n502), .A2(new_n503), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n510), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(G543), .B1(new_n506), .B2(new_n505), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G651), .B1(new_n518), .B2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  AND2_X1   g096(.A1(new_n512), .A2(G89), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(G76), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(KEYINPUT71), .B(G51), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n524), .A2(new_n523), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n528), .B1(new_n504), .B2(G63), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n526), .B1(new_n517), .B2(new_n527), .C1(new_n529), .C2(new_n525), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n522), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n512), .A2(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n510), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(new_n518), .B2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n532), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  NAND2_X1  g113(.A1(new_n504), .A2(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n525), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT72), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n512), .A2(G81), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n541), .A2(new_n542), .B1(G43), .B2(new_n518), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  INV_X1    g128(.A(G53), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n517), .A2(KEYINPUT9), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT9), .B1(new_n517), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT74), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n504), .B2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n507), .A2(new_n511), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI221_X1 g137(.A(new_n557), .B1(new_n525), .B2(new_n560), .C1(new_n561), .C2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G168), .ZN(G286));
  NAND2_X1  g139(.A1(new_n512), .A2(G87), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n504), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n566), .A2(G651), .B1(G49), .B2(new_n518), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(G73), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G61), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n510), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n518), .B2(G48), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n561), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g149(.A1(new_n574), .A2(KEYINPUT75), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(KEYINPUT75), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n525), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT76), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n579), .A2(KEYINPUT76), .B1(G47), .B2(new_n518), .ZN(new_n581));
  XNOR2_X1  g156(.A(KEYINPUT77), .B(G85), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n512), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n507), .A2(G92), .A3(new_n511), .ZN(new_n586));
  XOR2_X1   g161(.A(new_n586), .B(KEYINPUT10), .Z(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n510), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n518), .B2(G54), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT78), .ZN(new_n592));
  AND2_X1   g167(.A1(new_n587), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(G168), .B2(new_n596), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(G168), .B2(new_n596), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  XNOR2_X1  g176(.A(new_n546), .B(KEYINPUT73), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n596), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n587), .A2(new_n592), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n596), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n462), .A2(G135), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  INV_X1    g186(.A(G111), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G2105), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n483), .A2(new_n484), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n464), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n613), .B1(new_n615), .B2(G123), .ZN(new_n616));
  AND2_X1   g191(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2096), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n468), .A2(new_n465), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT79), .B(G2100), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n618), .A2(G2096), .ZN(new_n626));
  NAND4_X1  g201(.A1(new_n619), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XOR2_X1   g204(.A(G2427), .B(G2430), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT81), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n631), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n632), .A2(KEYINPUT14), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT82), .Z(new_n642));
  INV_X1    g217(.A(G14), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n639), .B2(new_n640), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT83), .ZN(new_n648));
  NOR2_X1   g223(.A1(G2072), .A2(G2078), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n442), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n648), .A2(new_n650), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n650), .B(KEYINPUT17), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n655), .B(new_n652), .C1(new_n648), .C2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n648), .A2(new_n651), .A3(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n654), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1961), .B(G1966), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1971), .B(G1976), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT19), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n663), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n664), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n670), .B(new_n672), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n667), .A2(new_n668), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT85), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT86), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT89), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(G303), .B2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G1971), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n686), .B1(new_n513), .B2(new_n519), .ZN(new_n692));
  OAI21_X1  g267(.A(G1971), .B1(new_n692), .B2(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n686), .A2(G6), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G305), .B2(G16), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT32), .B(G1981), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n694), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n686), .A2(G23), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(G288), .B2(G16), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n686), .B1(new_n565), .B2(new_n567), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n705), .A2(KEYINPUT33), .A3(new_n701), .ZN(new_n706));
  OAI21_X1  g281(.A(G1976), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(new_n703), .ZN(new_n708));
  INV_X1    g283(.A(G1976), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT33), .B1(new_n705), .B2(new_n701), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n697), .A2(new_n699), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n700), .A2(new_n712), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G25), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n615), .A2(G119), .ZN(new_n718));
  OAI21_X1  g293(.A(KEYINPUT87), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g295(.A1(KEYINPUT87), .A2(G95), .A3(G2105), .ZN(new_n721));
  OAI221_X1 g296(.A(G2104), .B1(G107), .B2(new_n464), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n462), .A2(G131), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n718), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n717), .B1(new_n725), .B2(new_n716), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT35), .B(G1991), .Z(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n726), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1986), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G24), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G290), .A2(KEYINPUT88), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n734));
  NAND4_X1  g309(.A1(new_n580), .A2(new_n581), .A3(new_n734), .A4(new_n583), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n730), .B(new_n732), .C1(new_n736), .C2(new_n686), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n686), .B1(new_n733), .B2(new_n735), .ZN(new_n738));
  OAI21_X1  g313(.A(G1986), .B1(new_n738), .B2(new_n731), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n729), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n715), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(KEYINPUT90), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n715), .A2(new_n743), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n700), .A2(new_n712), .A3(new_n714), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT34), .ZN(new_n747));
  AOI21_X1  g322(.A(KEYINPUT91), .B1(new_n745), .B2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n686), .A2(G19), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n548), .B2(new_n686), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G1341), .ZN(new_n753));
  INV_X1    g328(.A(G1341), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(new_n751), .C1(new_n548), .C2(new_n686), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n716), .A2(G26), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT28), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n462), .A2(G140), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n464), .A2(G116), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G128), .ZN(new_n762));
  OAI221_X1 g337(.A(new_n759), .B1(new_n760), .B2(new_n761), .C1(new_n762), .C2(new_n478), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT92), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n758), .B1(new_n764), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n686), .A2(G4), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n593), .B2(new_n686), .ZN(new_n769));
  INV_X1    g344(.A(G1348), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(G1348), .B(new_n768), .C1(new_n593), .C2(new_n686), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n750), .B1(new_n756), .B2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT97), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n773), .A2(new_n750), .A3(new_n753), .A4(new_n755), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n686), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n686), .ZN(new_n779));
  INV_X1    g354(.A(G1966), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT27), .B(G1996), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT94), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G141), .ZN(new_n786));
  INV_X1    g361(.A(new_n462), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n789), .A2(KEYINPUT26), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(KEYINPUT26), .ZN(new_n791));
  INV_X1    g366(.A(G129), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n790), .B(new_n791), .C1(new_n478), .C2(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(new_n716), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n716), .A2(G32), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n782), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n794), .B(KEYINPUT95), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n798), .B1(new_n800), .B2(G29), .ZN(new_n801));
  INV_X1    g376(.A(new_n782), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n686), .A2(G20), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT23), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G299), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  NOR2_X1   g383(.A1(G164), .A2(new_n716), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G27), .B2(new_n716), .ZN(new_n810));
  INV_X1    g385(.A(G2078), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n781), .A2(new_n804), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n716), .A2(G35), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G162), .B2(new_n716), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT29), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(G2090), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(G2090), .ZN(new_n818));
  NAND2_X1  g393(.A1(G160), .A2(G29), .ZN(new_n819));
  INV_X1    g394(.A(G34), .ZN(new_n820));
  AOI21_X1  g395(.A(G29), .B1(new_n820), .B2(KEYINPUT24), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(KEYINPUT24), .B2(new_n820), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n819), .A2(G2084), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n822), .ZN(new_n824));
  INV_X1    g399(.A(G2084), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n817), .A2(new_n818), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n716), .A2(G33), .ZN(new_n828));
  NAND2_X1  g403(.A1(G115), .A2(G2104), .ZN(new_n829));
  INV_X1    g404(.A(G127), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n614), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G2105), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT25), .Z(new_n834));
  INV_X1    g409(.A(G139), .ZN(new_n835));
  OAI211_X1 g410(.A(new_n832), .B(new_n834), .C1(new_n835), .C2(new_n787), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n828), .B1(new_n837), .B2(new_n716), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(G2072), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(G2072), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT31), .B(G11), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT30), .B(G28), .Z(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(G29), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n617), .B2(G29), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n839), .A2(new_n840), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n686), .A2(G5), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n846), .B1(G301), .B2(G16), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT96), .ZN(new_n848));
  INV_X1    g423(.A(G1961), .ZN(new_n849));
  OR3_X1    g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI22_X1  g425(.A1(new_n810), .A2(new_n811), .B1(new_n847), .B2(new_n849), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n845), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  NOR3_X1   g428(.A1(new_n813), .A2(new_n827), .A3(new_n853), .ZN(new_n854));
  NAND4_X1  g429(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n777), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT97), .B1(new_n856), .B2(new_n774), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n748), .A2(new_n749), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n715), .A2(new_n740), .A3(new_n743), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n743), .B1(new_n715), .B2(new_n740), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n747), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT91), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI211_X1 g438(.A(KEYINPUT91), .B(new_n747), .C1(new_n859), .C2(new_n860), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(KEYINPUT36), .A3(new_n864), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n858), .A2(new_n865), .ZN(G311));
  NAND2_X1  g441(.A1(new_n748), .A2(new_n749), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n855), .A2(new_n857), .ZN(new_n868));
  AND4_X1   g443(.A1(KEYINPUT98), .A2(new_n865), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT98), .B1(new_n858), .B2(new_n865), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(G150));
  AOI22_X1  g446(.A1(new_n512), .A2(G93), .B1(G55), .B2(new_n518), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  INV_X1    g448(.A(G67), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n510), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n525), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n879), .A2(G860), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n602), .A2(new_n879), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n879), .A2(new_n546), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n593), .A2(G559), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n889), .B(KEYINPUT100), .Z(new_n890));
  INV_X1    g465(.A(G860), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(new_n887), .B2(new_n888), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n881), .B1(new_n890), .B2(new_n892), .ZN(G145));
  AND2_X1   g468(.A1(new_n764), .A2(new_n500), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n764), .A2(new_n500), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(new_n796), .ZN(new_n897));
  NOR3_X1   g472(.A1(new_n894), .A2(new_n895), .A3(new_n800), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n837), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(KEYINPUT101), .ZN(new_n900));
  INV_X1    g475(.A(new_n794), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n894), .B2(new_n895), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n836), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n900), .B2(new_n903), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(G130), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n464), .A2(G118), .ZN(new_n909));
  OAI21_X1  g484(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n910));
  OAI22_X1  g485(.A1(new_n478), .A2(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n911), .B1(G142), .B2(new_n462), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(new_n621), .Z(new_n913));
  XOR2_X1   g488(.A(new_n724), .B(KEYINPUT102), .Z(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G160), .B(new_n617), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(new_n479), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n899), .B(new_n915), .C1(new_n905), .C2(new_n906), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT103), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n917), .A2(new_n923), .A3(new_n919), .A4(new_n920), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n919), .B1(new_n917), .B2(new_n920), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(G37), .ZN(new_n927));
  XNOR2_X1  g502(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n925), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n925), .B2(new_n927), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(G395));
  NAND2_X1  g506(.A1(new_n879), .A2(new_n596), .ZN(new_n932));
  XOR2_X1   g507(.A(G305), .B(G290), .Z(new_n933));
  XOR2_X1   g508(.A(G303), .B(G288), .Z(new_n934));
  XNOR2_X1  g509(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n935), .A2(KEYINPUT106), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT42), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n884), .B(new_n605), .Z(new_n938));
  OR3_X1    g513(.A1(new_n593), .A2(KEYINPUT105), .A3(G299), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT105), .B1(new_n593), .B2(G299), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n593), .A2(G299), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT41), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n939), .A2(new_n944), .A3(new_n940), .A4(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n942), .B2(new_n938), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n937), .B(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n932), .B1(new_n949), .B2(new_n596), .ZN(G295));
  OAI21_X1  g525(.A(new_n932), .B1(new_n949), .B2(new_n596), .ZN(G331));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  AOI21_X1  g527(.A(G168), .B1(new_n952), .B2(G301), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(new_n952), .B2(G301), .ZN(new_n954));
  NAND3_X1  g529(.A1(G168), .A2(G171), .A3(KEYINPUT107), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n884), .A2(new_n956), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n882), .A2(new_n883), .B1(new_n954), .B2(new_n955), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n959), .A3(new_n942), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n884), .A2(new_n956), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(new_n958), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n960), .B1(new_n946), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n935), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n960), .B(new_n935), .C1(new_n946), .C2(new_n962), .ZN(new_n966));
  INV_X1    g541(.A(G37), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(new_n966), .A3(new_n970), .A4(new_n967), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT44), .B1(new_n970), .B2(KEYINPUT108), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT109), .Z(new_n973));
  AND3_X1   g548(.A1(new_n969), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n969), .B2(new_n971), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(G1384), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n497), .A2(new_n499), .ZN(new_n978));
  INV_X1    g553(.A(new_n488), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n487), .B1(new_n468), .B2(new_n482), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n490), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n977), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G125), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n470), .B1(new_n614), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G2105), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n987), .A2(G40), .A3(new_n466), .A4(new_n463), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n984), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G1996), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n764), .B(new_n766), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n990), .B1(new_n993), .B2(new_n794), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT47), .Z(new_n996));
  NOR3_X1   g571(.A1(new_n990), .A2(G1986), .A3(G290), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT48), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n901), .A2(G1996), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n993), .B(new_n999), .C1(G1996), .C2(new_n800), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n724), .B(new_n728), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n998), .B1(new_n1002), .B2(new_n990), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n725), .A2(new_n727), .ZN(new_n1004));
  OAI22_X1  g579(.A1(new_n1000), .A2(new_n1004), .B1(G2067), .B2(new_n764), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n989), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n996), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n496), .B(KEYINPUT69), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n486), .A2(new_n488), .B1(new_n615), .B2(G126), .ZN(new_n1010));
  AOI21_X1  g585(.A(G1384), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n988), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n574), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n574), .A2(G1981), .ZN(new_n1018));
  OR3_X1    g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(new_n1013), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G288), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1021), .A2(new_n709), .A3(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1013), .B1(new_n1023), .B2(new_n1018), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1025), .B(KEYINPUT55), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n983), .A2(G1384), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n988), .B1(new_n500), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n984), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n690), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT110), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n988), .B1(new_n982), .B2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1034), .B(new_n977), .C1(new_n978), .C2(new_n981), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(G2090), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1031), .A2(KEYINPUT110), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1027), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1013), .B1(new_n709), .B2(G288), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1022), .A2(G1976), .ZN(new_n1041));
  OR3_X1    g616(.A1(new_n1040), .A2(new_n1041), .A3(KEYINPUT52), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1042), .A2(new_n1021), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1024), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1044), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1046), .A2(new_n1039), .ZN(new_n1047));
  OAI21_X1  g622(.A(G8), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n1026), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1028), .B1(new_n978), .B2(new_n981), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1012), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT45), .B1(new_n500), .B2(new_n977), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n780), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1030), .A2(KEYINPUT112), .A3(new_n780), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1012), .B1(new_n1011), .B2(new_n1034), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1035), .A2(new_n825), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT113), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(G2084), .B1(new_n1011), .B2(new_n1034), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1033), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1060), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1008), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(G168), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1047), .A2(new_n1049), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT111), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1011), .A2(new_n1070), .A3(new_n1034), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1033), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1031), .B1(new_n1073), .B2(G2090), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(G8), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(new_n1026), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1046), .A2(new_n1039), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1067), .B1(new_n1077), .B2(new_n1066), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1045), .B1(new_n1069), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1057), .A2(new_n1080), .A3(new_n1064), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1057), .B2(new_n1064), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G168), .A2(new_n1008), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT118), .B(KEYINPUT51), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(G8), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1085), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT112), .B1(new_n1030), .B2(new_n780), .ZN(new_n1092));
  AOI211_X1 g667(.A(new_n1054), .B(G1966), .C1(new_n984), .C2(new_n1029), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1058), .A2(new_n1059), .A3(KEYINPUT113), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1062), .B1(new_n1061), .B2(new_n1033), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1092), .A2(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT117), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1057), .A2(new_n1080), .A3(new_n1064), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1089), .B1(new_n1099), .B2(G8), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1088), .B1(new_n1091), .B2(new_n1100), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1065), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1065), .A2(KEYINPUT120), .A3(new_n1102), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1086), .B1(new_n1101), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1030), .B2(G1996), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n548), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT59), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n548), .A2(new_n1115), .A3(new_n1112), .ZN(new_n1116));
  AOI21_X1  g691(.A(G1348), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1109), .A2(G2067), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n604), .A2(KEYINPUT60), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1114), .A2(new_n1116), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1122));
  INV_X1    g697(.A(G1956), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1073), .A2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT57), .B1(new_n557), .B2(KEYINPUT114), .ZN(new_n1125));
  XNOR2_X1  g700(.A(G299), .B(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n984), .A2(new_n1029), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT116), .B1(KEYINPUT115), .B2(KEYINPUT61), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND4_X1   g708(.A1(new_n1122), .A2(new_n1129), .A3(new_n1130), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1036), .A2(new_n770), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1118), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n604), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n593), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1141), .B2(KEYINPUT60), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1121), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1126), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1140), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1144), .B1(new_n1145), .B2(new_n1129), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1077), .B1(new_n1143), .B2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n1030), .B2(G2078), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n984), .A2(new_n1029), .A3(KEYINPUT53), .A4(new_n811), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(G1961), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT122), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1035), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n849), .B1(new_n1058), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(new_n1159), .A3(new_n1153), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1152), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1149), .B1(new_n1161), .B2(G301), .ZN(new_n1162));
  NOR3_X1   g737(.A1(new_n1154), .A2(new_n1155), .A3(KEYINPUT122), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1159), .B1(new_n1158), .B2(new_n1153), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1151), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1162), .A2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1151), .A2(new_n1158), .A3(new_n1153), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1168), .A2(G171), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1148), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1171), .B1(new_n1165), .B2(G171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1161), .A2(KEYINPUT125), .A3(G301), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT126), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1151), .A2(KEYINPUT126), .A3(new_n1158), .A4(new_n1153), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1176), .A2(G171), .A3(new_n1177), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1178), .A2(KEYINPUT127), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT54), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1180), .B1(new_n1178), .B2(KEYINPUT127), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1174), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1147), .A2(new_n1170), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1079), .B1(new_n1108), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1047), .A2(new_n1167), .A3(new_n1076), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1086), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1008), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1084), .B1(new_n1187), .B2(new_n1089), .ZN(new_n1188));
  OAI21_X1  g763(.A(KEYINPUT119), .B1(new_n1083), .B2(new_n1008), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1087), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1186), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1185), .B1(new_n1192), .B2(KEYINPUT62), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1108), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1184), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g771(.A(G290), .B(new_n730), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n990), .B1(new_n1002), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1007), .B1(new_n1196), .B2(new_n1198), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g774(.A(G319), .ZN(new_n1201));
  NOR2_X1   g775(.A1(G227), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n645), .A2(new_n684), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g777(.A(new_n1203), .B1(new_n925), .B2(new_n927), .ZN(new_n1204));
  NAND2_X1  g778(.A1(new_n969), .A2(new_n971), .ZN(new_n1205));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1205), .ZN(G225));
  INV_X1    g780(.A(G225), .ZN(G308));
endmodule


