//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(G146), .C1(new_n188), .C2(KEYINPUT1), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n188), .A2(new_n190), .A3(G143), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n191), .A2(new_n193), .A3(new_n200), .ZN(new_n201));
  XNOR2_X1  g015(.A(G143), .B(G146), .ZN(new_n202));
  XNOR2_X1  g016(.A(KEYINPUT0), .B(G128), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n201), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n199), .B1(new_n198), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G224), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(G953), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n207), .B(KEYINPUT83), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n205), .B(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT76), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(G104), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT76), .B1(new_n213), .B2(G107), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n211), .A2(G104), .ZN(new_n215));
  OAI211_X1 g029(.A(G101), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n211), .A3(G104), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n213), .A2(G107), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G116), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT65), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G116), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n227), .A3(G119), .ZN(new_n228));
  INV_X1    g042(.A(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G116), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(KEYINPUT5), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n230), .A2(KEYINPUT5), .ZN(new_n232));
  INV_X1    g046(.A(G113), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(KEYINPUT2), .B(G113), .Z(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n228), .A3(new_n230), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n223), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n217), .A2(new_n219), .A3(new_n221), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(G101), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n239), .A2(G101), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n222), .A2(KEYINPUT4), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n237), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n236), .B1(new_n230), .B2(new_n228), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n238), .B1(new_n244), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT82), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n238), .B(KEYINPUT82), .C1(new_n244), .C2(new_n247), .ZN(new_n251));
  XNOR2_X1  g065(.A(G110), .B(G122), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n238), .B(new_n252), .C1(new_n244), .C2(new_n247), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT6), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n252), .B1(new_n248), .B2(new_n249), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n258), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n209), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(G210), .B1(G237), .B2(G902), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT7), .B1(new_n206), .B2(G953), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n205), .B(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n235), .A2(new_n237), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(new_n223), .ZN(new_n266));
  XOR2_X1   g080(.A(new_n252), .B(KEYINPUT8), .Z(new_n267));
  OAI211_X1 g081(.A(new_n264), .B(new_n255), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n260), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n209), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n258), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n258), .A2(new_n251), .B1(KEYINPUT6), .B2(new_n255), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n270), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n261), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(G128), .B(G143), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n225), .A2(new_n227), .A3(G122), .ZN(new_n283));
  OR2_X1    g097(.A1(new_n224), .A2(G122), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n285), .A2(KEYINPUT14), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT14), .ZN(new_n287));
  OAI21_X1  g101(.A(G107), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  OAI221_X1 g102(.A(new_n282), .B1(G107), .B2(new_n285), .C1(new_n286), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(KEYINPUT87), .C1(G128), .C2(new_n192), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT13), .B1(new_n192), .B2(G128), .ZN(new_n292));
  OAI221_X1 g106(.A(G134), .B1(KEYINPUT87), .B2(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n280), .A2(new_n281), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n211), .B1(new_n283), .B2(new_n284), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n285), .A2(G107), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  INV_X1    g112(.A(G217), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n298), .A2(new_n299), .A3(G953), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n289), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n300), .B1(new_n289), .B2(new_n297), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  OR3_X1    g119(.A1(new_n303), .A2(G902), .A3(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n305), .B1(new_n303), .B2(G902), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G952), .ZN(new_n309));
  AOI211_X1 g123(.A(G953), .B(new_n309), .C1(G234), .C2(G237), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(KEYINPUT67), .A2(G953), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT67), .A2(G953), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n269), .B1(G234), .B2(G237), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT21), .B(G898), .Z(new_n319));
  OAI21_X1  g133(.A(new_n311), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n320), .B(KEYINPUT88), .Z(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n308), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(KEYINPUT67), .A2(G953), .ZN(new_n324));
  INV_X1    g138(.A(G237), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT67), .A2(G953), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(G214), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT84), .B(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  OR2_X1    g143(.A1(KEYINPUT84), .A2(G143), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n314), .A2(G214), .A3(new_n325), .A4(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G131), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT17), .ZN(new_n334));
  INV_X1    g148(.A(G131), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n329), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT74), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n198), .A3(G140), .ZN(new_n339));
  INV_X1    g153(.A(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G125), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n198), .A2(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT16), .B(new_n339), .C1(new_n343), .C2(new_n338), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT16), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n190), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n332), .A2(KEYINPUT17), .A3(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n190), .A3(new_n346), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT18), .ZN(new_n352));
  AOI211_X1 g166(.A(new_n352), .B(new_n335), .C1(new_n329), .C2(new_n331), .ZN(new_n353));
  NAND2_X1  g167(.A1(KEYINPUT18), .A2(G131), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n329), .A2(new_n331), .A3(new_n354), .ZN(new_n355));
  OAI211_X1 g169(.A(G146), .B(new_n339), .C1(new_n343), .C2(new_n338), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n341), .A2(new_n342), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n190), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT85), .B1(new_n353), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n332), .A2(KEYINPUT18), .A3(G131), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT85), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n362), .A2(new_n363), .A3(new_n355), .A4(new_n359), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n337), .A2(new_n351), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(G113), .B(G122), .ZN(new_n366));
  XNOR2_X1  g180(.A(new_n366), .B(new_n213), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n361), .A2(new_n364), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n337), .A2(new_n350), .A3(new_n348), .A4(new_n349), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT86), .A4(new_n367), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n368), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(G475), .B1(new_n375), .B2(G902), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT20), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n333), .A2(new_n336), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n357), .A2(KEYINPUT19), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n339), .B1(new_n343), .B2(new_n338), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n379), .B1(new_n380), .B2(KEYINPUT19), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n378), .B(new_n348), .C1(G146), .C2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n367), .B1(new_n369), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT86), .B1(new_n365), .B2(new_n367), .ZN(new_n385));
  INV_X1    g199(.A(new_n374), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n377), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n383), .B1(new_n373), .B2(new_n374), .ZN(new_n390));
  INV_X1    g204(.A(new_n388), .ZN(new_n391));
  NOR3_X1   g205(.A1(new_n390), .A2(KEYINPUT20), .A3(new_n391), .ZN(new_n392));
  OAI211_X1 g206(.A(new_n323), .B(new_n376), .C1(new_n389), .C2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT81), .ZN(new_n395));
  OAI21_X1  g209(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G469), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n269), .ZN(new_n399));
  INV_X1    g213(.A(new_n204), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(new_n241), .C1(new_n242), .C2(new_n243), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n197), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n216), .A2(new_n222), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n195), .A2(new_n196), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(KEYINPUT77), .B2(new_n194), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT77), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n202), .A2(new_n406), .A3(new_n189), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n403), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n401), .B(new_n402), .C1(new_n408), .C2(KEYINPUT10), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT11), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n281), .B2(G137), .ZN(new_n411));
  INV_X1    g225(.A(G137), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT11), .A3(G134), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n281), .A2(G137), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G131), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n411), .A2(new_n413), .A3(new_n335), .A4(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT78), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT79), .B1(new_n409), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n194), .A2(KEYINPUT77), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n421), .A2(new_n407), .A3(new_n195), .A4(new_n196), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n223), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT10), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n197), .A2(KEYINPUT10), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n423), .A2(new_n424), .B1(new_n425), .B2(new_n223), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n418), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT79), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n426), .A2(new_n428), .A3(new_n429), .A4(new_n401), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT80), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n416), .B2(new_n417), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n197), .B1(new_n222), .B2(new_n216), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n433), .B1(new_n408), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT12), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT12), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n433), .C1(new_n408), .C2(new_n434), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n431), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n314), .A2(G227), .ZN(new_n442));
  XOR2_X1   g256(.A(G110), .B(G140), .Z(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n420), .B2(new_n430), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n409), .A2(new_n418), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n441), .A2(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n399), .B1(new_n447), .B2(G469), .ZN(new_n448));
  INV_X1    g262(.A(new_n444), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n431), .A2(new_n440), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n449), .B1(new_n431), .B2(new_n446), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n398), .B(new_n269), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n395), .B(new_n397), .C1(new_n448), .C2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n431), .A2(new_n446), .A3(new_n449), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n439), .B1(new_n430), .B2(new_n420), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n454), .B(G469), .C1(new_n449), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n399), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n452), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT81), .B1(new_n458), .B2(new_n396), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n279), .B(new_n394), .C1(new_n453), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n188), .A2(G119), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n229), .A2(G128), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT24), .B(G110), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT23), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n229), .B2(G128), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n463), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n470), .A2(KEYINPUT73), .ZN(new_n471));
  INV_X1    g285(.A(G110), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n470), .B2(KEYINPUT73), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n466), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n350), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n474), .B1(new_n475), .B2(new_n347), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(new_n465), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n477), .B1(new_n470), .B2(G110), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n348), .A2(new_n358), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n314), .A2(G221), .A3(G234), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT22), .B(G137), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n476), .A2(new_n479), .A3(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n269), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT25), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n485), .A2(KEYINPUT25), .A3(new_n269), .A4(new_n486), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n299), .B1(G234), .B2(new_n269), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n485), .A2(new_n486), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n492), .A2(G902), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT75), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(G472), .A2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT26), .B(G101), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n314), .A2(G210), .A3(new_n325), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT27), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n503), .A2(KEYINPUT27), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n504), .A3(new_n501), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n511));
  INV_X1    g325(.A(new_n247), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n281), .A2(G137), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n412), .A2(G134), .ZN(new_n514));
  OAI21_X1  g328(.A(G131), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n189), .A2(new_n191), .A3(new_n193), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n417), .B(new_n515), .C1(new_n516), .C2(new_n404), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n204), .B1(new_n417), .B2(new_n416), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT64), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n418), .A2(new_n519), .A3(new_n400), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n418), .A2(new_n400), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n418), .A2(KEYINPUT66), .A3(new_n400), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n525), .A2(new_n247), .A3(new_n517), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n511), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n228), .A2(new_n230), .ZN(new_n529));
  INV_X1    g343(.A(new_n236), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n517), .A2(new_n531), .A3(new_n237), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n511), .B1(new_n532), .B2(new_n518), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT68), .B(new_n511), .C1(new_n532), .C2(new_n518), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n510), .B1(new_n528), .B2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n539), .B1(new_n520), .B2(new_n521), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n525), .A2(KEYINPUT30), .A3(new_n517), .A4(new_n526), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n512), .A3(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n418), .A2(KEYINPUT66), .A3(new_n400), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT66), .B1(new_n418), .B2(new_n400), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n543), .A2(new_n544), .A3(new_n532), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n542), .A2(KEYINPUT31), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(KEYINPUT31), .B1(new_n542), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n538), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT69), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(KEYINPUT69), .B(new_n538), .C1(new_n547), .C2(new_n548), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n500), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n535), .A2(new_n536), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n510), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n525), .A2(new_n517), .A3(new_n526), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n545), .B1(new_n512), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n554), .B(new_n556), .C1(new_n558), .C2(new_n511), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n557), .A2(new_n512), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n527), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT28), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n564), .A2(KEYINPUT72), .A3(new_n554), .A4(new_n556), .ZN(new_n565));
  AOI21_X1  g379(.A(G902), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n542), .A2(new_n527), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(new_n510), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT71), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n528), .A2(new_n537), .ZN(new_n570));
  INV_X1    g384(.A(new_n510), .ZN(new_n571));
  AOI21_X1  g385(.A(KEYINPUT29), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT71), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n567), .A2(new_n573), .A3(new_n510), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n566), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n553), .A2(KEYINPUT32), .B1(new_n576), .B2(G472), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n542), .A2(new_n546), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT31), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n542), .A2(KEYINPUT31), .A3(new_n546), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(KEYINPUT69), .B1(new_n582), .B2(new_n538), .ZN(new_n583));
  INV_X1    g397(.A(new_n552), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n499), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n498), .B1(new_n577), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n461), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  OAI21_X1  g405(.A(new_n279), .B1(new_n453), .B2(new_n459), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n498), .A2(new_n322), .ZN(new_n593));
  INV_X1    g407(.A(G472), .ZN(new_n594));
  AOI21_X1  g408(.A(G902), .B1(new_n551), .B2(new_n552), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n593), .B(new_n585), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n303), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n303), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n601), .A3(G478), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n304), .A3(new_n269), .ZN(new_n603));
  NAND2_X1  g417(.A1(G478), .A2(G902), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n387), .A2(new_n377), .A3(new_n388), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT20), .B1(new_n390), .B2(new_n391), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI211_X1 g422(.A(KEYINPUT89), .B(new_n605), .C1(new_n608), .C2(new_n376), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT89), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n376), .B1(new_n389), .B2(new_n392), .ZN(new_n611));
  INV_X1    g425(.A(new_n605), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n597), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT90), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT34), .B(G104), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n606), .A2(new_n607), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n389), .A2(KEYINPUT91), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n376), .A4(new_n308), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n592), .A2(new_n596), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(KEYINPUT35), .B(G107), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  OAI21_X1  g440(.A(new_n480), .B1(KEYINPUT36), .B2(new_n484), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n476), .A2(new_n479), .A3(new_n628), .A4(new_n483), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n496), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT92), .ZN(new_n631));
  INV_X1    g445(.A(new_n492), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n632), .B1(new_n489), .B2(new_n490), .ZN(new_n633));
  OAI21_X1  g447(.A(KEYINPUT93), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT92), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n630), .B(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT93), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n493), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n639), .B(new_n585), .C1(new_n594), .C2(new_n595), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n460), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT37), .B(G110), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  NAND2_X1  g457(.A1(new_n634), .A2(new_n638), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n577), .B2(new_n588), .ZN(new_n645));
  INV_X1    g459(.A(new_n452), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n456), .A2(new_n457), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n396), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n395), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n458), .A2(KEYINPUT81), .A3(new_n396), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n278), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(G900), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n310), .B1(new_n317), .B2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n623), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n645), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT94), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n645), .A2(new_n651), .A3(new_n657), .A4(new_n654), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT95), .B(G128), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G30));
  NAND2_X1  g475(.A1(new_n649), .A2(new_n650), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n653), .B(KEYINPUT39), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n271), .A2(new_n277), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT38), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(KEYINPUT32), .B(new_n499), .C1(new_n583), .C2(new_n584), .ZN(new_n669));
  INV_X1    g483(.A(new_n578), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n563), .A2(new_n510), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(KEYINPUT96), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n671), .A2(KEYINPUT96), .ZN(new_n673));
  AOI21_X1  g487(.A(G902), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n588), .B(new_n669), .C1(new_n594), .C2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n493), .A2(new_n636), .ZN(new_n676));
  INV_X1    g490(.A(new_n187), .ZN(new_n677));
  INV_X1    g491(.A(new_n308), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n611), .A2(new_n668), .A3(new_n675), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n664), .A2(KEYINPUT40), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n665), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  INV_X1    g497(.A(new_n653), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n611), .A2(new_n612), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n645), .A2(new_n651), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT97), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n645), .A2(new_n651), .A3(KEYINPUT97), .A4(new_n686), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NOR2_X1   g506(.A1(new_n278), .A2(new_n322), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n609), .B2(new_n613), .ZN(new_n694));
  INV_X1    g508(.A(new_n498), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n431), .A2(new_n446), .ZN(new_n696));
  AOI22_X1  g510(.A1(new_n696), .A2(new_n444), .B1(new_n445), .B2(new_n440), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n396), .A3(new_n452), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n537), .B1(new_n563), .B2(KEYINPUT28), .ZN(new_n701));
  AOI21_X1  g515(.A(KEYINPUT72), .B1(new_n701), .B2(new_n556), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n511), .B1(new_n562), .B2(new_n527), .ZN(new_n703));
  INV_X1    g517(.A(new_n556), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n703), .A2(new_n704), .A3(new_n537), .A4(new_n560), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n269), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n517), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n523), .B2(KEYINPUT64), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n518), .A2(new_n519), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n247), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT28), .B1(new_n710), .B2(new_n545), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(new_n554), .A3(new_n571), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n555), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n573), .B1(new_n567), .B2(new_n510), .ZN(new_n714));
  AOI211_X1 g528(.A(KEYINPUT71), .B(new_n571), .C1(new_n542), .C2(new_n527), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n669), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n553), .A2(new_n586), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n695), .B(new_n700), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n694), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NOR3_X1   g537(.A1(new_n623), .A2(new_n278), .A3(new_n322), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n589), .A2(new_n724), .A3(new_n700), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  OAI211_X1 g540(.A(new_n669), .B(new_n717), .C1(new_n553), .C2(new_n586), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n699), .A2(new_n278), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n394), .A3(new_n639), .A4(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NOR3_X1   g544(.A1(new_n699), .A2(new_n278), .A3(new_n322), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n269), .B1(new_n583), .B2(new_n584), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n582), .B1(new_n571), .B2(new_n701), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n732), .A2(G472), .B1(new_n499), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n678), .B1(new_n608), .B2(new_n376), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n731), .A2(new_n734), .A3(new_n695), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  NAND2_X1  g551(.A1(new_n733), .A2(new_n499), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(new_n676), .C1(new_n595), .C2(new_n594), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n686), .A3(new_n728), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G125), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n456), .A2(KEYINPUT98), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n441), .A2(new_n444), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT98), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n746), .A3(G469), .A4(new_n454), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n744), .A2(new_n452), .A3(new_n457), .A4(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n262), .B1(new_n260), .B2(new_n270), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n275), .A2(new_n261), .A3(new_n276), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n187), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n751), .A3(new_n396), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT99), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT99), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n748), .A2(new_n751), .A3(new_n754), .A4(new_n396), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n685), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n553), .A2(KEYINPUT32), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n498), .B1(new_n757), .B2(new_n577), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n743), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n755), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n760), .A2(new_n589), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT100), .B(G131), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G33));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n589), .A3(new_n654), .ZN(new_n766));
  XOR2_X1   g580(.A(KEYINPUT101), .B(G134), .Z(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G36));
  OR2_X1    g582(.A1(new_n447), .A2(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n447), .A2(KEYINPUT45), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(G469), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT102), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n399), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n452), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n396), .B(new_n663), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  INV_X1    g592(.A(new_n611), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n612), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT43), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n780), .B1(KEYINPUT103), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n782), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT104), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n595), .A2(new_n594), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n553), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n789), .B1(new_n493), .B2(new_n636), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n777), .B1(new_n778), .B2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n751), .B(KEYINPUT105), .Z(new_n793));
  OAI211_X1 g607(.A(new_n792), .B(new_n793), .C1(new_n778), .C2(new_n791), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  OAI21_X1  g609(.A(new_n396), .B1(new_n775), .B2(new_n776), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT47), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g612(.A(KEYINPUT47), .B(new_n396), .C1(new_n775), .C2(new_n776), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n751), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n727), .A2(new_n685), .A3(new_n695), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(KEYINPUT106), .B(G140), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n803), .B(new_n804), .ZN(G42));
  NAND3_X1  g619(.A1(new_n695), .A2(new_n396), .A3(new_n187), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n698), .A2(new_n452), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n806), .B(new_n780), .C1(KEYINPUT49), .C2(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT107), .Z(new_n809));
  NOR2_X1   g623(.A1(new_n807), .A2(KEYINPUT49), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(KEYINPUT108), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n667), .B1(new_n813), .B2(new_n810), .ZN(new_n814));
  OR4_X1    g628(.A1(new_n675), .A2(new_n809), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n668), .A2(new_n187), .A3(new_n699), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n734), .A2(new_n695), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n784), .A2(new_n816), .A3(new_n310), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT50), .B1(new_n819), .B2(KEYINPUT115), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT116), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n822), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n825), .A3(new_n820), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n801), .A2(new_n311), .A3(new_n699), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n784), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n740), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n695), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n675), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n779), .A3(new_n605), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n698), .A2(new_n397), .A3(new_n452), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n798), .A2(new_n799), .A3(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n784), .A2(new_n310), .A3(new_n818), .A4(new_n793), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT114), .Z(new_n838));
  AOI21_X1  g652(.A(new_n834), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n827), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n829), .A2(new_n758), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(KEYINPUT48), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n784), .A2(new_n310), .A3(new_n728), .A4(new_n818), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n309), .B(G953), .C1(new_n832), .C2(new_n615), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n821), .A2(new_n841), .A3(new_n822), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n839), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT51), .B1(new_n827), .B2(new_n839), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n836), .A2(new_n838), .ZN(new_n853));
  INV_X1    g667(.A(new_n834), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n849), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT117), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT53), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n779), .A2(new_n308), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n592), .A2(new_n596), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT109), .B1(new_n862), .B2(new_n641), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n611), .A2(new_n612), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n597), .A2(new_n865), .B1(new_n461), .B2(new_n589), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n651), .A2(new_n394), .A3(new_n789), .A4(new_n639), .ZN(new_n867));
  INV_X1    g681(.A(new_n596), .ZN(new_n868));
  INV_X1    g682(.A(new_n861), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n651), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT109), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n863), .A2(new_n866), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n760), .A2(new_n686), .A3(new_n740), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n376), .A2(new_n678), .A3(new_n684), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n801), .A2(new_n644), .A3(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n621), .A2(new_n622), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(new_n662), .A3(new_n727), .A4(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n766), .A2(new_n874), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n748), .A2(new_n396), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n735), .A2(new_n279), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n676), .A2(new_n653), .ZN(new_n883));
  AND4_X1   g697(.A1(new_n675), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n884), .B1(new_n689), .B2(new_n690), .ZN(new_n885));
  INV_X1    g699(.A(new_n741), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n656), .B2(new_n658), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT52), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n759), .A2(new_n762), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n721), .A2(new_n725), .A3(new_n729), .A4(new_n736), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n880), .A2(new_n889), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n885), .B2(new_n887), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n860), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n729), .B(new_n736), .C1(new_n694), .C2(new_n720), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n589), .A2(new_n700), .A3(new_n724), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n763), .A2(new_n898), .A3(KEYINPUT53), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n766), .A2(new_n874), .A3(new_n878), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n872), .A3(new_n863), .A4(new_n866), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT112), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n885), .A2(new_n887), .ZN(new_n904));
  XOR2_X1   g718(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n863), .A2(new_n866), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n907), .A2(KEYINPUT112), .A3(new_n872), .A4(new_n900), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(new_n889), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT54), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n895), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n906), .A2(new_n889), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n880), .A2(new_n892), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT110), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n880), .A2(new_n892), .A3(KEYINPUT110), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n912), .A2(new_n915), .A3(new_n860), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n904), .A2(KEYINPUT52), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(new_n892), .A3(new_n880), .A4(new_n889), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n917), .B1(new_n860), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n911), .B1(new_n921), .B2(new_n910), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT113), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT113), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n924), .B(new_n911), .C1(new_n921), .C2(new_n910), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n859), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n815), .B1(new_n926), .B2(new_n927), .ZN(G75));
  NOR2_X1   g742(.A1(new_n314), .A2(G952), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n895), .A2(new_n909), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT56), .B1(new_n933), .B2(G210), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n273), .A2(new_n274), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n209), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n275), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT119), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n930), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n941), .B1(new_n934), .B2(new_n940), .ZN(G51));
  INV_X1    g756(.A(new_n773), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT121), .B1(new_n932), .B2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT121), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n931), .A2(new_n945), .A3(G902), .A4(new_n773), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT120), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n931), .A2(KEYINPUT54), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n911), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n399), .B(KEYINPUT57), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n697), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n947), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n697), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n949), .A2(new_n911), .ZN(new_n955));
  INV_X1    g769(.A(new_n951), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT120), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n929), .B1(new_n953), .B2(new_n958), .ZN(G54));
  NAND3_X1  g773(.A1(new_n933), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n390), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n390), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n929), .ZN(G60));
  AND2_X1   g777(.A1(new_n599), .A2(new_n601), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n604), .B(KEYINPUT59), .Z(new_n965));
  OR2_X1    g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n930), .B1(new_n955), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n965), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n923), .A2(new_n925), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n967), .B1(new_n969), .B2(new_n964), .ZN(G63));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n895), .B2(new_n909), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n627), .A2(new_n629), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n929), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  INV_X1    g790(.A(new_n494), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n901), .A2(new_n902), .ZN(new_n978));
  INV_X1    g792(.A(new_n899), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n908), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI22_X1  g794(.A1(new_n980), .A2(new_n912), .B1(new_n919), .B2(new_n860), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n981), .B2(new_n972), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n975), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n976), .B1(new_n975), .B2(new_n982), .ZN(new_n984));
  INV_X1    g798(.A(new_n972), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n931), .A2(new_n974), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(KEYINPUT122), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT61), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n983), .A2(new_n984), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT61), .B1(new_n986), .B2(KEYINPUT122), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n986), .A2(new_n930), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n973), .A2(new_n494), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT123), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n975), .A2(new_n982), .A3(new_n976), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n991), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n990), .A2(new_n996), .ZN(G66));
  NOR2_X1   g811(.A1(new_n873), .A2(new_n891), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n998), .B(KEYINPUT124), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n319), .A2(G224), .ZN(new_n1000));
  AOI22_X1  g814(.A1(new_n999), .A2(new_n314), .B1(G953), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n935), .B1(G898), .B2(new_n314), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1001), .B(new_n1002), .Z(G69));
  NAND2_X1  g817(.A1(new_n540), .A2(new_n541), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(new_n381), .Z(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT125), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n801), .B1(new_n861), .B2(new_n864), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n589), .A3(new_n662), .A4(new_n663), .ZN(new_n1008));
  AND2_X1   g822(.A1(new_n794), .A2(new_n1008), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n887), .A2(new_n691), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n682), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1011), .A2(KEYINPUT62), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(KEYINPUT62), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1009), .A2(new_n803), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1006), .B1(new_n1014), .B2(new_n314), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n314), .B1(G227), .B2(G900), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n763), .A2(new_n766), .ZN(new_n1017));
  INV_X1    g831(.A(new_n777), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n758), .A2(new_n882), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n794), .A2(new_n1020), .A3(new_n803), .A4(new_n1010), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n315), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1005), .B1(G900), .B2(new_n315), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  OR3_X1    g839(.A1(new_n1015), .A2(new_n1016), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1016), .B1(new_n1015), .B2(new_n1025), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(G72));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT63), .ZN(new_n1030));
  XOR2_X1   g844(.A(new_n1030), .B(KEYINPUT126), .Z(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n1014), .B2(new_n999), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1032), .A2(new_n571), .A3(new_n567), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n714), .A2(new_n715), .A3(new_n670), .ZN(new_n1034));
  OR3_X1    g848(.A1(new_n921), .A2(new_n1030), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1031), .B1(new_n1021), .B2(new_n999), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n567), .A2(new_n571), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT127), .Z(new_n1038));
  AOI21_X1  g852(.A(new_n929), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1033), .A2(new_n1035), .A3(new_n1039), .ZN(G57));
endmodule


