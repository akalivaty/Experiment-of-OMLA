//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT66), .ZN(new_n203));
  OAI22_X1  g002(.A1(new_n202), .A2(KEYINPUT24), .B1(new_n203), .B2(KEYINPUT25), .ZN(new_n204));
  XOR2_X1   g003(.A(G183gat), .B(G190gat), .Z(new_n205));
  AOI21_X1  g004(.A(new_n204), .B1(new_n205), .B2(KEYINPUT24), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT65), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(KEYINPUT25), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n212), .B(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT26), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n221), .A2(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n219), .A2(KEYINPUT67), .A3(new_n222), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n214), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT70), .ZN(new_n228));
  XOR2_X1   g027(.A(G113gat), .B(G120gat), .Z(new_n229));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G127gat), .ZN(new_n232));
  INV_X1    g031(.A(G127gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G134gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n229), .B(new_n230), .C1(KEYINPUT69), .C2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  INV_X1    g036(.A(new_n235), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n237), .ZN(new_n240));
  XNOR2_X1  g039(.A(G113gat), .B(G120gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT69), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT1), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n228), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n240), .A2(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n238), .A2(new_n242), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n241), .A2(KEYINPUT1), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n247), .A2(new_n248), .B1(KEYINPUT68), .B2(new_n235), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n249), .A3(KEYINPUT70), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n227), .A2(new_n251), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n245), .A2(new_n250), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n253), .A2(new_n214), .A3(new_n225), .A4(new_n226), .ZN(new_n254));
  INV_X1    g053(.A(G227gat), .ZN(new_n255));
  INV_X1    g054(.A(G233gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(new_n254), .A3(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT34), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n252), .B2(new_n254), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT32), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n262), .A2(KEYINPUT33), .ZN(new_n265));
  XOR2_X1   g064(.A(G15gat), .B(G43gat), .Z(new_n266));
  XNOR2_X1  g065(.A(G71gat), .B(G99gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT32), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n254), .ZN(new_n271));
  AOI221_X4 g070(.A(new_n270), .B1(KEYINPUT33), .B2(new_n268), .C1(new_n271), .C2(new_n257), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n261), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n269), .A2(new_n261), .A3(new_n273), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n268), .B1(new_n262), .B2(KEYINPUT33), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n262), .A2(new_n270), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n260), .B1(new_n279), .B2(new_n272), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n276), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT36), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(new_n276), .ZN(new_n286));
  OAI21_X1  g085(.A(KEYINPUT36), .B1(new_n286), .B2(new_n274), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(G78gat), .B(G106gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(G22gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(G197gat), .ZN(new_n292));
  INV_X1    g091(.A(G204gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G211gat), .ZN(new_n295));
  INV_X1    g094(.A(G218gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n294), .B1(KEYINPUT22), .B2(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(G211gat), .B(G218gat), .Z(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(G141gat), .B(G148gat), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT2), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n302), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n304), .A2(new_n305), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n309));
  AOI22_X1  g108(.A1(new_n309), .A2(new_n303), .B1(G155gat), .B2(G162gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n308), .ZN(new_n312));
  OAI211_X1 g111(.A(new_n312), .B(new_n302), .C1(new_n303), .C2(new_n306), .ZN(new_n313));
  AND2_X1   g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT79), .B(KEYINPUT3), .Z(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n313), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n317), .A3(new_n320), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(G228gat), .A3(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n315), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n320), .A2(new_n325), .B1(G228gat), .B2(G233gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n319), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT31), .B(G50gat), .Z(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n329), .B1(new_n324), .B2(new_n327), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n291), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n332), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n334), .A2(new_n290), .A3(new_n330), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT29), .B1(new_n214), .B2(new_n223), .ZN(new_n338));
  NAND2_X1  g137(.A1(G226gat), .A2(G233gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT73), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n227), .A2(KEYINPUT74), .A3(new_n340), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT74), .B1(new_n227), .B2(new_n340), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n342), .B(new_n300), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n340), .B1(new_n227), .B2(new_n317), .ZN(new_n347));
  INV_X1    g146(.A(new_n340), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n214), .B2(new_n223), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n301), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(KEYINPUT75), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n345), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n341), .B1(new_n352), .B2(new_n343), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n300), .ZN(new_n355));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT76), .ZN(new_n357));
  XNOR2_X1  g156(.A(G64gat), .B(G92gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n351), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n360), .B1(new_n351), .B2(new_n355), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(KEYINPUT30), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n351), .A2(new_n355), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n359), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT77), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT77), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n363), .A2(new_n369), .A3(KEYINPUT30), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n364), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(G225gat), .A2(G233gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n372), .B(KEYINPUT81), .Z(new_n373));
  NOR2_X1   g172(.A1(new_n239), .A2(new_n244), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n316), .A2(new_n374), .A3(new_n321), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n316), .A2(KEYINPUT80), .A3(new_n374), .A4(new_n321), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n380));
  NAND3_X1  g179(.A1(new_n253), .A2(new_n314), .A3(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n314), .B1(new_n244), .B2(new_n239), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT5), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT88), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n379), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n379), .B2(new_n384), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n374), .A2(new_n320), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n382), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n373), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(KEYINPUT85), .A3(new_n373), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT5), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT86), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n245), .A2(new_n250), .A3(new_n314), .ZN(new_n398));
  INV_X1    g197(.A(new_n380), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n398), .A2(KEYINPUT83), .A3(new_n399), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n402), .B(new_n403), .C1(KEYINPUT4), .C2(new_n382), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT84), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n379), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n393), .A2(KEYINPUT86), .A3(KEYINPUT5), .A4(new_n394), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n404), .B2(new_n379), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n388), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G1gat), .B(G29gat), .Z(new_n411));
  XNOR2_X1  g210(.A(G57gat), .B(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n377), .A2(new_n378), .B1(new_n381), .B2(new_n383), .ZN(new_n418));
  INV_X1    g217(.A(new_n373), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT39), .B1(new_n390), .B2(new_n373), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OR3_X1    g221(.A1(new_n418), .A2(KEYINPUT39), .A3(new_n419), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n415), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT40), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n422), .A2(KEYINPUT40), .A3(new_n415), .A4(new_n423), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n417), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n337), .B1(new_n371), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT37), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n359), .B1(new_n365), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n431), .B1(new_n430), .B2(new_n365), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(KEYINPUT38), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT89), .B1(new_n353), .B2(new_n300), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n342), .B1(new_n344), .B2(new_n345), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n301), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n347), .A2(new_n349), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n434), .B(new_n437), .C1(new_n301), .C2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT38), .B1(new_n439), .B2(KEYINPUT37), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n363), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n410), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT6), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n415), .B(new_n388), .C1(new_n408), .C2(new_n409), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n417), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n433), .A2(new_n441), .A3(new_n442), .A4(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n288), .B1(new_n429), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n361), .B1(new_n366), .B2(new_n367), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n369), .B1(new_n363), .B2(KEYINPUT30), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n366), .A2(KEYINPUT77), .A3(new_n367), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n445), .A2(new_n442), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n337), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n336), .A2(new_n280), .A3(new_n276), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n451), .A2(new_n452), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT35), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT35), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n336), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n459), .B1(new_n445), .B2(new_n442), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n283), .A2(KEYINPUT90), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT90), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n275), .A2(new_n282), .A3(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n460), .A2(new_n451), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n447), .A2(new_n454), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT94), .ZN(new_n466));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467));
  INV_X1    g266(.A(G1gat), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(KEYINPUT16), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n467), .A2(new_n468), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n466), .B(G8gat), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT95), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n467), .A2(new_n468), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n467), .A2(KEYINPUT16), .A3(new_n468), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n466), .A2(G8gat), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n466), .A2(G8gat), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n471), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n472), .B1(new_n471), .B2(new_n477), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(G29gat), .A2(G36gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(KEYINPUT14), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT92), .B(G29gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n482), .B1(G36gat), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n485), .B(new_n488), .C1(KEYINPUT93), .C2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n481), .B(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G36gat), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n488), .B(new_n492), .C1(new_n493), .C2(new_n483), .ZN(new_n494));
  INV_X1    g293(.A(new_n489), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n492), .B(KEYINPUT93), .C1(new_n493), .C2(new_n483), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n490), .A2(KEYINPUT17), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT17), .B1(new_n490), .B2(new_n497), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n480), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(G229gat), .A2(G233gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT96), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n490), .A2(new_n497), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n471), .A2(new_n477), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n500), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT97), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n507), .A2(KEYINPUT18), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n503), .B(new_n504), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n502), .B(KEYINPUT13), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n508), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n500), .A2(new_n502), .A3(new_n505), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G197gat), .ZN(new_n518));
  XOR2_X1   g317(.A(KEYINPUT11), .B(G169gat), .Z(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n520), .B(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n516), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n509), .A2(new_n522), .A3(new_n513), .A4(new_n515), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n465), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G57gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(G64gat), .ZN(new_n530));
  INV_X1    g329(.A(G64gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G57gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G71gat), .A2(G78gat), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n537), .A2(KEYINPUT98), .ZN(new_n538));
  NOR2_X1   g337(.A1(G71gat), .A2(G78gat), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n539), .B1(KEYINPUT98), .B2(new_n537), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542));
  AND4_X1   g341(.A1(KEYINPUT99), .A2(new_n533), .A3(new_n542), .A4(new_n535), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n534), .B1(new_n530), .B2(new_n532), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT99), .B1(new_n544), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n541), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT101), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n542), .A3(new_n535), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n544), .A2(KEYINPUT99), .A3(new_n542), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n553), .A2(KEYINPUT101), .A3(new_n541), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n548), .A2(KEYINPUT21), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n504), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT102), .Z(new_n557));
  AOI21_X1  g356(.A(KEYINPUT21), .B1(new_n553), .B2(new_n541), .ZN(new_n558));
  AND2_X1   g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(new_n233), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n557), .A2(new_n561), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT100), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(G155gat), .ZN(new_n567));
  XOR2_X1   g366(.A(G183gat), .B(G211gat), .Z(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n562), .A2(new_n563), .A3(new_n569), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G99gat), .B(G106gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G99gat), .A2(G106gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT104), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT8), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT104), .B1(G99gat), .B2(G106gat), .ZN(new_n580));
  NOR3_X1   g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT103), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(KEYINPUT103), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n575), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n579), .B1(new_n576), .B2(new_n577), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n588), .B1(new_n577), .B2(new_n576), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n589), .A2(new_n574), .A3(new_n584), .A4(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(KEYINPUT105), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n498), .B2(new_n499), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n490), .A2(new_n497), .A3(new_n590), .A4(new_n587), .ZN(new_n594));
  NAND3_X1  g393(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n594), .A2(KEYINPUT106), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(KEYINPUT106), .B1(new_n594), .B2(new_n595), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(G190gat), .B(G218gat), .Z(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n599), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n604), .B(new_n593), .C1(new_n596), .C2(new_n597), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n603), .B1(new_n600), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n573), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n587), .A2(new_n590), .A3(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n548), .A2(new_n554), .A3(new_n612), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n613), .A2(KEYINPUT107), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT107), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n548), .A2(new_n554), .A3(new_n615), .A4(new_n612), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n546), .A2(new_n591), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n553), .A2(new_n541), .A3(new_n590), .A4(new_n587), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n611), .B1(new_n614), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n617), .A2(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(new_n611), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  NAND3_X1  g427(.A1(new_n622), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n628), .B1(new_n622), .B2(new_n625), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n610), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n452), .B(KEYINPUT108), .Z(new_n635));
  NAND3_X1  g434(.A1(new_n528), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT109), .B(G1gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(G1324gat));
  NAND3_X1  g437(.A1(new_n528), .A2(new_n371), .A3(new_n634), .ZN(new_n639));
  XNOR2_X1  g438(.A(KEYINPUT16), .B(G8gat), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT110), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT42), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(KEYINPUT110), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(G8gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(G1325gat));
  INV_X1    g446(.A(G15gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n461), .A2(new_n463), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n528), .A2(new_n648), .A3(new_n650), .A4(new_n634), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n528), .A2(new_n634), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n652), .A2(new_n288), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n651), .B1(new_n653), .B2(new_n648), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n337), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(G1327gat));
  NOR3_X1   g456(.A1(new_n573), .A2(new_n609), .A3(new_n633), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n528), .A2(new_n483), .A3(new_n635), .A4(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(KEYINPUT111), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(KEYINPUT111), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT45), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n465), .B2(new_n609), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n429), .A2(new_n446), .ZN(new_n667));
  INV_X1    g466(.A(new_n288), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n454), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n457), .A2(new_n464), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n671), .A2(KEYINPUT44), .A3(new_n608), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n573), .A2(new_n527), .A3(new_n633), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n673), .A2(new_n635), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n484), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n660), .A2(KEYINPUT45), .A3(new_n661), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n664), .A2(new_n676), .A3(new_n677), .ZN(G1328gat));
  NOR2_X1   g477(.A1(new_n451), .A2(G36gat), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n671), .A2(new_n526), .A3(new_n658), .A4(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT46), .Z(new_n681));
  NAND4_X1  g480(.A1(new_n666), .A2(new_n672), .A3(new_n371), .A4(new_n674), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(G36gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT112), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT112), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n681), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(G1329gat));
  AND2_X1   g487(.A1(new_n528), .A2(new_n658), .ZN(new_n689));
  INV_X1    g488(.A(G43gat), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n690), .A3(new_n650), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n666), .A2(new_n672), .A3(new_n288), .A4(new_n674), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G43gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1330gat));
  INV_X1    g495(.A(G50gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n689), .A2(new_n697), .A3(new_n337), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n666), .A2(new_n672), .A3(new_n337), .A4(new_n674), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G50gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT48), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1331gat));
  NAND3_X1  g502(.A1(new_n573), .A2(new_n609), .A3(new_n633), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n465), .A2(new_n526), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n635), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g506(.A(new_n451), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT113), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n705), .A2(new_n711), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1333gat));
  INV_X1    g514(.A(G71gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n705), .A2(new_n716), .A3(new_n650), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n705), .A2(new_n288), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n717), .B1(new_n718), .B2(new_n716), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1334gat));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n337), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g522(.A1(new_n573), .A2(new_n526), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n632), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n673), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n635), .ZN(new_n728));
  OAI21_X1  g527(.A(G85gat), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n671), .A2(new_n608), .A3(new_n724), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT51), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n609), .B1(new_n669), .B2(new_n670), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n724), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n728), .A2(G85gat), .A3(new_n632), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT114), .Z(new_n738));
  OAI21_X1  g537(.A(new_n729), .B1(new_n736), .B2(new_n738), .ZN(G1336gat));
  NOR2_X1   g538(.A1(new_n451), .A2(new_n632), .ZN(new_n740));
  AOI21_X1  g539(.A(G92gat), .B1(new_n735), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(KEYINPUT115), .ZN(new_n743));
  INV_X1    g542(.A(G92gat), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n451), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n666), .A2(new_n672), .A3(new_n726), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n742), .A2(KEYINPUT115), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n741), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n743), .ZN(new_n750));
  NOR4_X1   g549(.A1(new_n465), .A2(new_n731), .A3(new_n609), .A4(new_n725), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT51), .B1(new_n733), .B2(new_n724), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n740), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n744), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n746), .A2(new_n747), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n749), .A2(new_n756), .ZN(G1337gat));
  OAI21_X1  g556(.A(G99gat), .B1(new_n727), .B2(new_n668), .ZN(new_n758));
  OR3_X1    g557(.A1(new_n649), .A2(G99gat), .A3(new_n632), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n736), .B2(new_n759), .ZN(G1338gat));
  NOR3_X1   g559(.A1(new_n336), .A2(G106gat), .A3(new_n632), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n735), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n666), .A2(new_n672), .A3(new_n337), .A4(new_n726), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G106gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n762), .A2(KEYINPUT116), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT53), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n762), .B(new_n764), .C1(KEYINPUT116), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1339gat));
  NAND4_X1  g569(.A1(new_n573), .A2(new_n527), .A3(new_n609), .A4(new_n632), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n613), .A2(KEYINPUT107), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n624), .A3(new_n620), .A4(new_n616), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n622), .A2(KEYINPUT54), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n776), .B(new_n611), .C1(new_n614), .C2(new_n621), .ZN(new_n777));
  INV_X1    g576(.A(new_n628), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n777), .A2(KEYINPUT117), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT117), .B1(new_n777), .B2(new_n778), .ZN(new_n780));
  OAI211_X1 g579(.A(KEYINPUT55), .B(new_n775), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n629), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n775), .B1(new_n779), .B2(new_n780), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n510), .A2(new_n512), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n502), .B1(new_n500), .B2(new_n505), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n520), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n525), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n782), .A2(new_n608), .A3(new_n785), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n632), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n783), .A2(new_n784), .B1(new_n524), .B2(new_n525), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n782), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n609), .B1(new_n794), .B2(KEYINPUT118), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n785), .A2(new_n526), .A3(new_n629), .A4(new_n781), .ZN(new_n796));
  INV_X1    g595(.A(new_n792), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n796), .A2(KEYINPUT118), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n791), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n573), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n772), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n337), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n803), .A2(new_n451), .A3(new_n650), .A4(new_n635), .ZN(new_n804));
  OAI21_X1  g603(.A(G113gat), .B1(new_n804), .B2(new_n527), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n803), .A2(new_n635), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n451), .A2(new_n280), .A3(new_n276), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n527), .A2(G113gat), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT119), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n805), .B1(new_n809), .B2(new_n811), .ZN(G1340gat));
  INV_X1    g611(.A(G120gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n804), .A2(new_n813), .A3(new_n632), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n808), .A2(new_n633), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n814), .B1(new_n813), .B2(new_n815), .ZN(G1341gat));
  OAI21_X1  g615(.A(new_n233), .B1(new_n809), .B2(new_n801), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n233), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OR3_X1    g618(.A1(new_n804), .A2(KEYINPUT120), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT120), .B1(new_n804), .B2(new_n819), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n817), .A2(new_n820), .A3(new_n821), .ZN(G1342gat));
  NAND2_X1  g621(.A1(new_n608), .A2(new_n231), .ZN(new_n823));
  OR3_X1    g622(.A1(new_n809), .A2(KEYINPUT56), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G134gat), .B1(new_n804), .B2(new_n609), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT56), .B1(new_n809), .B2(new_n823), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(G1343gat));
  AOI21_X1  g626(.A(new_n608), .B1(new_n796), .B2(new_n797), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n785), .A2(new_n608), .A3(new_n790), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n781), .A2(new_n629), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n801), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n771), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n336), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT121), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n834), .B1(new_n802), .B2(new_n336), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n728), .A2(new_n371), .A3(new_n288), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n526), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(G141gat), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n802), .A2(new_n336), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n840), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(G141gat), .A3(new_n527), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(G141gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n841), .B2(new_n526), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT58), .B1(new_n851), .B2(new_n847), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n849), .A2(new_n852), .ZN(G1344gat));
  OAI21_X1  g652(.A(KEYINPUT59), .B1(new_n846), .B2(new_n632), .ZN(new_n854));
  INV_X1    g653(.A(G148gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n633), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(KEYINPUT59), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n854), .A2(new_n855), .B1(new_n857), .B2(new_n839), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n336), .B1(new_n832), .B2(new_n771), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(KEYINPUT57), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n791), .B1(new_n794), .B2(new_n608), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n772), .B1(new_n862), .B2(new_n801), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT123), .B(new_n834), .C1(new_n863), .C2(new_n336), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n835), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n802), .B2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n796), .A2(new_n797), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n609), .A3(new_n798), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n573), .B1(new_n872), .B2(new_n791), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n868), .B(new_n835), .C1(new_n873), .C2(new_n772), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n865), .A2(new_n867), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n875), .A2(new_n633), .A3(new_n840), .ZN(new_n876));
  NAND2_X1  g675(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n858), .B1(new_n876), .B2(new_n877), .ZN(G1345gat));
  AOI21_X1  g677(.A(new_n304), .B1(new_n841), .B2(new_n573), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n846), .A2(G155gat), .A3(new_n801), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n879), .A2(new_n880), .ZN(G1346gat));
  AOI21_X1  g680(.A(new_n305), .B1(new_n841), .B2(new_n608), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n846), .A2(G162gat), .A3(new_n609), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n882), .A2(new_n883), .ZN(G1347gat));
  NOR3_X1   g683(.A1(new_n635), .A2(new_n451), .A3(new_n649), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n803), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(KEYINPUT124), .A3(new_n803), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(G169gat), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n527), .ZN(new_n892));
  INV_X1    g691(.A(new_n802), .ZN(new_n893));
  AND4_X1   g692(.A1(new_n371), .A2(new_n893), .A3(new_n455), .A4(new_n728), .ZN(new_n894));
  AOI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n526), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n892), .A2(new_n895), .ZN(G1348gat));
  OAI21_X1  g695(.A(G176gat), .B1(new_n890), .B2(new_n632), .ZN(new_n897));
  INV_X1    g696(.A(G176gat), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n894), .A2(new_n898), .A3(new_n633), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1349gat));
  OAI21_X1  g699(.A(G183gat), .B1(new_n890), .B2(new_n801), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n215), .A3(new_n573), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT60), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT60), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n894), .A2(new_n216), .A3(new_n608), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n608), .A3(new_n889), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n910));
  AND3_X1   g709(.A1(new_n909), .A2(new_n910), .A3(G190gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n909), .B2(G190gat), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n635), .A2(new_n451), .A3(new_n288), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n845), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(G197gat), .A3(new_n527), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n916), .B(KEYINPUT125), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n875), .A2(new_n526), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G197gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1352gat));
  INV_X1    g719(.A(new_n915), .ZN(new_n921));
  AOI21_X1  g720(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n633), .A3(new_n922), .ZN(new_n923));
  NOR2_X1   g722(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AND3_X1   g724(.A1(new_n875), .A2(new_n633), .A3(new_n914), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n293), .B2(new_n926), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n921), .A2(new_n295), .A3(new_n573), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT127), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n875), .A2(new_n914), .A3(new_n929), .A4(new_n573), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n930), .A2(G211gat), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n875), .A2(new_n573), .A3(new_n914), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT127), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  AND4_X1   g733(.A1(KEYINPUT63), .A2(new_n933), .A3(G211gat), .A4(new_n930), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n928), .B1(new_n934), .B2(new_n935), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n921), .A2(new_n296), .A3(new_n608), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n875), .A2(new_n608), .A3(new_n914), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n296), .ZN(G1355gat));
endmodule


