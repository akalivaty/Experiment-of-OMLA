//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:29 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g043(.A1(new_n468), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n468), .A2(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n467), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n477), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(new_n480), .A2(G138), .ZN(new_n486));
  XOR2_X1   g061(.A(KEYINPUT69), .B(KEYINPUT4), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n480), .B(G138), .C1(KEYINPUT69), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n477), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n463), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G102), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G50), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT70), .A2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT70), .A2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT5), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n507), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT70), .B(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT71), .B1(new_n514), .B2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g090(.A(new_n504), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(new_n502), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n513), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n506), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n513), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G62), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  XOR2_X1   g100(.A(new_n525), .B(KEYINPUT72), .Z(new_n526));
  AOI21_X1  g101(.A(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(G166));
  NAND2_X1  g103(.A1(new_n518), .A2(G89), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n531), .B(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n505), .A2(G51), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n529), .A2(new_n530), .A3(new_n532), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AND2_X1   g110(.A1(new_n523), .A2(G64), .ZN(new_n536));
  AND2_X1   g111(.A1(G77), .A2(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(G651), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n505), .A2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n518), .A2(G90), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n501), .ZN(new_n545));
  NAND2_X1  g120(.A1(KEYINPUT70), .A2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g122(.A(KEYINPUT71), .B1(new_n547), .B2(new_n511), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n510), .A2(new_n507), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n548), .A2(G56), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(G68), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n517), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n548), .A2(G81), .A3(new_n553), .A4(new_n549), .ZN(new_n554));
  XNOR2_X1  g129(.A(KEYINPUT73), .B(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n505), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n554), .A2(KEYINPUT74), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(KEYINPUT74), .B1(new_n554), .B2(new_n556), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n562), .A2(new_n565), .ZN(G188));
  NAND3_X1  g141(.A1(new_n548), .A2(G65), .A3(new_n549), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G651), .B1(G91), .B2(new_n518), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT76), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n572));
  NOR2_X1   g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n505), .B2(G53), .ZN(new_n574));
  OAI211_X1 g149(.A(G53), .B(G543), .C1(new_n516), .C2(new_n502), .ZN(new_n575));
  XNOR2_X1  g150(.A(KEYINPUT75), .B(KEYINPUT9), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n571), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n575), .B1(new_n572), .B2(KEYINPUT9), .ZN(new_n579));
  INV_X1    g154(.A(new_n576), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n505), .A2(new_n580), .A3(G53), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n579), .A2(new_n581), .A3(KEYINPUT76), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g158(.A(KEYINPUT77), .B1(new_n570), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n513), .A2(new_n515), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n568), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n518), .A2(G91), .ZN(new_n589));
  AND4_X1   g164(.A1(KEYINPUT77), .A2(new_n588), .A3(new_n589), .A4(new_n583), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n584), .A2(new_n590), .ZN(G299));
  INV_X1    g166(.A(G166), .ZN(G303));
  NAND2_X1  g167(.A1(new_n518), .A2(G87), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT78), .Z(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n505), .A2(G49), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(new_n518), .A2(G86), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n523), .A2(G61), .ZN(new_n601));
  INV_X1    g176(.A(G73), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n501), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G48), .B2(new_n505), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(G305));
  AOI22_X1  g180(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n606), .A2(new_n522), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n505), .A2(G47), .ZN(new_n608));
  INV_X1    g183(.A(G85), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n519), .B2(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(G290));
  NAND2_X1  g187(.A1(G301), .A2(G868), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n548), .A2(G92), .A3(new_n553), .A4(new_n549), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n505), .A2(G54), .ZN(new_n619));
  AND3_X1   g194(.A1(new_n548), .A2(G66), .A3(new_n549), .ZN(new_n620));
  AND2_X1   g195(.A1(G79), .A2(G543), .ZN(new_n621));
  OAI21_X1  g196(.A(G651), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(KEYINPUT80), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT80), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n613), .B1(new_n629), .B2(G868), .ZN(G284));
  OAI21_X1  g205(.A(new_n613), .B1(new_n629), .B2(G868), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  INV_X1    g207(.A(G299), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G297));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n629), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(G868), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n641));
  XNOR2_X1  g216(.A(G323), .B(new_n641), .ZN(G282));
  NAND2_X1  g217(.A1(new_n468), .A2(new_n495), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2100), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n478), .A2(G123), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n480), .A2(G135), .ZN(new_n649));
  NOR2_X1   g224(.A1(G99), .A2(G2105), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(new_n477), .B2(G111), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n653), .ZN(G156));
  XOR2_X1   g229(.A(KEYINPUT15), .B(G2435), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2438), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT14), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(KEYINPUT85), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n658), .A2(new_n659), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G1348), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2451), .B(G2454), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT84), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n664), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT86), .B(G1341), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G14), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n677), .A2(new_n678), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT17), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT18), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n684), .B(new_n685), .C1(new_n683), .C2(new_n679), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n685), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(G2096), .B(G2100), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XOR2_X1   g264(.A(G1971), .B(G1976), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1956), .B(G2474), .Z(new_n693));
  XOR2_X1   g268(.A(G1961), .B(G1966), .Z(new_n694));
  AND2_X1   g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT88), .Z(new_n697));
  OR2_X1    g272(.A1(new_n697), .A2(KEYINPUT20), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(KEYINPUT20), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n693), .A2(new_n694), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n692), .A2(new_n700), .ZN(new_n701));
  OR3_X1    g276(.A1(new_n692), .A2(new_n700), .A3(new_n695), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1986), .B(G1996), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1981), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1991), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n705), .B(new_n708), .ZN(G229));
  AND2_X1   g284(.A1(KEYINPUT89), .A2(G16), .ZN(new_n710));
  NOR2_X1   g285(.A1(KEYINPUT89), .A2(G16), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G24), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n611), .B(KEYINPUT91), .Z(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n713), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT92), .B(G1986), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n478), .A2(G119), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G131), .ZN(new_n724));
  OR2_X1    g299(.A1(G95), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G107), .C2(new_n477), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n722), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT35), .B(G1991), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n719), .A2(new_n720), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n713), .A2(G22), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G166), .B2(new_n713), .ZN(new_n734));
  MUX2_X1   g309(.A(new_n733), .B(new_n734), .S(KEYINPUT94), .Z(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1971), .Z(new_n736));
  INV_X1    g311(.A(G16), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G6), .ZN(new_n738));
  INV_X1    g313(.A(G305), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n738), .B1(new_n739), .B2(new_n737), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT32), .B(G1981), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n737), .A2(G23), .ZN(new_n743));
  INV_X1    g318(.A(G288), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n737), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT33), .B(G1976), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT93), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n736), .A2(new_n742), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n732), .B1(new_n749), .B2(KEYINPUT34), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n750), .B1(KEYINPUT34), .B2(new_n749), .C1(new_n730), .C2(new_n729), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT36), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n713), .A2(G19), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n560), .B2(new_n713), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT95), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(G1341), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n713), .A2(KEYINPUT23), .A3(G20), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G20), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n712), .B2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n757), .B(new_n760), .C1(new_n633), .C2(new_n737), .ZN(new_n761));
  INV_X1    g336(.A(G1956), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT31), .B(G11), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT102), .B(G28), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT30), .ZN(new_n766));
  MUX2_X1   g341(.A(new_n766), .B(new_n652), .S(G29), .Z(new_n767));
  NAND2_X1  g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(KEYINPUT24), .A2(G34), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n769), .A2(new_n770), .A3(G29), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n475), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n764), .B(new_n767), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n480), .A2(G139), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT99), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  OR3_X1    g352(.A1(new_n777), .A2(KEYINPUT100), .A3(new_n477), .ZN(new_n778));
  OAI21_X1  g353(.A(KEYINPUT100), .B1(new_n777), .B2(new_n477), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT98), .B(KEYINPUT25), .Z(new_n780));
  NAND2_X1  g355(.A1(new_n495), .A2(G103), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND4_X1  g357(.A1(new_n776), .A2(new_n778), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G33), .B(new_n783), .S(G29), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2072), .ZN(new_n785));
  AOI211_X1 g360(.A(new_n774), .B(new_n785), .C1(new_n773), .C2(new_n772), .ZN(new_n786));
  AOI22_X1  g361(.A1(G129), .A2(new_n478), .B1(new_n480), .B2(G141), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n495), .A2(G105), .ZN(new_n788));
  NAND3_X1  g363(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT26), .Z(new_n790));
  NAND3_X1  g365(.A1(new_n787), .A2(new_n788), .A3(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G32), .B(new_n791), .S(G29), .Z(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT27), .B(G1996), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n721), .A2(G26), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n480), .A2(G140), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT96), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n478), .A2(G128), .ZN(new_n798));
  NOR2_X1   g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI21_X1  g374(.A(G2104), .B1(new_n477), .B2(G116), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(G29), .ZN(new_n802));
  MUX2_X1   g377(.A(new_n795), .B(new_n802), .S(KEYINPUT28), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT97), .B(G2067), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n786), .A2(new_n794), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n721), .A2(G35), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G162), .B2(new_n721), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT29), .Z(new_n809));
  INV_X1    g384(.A(G2090), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT104), .Z(new_n812));
  NAND2_X1  g387(.A1(new_n721), .A2(G27), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G164), .B2(new_n721), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(G2078), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n737), .A2(G5), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G171), .B2(new_n737), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT103), .B(G1961), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G16), .A2(G21), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G168), .B2(G16), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(G1966), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G2078), .B2(new_n814), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n819), .B(new_n823), .C1(new_n810), .C2(new_n809), .ZN(new_n824));
  NOR4_X1   g399(.A1(new_n806), .A2(new_n812), .A3(new_n815), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n821), .A2(G1966), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT101), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n737), .A2(G4), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n629), .B2(new_n737), .ZN(new_n829));
  INV_X1    g404(.A(G1348), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  AND4_X1   g406(.A1(new_n763), .A2(new_n825), .A3(new_n827), .A4(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n752), .A2(new_n756), .A3(new_n832), .ZN(G150));
  INV_X1    g408(.A(G150), .ZN(G311));
  NOR2_X1   g409(.A1(new_n628), .A2(new_n636), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT105), .B(KEYINPUT38), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n548), .A2(G67), .A3(new_n549), .ZN(new_n839));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n522), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g416(.A1(new_n548), .A2(G93), .A3(new_n553), .A4(new_n549), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n505), .A2(G55), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n559), .A2(new_n845), .ZN(new_n846));
  OAI221_X1 g421(.A(new_n552), .B1(new_n841), .B2(new_n844), .C1(new_n557), .C2(new_n558), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n838), .B(new_n848), .Z(new_n849));
  NOR2_X1   g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT106), .Z(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n513), .A2(new_n515), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n840), .ZN(new_n854));
  OAI21_X1  g429(.A(G651), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(new_n843), .A3(new_n842), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G860), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT107), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n851), .A2(new_n859), .ZN(G145));
  AND2_X1   g435(.A1(new_n492), .A2(new_n493), .ZN(new_n861));
  OAI211_X1 g436(.A(KEYINPUT108), .B(new_n496), .C1(new_n861), .C2(new_n477), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT108), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n494), .B2(new_n497), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n862), .A2(new_n864), .B1(new_n488), .B2(new_n490), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n801), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n791), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n783), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n478), .A2(G130), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n480), .A2(G142), .ZN(new_n871));
  NOR2_X1   g446(.A1(G106), .A2(G2105), .ZN(new_n872));
  OAI21_X1  g447(.A(G2104), .B1(new_n477), .B2(G118), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n870), .B(new_n871), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n644), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n727), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n475), .B(new_n652), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n484), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n869), .A2(KEYINPUT109), .A3(new_n876), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n877), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n882), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g463(.A(new_n638), .B(new_n848), .Z(new_n889));
  OAI21_X1  g464(.A(new_n623), .B1(new_n584), .B2(new_n590), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n588), .A2(new_n583), .A3(new_n589), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT77), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n570), .A2(KEYINPUT77), .A3(new_n583), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n625), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n890), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n890), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n890), .A2(new_n895), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n900), .B1(new_n901), .B2(new_n889), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(G290), .A2(new_n604), .A3(new_n600), .ZN(new_n905));
  NAND2_X1  g480(.A1(G305), .A2(new_n611), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(G288), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(G288), .B1(new_n905), .B2(new_n906), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT110), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n911));
  NAND2_X1  g486(.A1(G166), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT111), .B1(new_n521), .B2(new_n527), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n910), .A3(new_n913), .ZN(new_n915));
  OAI22_X1  g490(.A1(new_n908), .A2(new_n909), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n909), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n907), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n902), .A2(new_n903), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n904), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n920), .B1(new_n904), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G868), .B2(new_n845), .ZN(G295));
  OAI21_X1  g500(.A(new_n924), .B1(G868), .B2(new_n845), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n846), .A2(G301), .A3(new_n847), .ZN(new_n928));
  AOI21_X1  g503(.A(G301), .B1(new_n846), .B2(new_n847), .ZN(new_n929));
  OAI21_X1  g504(.A(G286), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n559), .A2(new_n845), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n554), .A2(new_n556), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT74), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n554), .A2(KEYINPUT74), .A3(new_n556), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n856), .B1(new_n936), .B2(new_n552), .ZN(new_n937));
  OAI21_X1  g512(.A(G171), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n846), .A2(new_n847), .A3(G301), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(G168), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(new_n940), .A3(new_n901), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT114), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT114), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n930), .A2(new_n940), .A3(new_n943), .A4(new_n901), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n930), .A2(new_n940), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n898), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n916), .A2(new_n919), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n945), .A2(new_n898), .A3(KEYINPUT112), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n951), .A2(new_n920), .A3(new_n941), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(G37), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n949), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT115), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT115), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n949), .A2(new_n953), .A3(new_n957), .A4(new_n954), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n927), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n951), .A2(new_n941), .A3(new_n952), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n916), .A2(new_n919), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n962), .A2(new_n951), .A3(new_n941), .A4(new_n952), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n954), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n966), .A2(new_n927), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n959), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT116), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n949), .A2(new_n953), .A3(new_n927), .A4(new_n954), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n968), .A2(new_n969), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n969), .B1(new_n968), .B2(new_n974), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(G397));
  NOR2_X1   g552(.A1(new_n865), .A2(G1384), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n470), .A2(G40), .A3(new_n474), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n801), .B(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n791), .B(G1996), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n727), .A2(new_n730), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT126), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g565(.A1(new_n801), .A2(G2067), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n982), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n982), .A2(G1996), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT46), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n993), .B(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n982), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n985), .B2(new_n791), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n996), .B(new_n998), .C1(new_n994), .C2(KEYINPUT46), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(KEYINPUT47), .Z(new_n1000));
  INV_X1    g575(.A(new_n730), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n987), .B1(new_n1001), .B2(new_n728), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n997), .B1(new_n1002), .B2(new_n988), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n982), .A2(G290), .A3(G1986), .ZN(new_n1004));
  XOR2_X1   g579(.A(new_n1004), .B(KEYINPUT48), .Z(new_n1005));
  AOI211_X1 g580(.A(new_n992), .B(new_n1000), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1981), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n739), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n604), .A2(new_n598), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(G1981), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT49), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n978), .A2(new_n981), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT117), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT117), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1976), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1015), .B1(G288), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT52), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n744), .A2(G1976), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1024), .A2(new_n1022), .A3(KEYINPUT52), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n499), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n980), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1026), .A2(new_n981), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1031), .A2(G1971), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n978), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n981), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G2090), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1014), .B1(new_n1032), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(G166), .A2(new_n1014), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT55), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .A4(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n980), .B1(new_n865), .B2(G1384), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n981), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT118), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n1027), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1044), .A2(new_n1048), .A3(new_n981), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1966), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1036), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1050), .A2(new_n1051), .B1(new_n1052), .B2(new_n773), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(new_n1014), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G168), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT63), .B1(new_n1043), .B2(new_n1055), .ZN(new_n1056));
  AOI211_X1 g631(.A(G1976), .B(G288), .C1(new_n1018), .C2(new_n1019), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1008), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1015), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n499), .A2(new_n1033), .A3(new_n1027), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n981), .B(new_n1061), .C1(new_n978), .C2(new_n1033), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1032), .B1(G2090), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1041), .B1(new_n1063), .B2(G8), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1064), .A2(KEYINPUT63), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1060), .B1(new_n1065), .B2(new_n1055), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1066), .A2(new_n1020), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1056), .A2(new_n1059), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1020), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(G8), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1054), .A2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1071), .B(KEYINPUT121), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1052), .A2(new_n773), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1076), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT122), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1075), .B1(new_n1053), .B2(new_n1014), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT51), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1074), .B1(new_n1081), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1053), .A2(new_n1071), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1070), .B(KEYINPUT62), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1084), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1083), .B1(new_n1082), .B2(KEYINPUT51), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1088), .A2(new_n1089), .B1(new_n1054), .B2(new_n1073), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1086), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G2078), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1046), .A2(new_n1094), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT123), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT53), .B1(new_n1095), .B2(KEYINPUT123), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n1031), .B2(new_n1094), .ZN(new_n1099));
  INV_X1    g674(.A(G1961), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1099), .B1(new_n1100), .B2(new_n1036), .ZN(new_n1101));
  AOI21_X1  g676(.A(G301), .B1(new_n1098), .B2(new_n1101), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n1070), .A2(KEYINPUT62), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1087), .A2(new_n1093), .A3(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1045), .A2(KEYINPUT124), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1107), .B1(new_n1045), .B2(KEYINPUT124), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1106), .A2(new_n1108), .A3(new_n1094), .A4(new_n1026), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1101), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(G171), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1101), .B(G301), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1112), .A2(KEYINPUT54), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1062), .A2(new_n762), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT56), .B(G2072), .Z(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1026), .A2(new_n1029), .A3(new_n981), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n579), .B2(new_n581), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n570), .A2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1119), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1118), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1122), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1036), .A2(new_n830), .B1(new_n1013), .B2(new_n983), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n628), .A2(KEYINPUT60), .ZN(new_n1128));
  AOI22_X1  g703(.A1(new_n1126), .A2(KEYINPUT61), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT61), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT120), .B1(new_n1118), .B2(new_n1122), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1114), .A2(new_n1117), .A3(new_n1124), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1130), .B1(new_n1134), .B2(new_n1125), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1127), .A2(new_n628), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1127), .A2(new_n628), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT60), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(KEYINPUT58), .B(G1341), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n1030), .A2(G1996), .B1(new_n1013), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n560), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT59), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1129), .A2(new_n1135), .A3(new_n1138), .A4(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1131), .B(new_n1133), .C1(new_n1137), .C2(new_n1125), .ZN(new_n1144));
  AOI22_X1  g719(.A1(new_n1111), .A2(new_n1113), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1110), .A2(G171), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1147), .B1(new_n1102), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1069), .B1(new_n1105), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1064), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1068), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1002), .A2(new_n988), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n611), .B(G1986), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n982), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1006), .B1(new_n1153), .B2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g732(.A1(G229), .A2(new_n461), .ZN(new_n1159));
  NOR2_X1   g733(.A1(G401), .A2(G227), .ZN(new_n1160));
  NAND4_X1  g734(.A1(new_n887), .A2(new_n972), .A3(new_n1159), .A4(new_n1160), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


