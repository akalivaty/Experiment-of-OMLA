//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n806,
    new_n808, new_n809, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  INV_X1    g004(.A(G8gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT96), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n208), .A2(new_n209), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  OR3_X1    g012(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  OAI221_X1 g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT15), .C2(new_n208), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT98), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(KEYINPUT97), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n214), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n215), .A2(KEYINPUT97), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n223), .A2(new_n224), .B1(new_n217), .B2(new_n218), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n213), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n207), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n226), .ZN(new_n228));
  XNOR2_X1  g027(.A(new_n228), .B(KEYINPUT17), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n227), .B1(new_n229), .B2(new_n207), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  AND2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OR2_X1    g031(.A1(new_n232), .A2(KEYINPUT18), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(KEYINPUT18), .ZN(new_n234));
  XOR2_X1   g033(.A(new_n228), .B(new_n207), .Z(new_n235));
  XOR2_X1   g034(.A(new_n231), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n233), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G113gat), .B(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XOR2_X1   g039(.A(KEYINPUT11), .B(G169gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n242), .B(KEYINPUT12), .Z(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n243), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n233), .A2(new_n245), .A3(new_n234), .A4(new_n237), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G226gat), .ZN(new_n249));
  INV_X1    g048(.A(G233gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(KEYINPUT65), .B(G176gat), .ZN(new_n253));
  INV_X1    g052(.A(G169gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n253), .A2(KEYINPUT23), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G183gat), .ZN(new_n258));
  INV_X1    g057(.A(G190gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G183gat), .A2(G190gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(KEYINPUT24), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G169gat), .A2(G176gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(KEYINPUT23), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n261), .A2(KEYINPUT24), .ZN(new_n265));
  INV_X1    g064(.A(G176gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n253), .A2(KEYINPUT66), .A3(KEYINPUT23), .A4(new_n254), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n257), .A2(new_n262), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n271), .B1(new_n263), .B2(KEYINPUT23), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n262), .A3(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n263), .A2(KEYINPUT26), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(new_n267), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n263), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT27), .B(G183gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(KEYINPUT28), .A3(new_n259), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n258), .A2(KEYINPUT27), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT67), .ZN(new_n283));
  AOI21_X1  g082(.A(G190gat), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n258), .A2(KEYINPUT67), .A3(KEYINPUT27), .ZN(new_n285));
  XNOR2_X1  g084(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n284), .B(new_n285), .C1(new_n258), .C2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT69), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT27), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n283), .B1(new_n290), .B2(G183gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(new_n259), .A3(new_n285), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(KEYINPUT68), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT27), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n258), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(KEYINPUT69), .B(new_n288), .C1(new_n292), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n281), .B1(new_n289), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT70), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n279), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n281), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n288), .B1(new_n292), .B2(new_n296), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI211_X1 g104(.A(new_n300), .B(new_n302), .C1(new_n305), .C2(new_n297), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n275), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n252), .B1(new_n308), .B2(KEYINPUT29), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n310));
  OR2_X1    g109(.A1(new_n310), .A2(KEYINPUT80), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(KEYINPUT80), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G211gat), .B(G218gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n314), .B(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n272), .A2(new_n274), .ZN(new_n318));
  INV_X1    g117(.A(new_n279), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n302), .B1(new_n305), .B2(new_n297), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT70), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n318), .B1(new_n321), .B2(new_n306), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n323));
  AND3_X1   g122(.A1(new_n322), .A2(new_n323), .A3(new_n251), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n322), .B2(new_n251), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n309), .B(new_n317), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n308), .A2(new_n252), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n251), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n316), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n326), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n331), .A2(KEYINPUT37), .ZN(new_n332));
  XOR2_X1   g131(.A(G8gat), .B(G36gat), .Z(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(KEYINPUT82), .ZN(new_n334));
  XNOR2_X1  g133(.A(G64gat), .B(G92gat), .ZN(new_n335));
  XOR2_X1   g134(.A(new_n334), .B(new_n335), .Z(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n331), .B2(KEYINPUT37), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT38), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT38), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(new_n337), .C1(new_n331), .C2(KEYINPUT37), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT81), .B1(new_n308), .B2(new_n252), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n323), .A3(new_n251), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n329), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT94), .B1(new_n345), .B2(new_n317), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n309), .B1(new_n324), .B2(new_n325), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n316), .ZN(new_n349));
  OAI211_X1 g148(.A(new_n309), .B(new_n317), .C1(new_n252), .C2(new_n308), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT37), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G155gat), .ZN(new_n354));
  INV_X1    g153(.A(G162gat), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT84), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n357), .B1(G155gat), .B2(G162gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G141gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G148gat), .ZN(new_n362));
  INV_X1    g161(.A(G148gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(G141gat), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT2), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  OR2_X1    g164(.A1(new_n360), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(KEYINPUT85), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT85), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G148gat), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n367), .A2(new_n369), .A3(G141gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n362), .ZN(new_n371));
  OR2_X1    g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n359), .B1(new_n372), .B2(KEYINPUT2), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n366), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(G120gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G113gat), .ZN(new_n377));
  INV_X1    g176(.A(G113gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G120gat), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT1), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(G134gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT72), .B1(new_n381), .B2(G127gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT72), .ZN(new_n383));
  INV_X1    g182(.A(G127gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(G134gat), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT71), .B(G134gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G127gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n380), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT73), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n381), .A2(G127gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n384), .A2(G134gat), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT73), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n392), .A2(new_n395), .A3(new_n380), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n375), .B1(new_n389), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n386), .A2(new_n388), .ZN(new_n398));
  INV_X1    g197(.A(new_n380), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n392), .A2(new_n395), .A3(new_n380), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n374), .A3(new_n366), .A4(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n397), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n400), .A2(new_n401), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT86), .A3(new_n375), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT5), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n375), .A2(KEYINPUT3), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT3), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n366), .A2(new_n374), .A3(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n413), .A3(new_n407), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n402), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n396), .A2(new_n389), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n374), .A4(new_n366), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n414), .A2(new_n416), .A3(new_n418), .A4(new_n405), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT5), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND3_X1  g227(.A1(new_n420), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT93), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n420), .A2(new_n423), .ZN(new_n431));
  INV_X1    g230(.A(new_n428), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XOR2_X1   g232(.A(KEYINPUT88), .B(KEYINPUT6), .Z(new_n434));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n420), .A2(new_n423), .A3(new_n435), .A4(new_n428), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n430), .A2(new_n433), .A3(new_n434), .A4(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n429), .A2(new_n434), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n326), .A2(new_n330), .A3(new_n336), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT95), .B1(new_n353), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n443), .B(new_n440), .C1(new_n342), .C2(new_n352), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n339), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(G78gat), .B(G106gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT31), .B(G50gat), .ZN(new_n447));
  XOR2_X1   g246(.A(new_n446), .B(new_n447), .Z(new_n448));
  OAI21_X1  g247(.A(new_n412), .B1(new_n316), .B2(KEYINPUT29), .ZN(new_n449));
  AND2_X1   g248(.A1(new_n449), .A2(new_n375), .ZN(new_n450));
  NAND2_X1  g249(.A1(G228gat), .A2(G233gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n413), .A2(new_n328), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n317), .B1(new_n453), .B2(KEYINPUT89), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(KEYINPUT89), .B2(new_n453), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n453), .A2(new_n316), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n451), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(G22gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n448), .B1(new_n460), .B2(KEYINPUT90), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(G22gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n460), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT90), .A3(new_n462), .A4(new_n448), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n414), .A2(new_n416), .A3(new_n418), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(new_n406), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n471), .A2(KEYINPUT39), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n432), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n404), .A2(new_n408), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n476), .A2(new_n406), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n476), .A2(KEYINPUT92), .A3(new_n406), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT39), .B(new_n471), .C1(new_n479), .C2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n469), .B1(new_n475), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n473), .A2(new_n474), .ZN(new_n483));
  AOI21_X1  g282(.A(KEYINPUT91), .B1(new_n472), .B2(new_n432), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n481), .B(new_n469), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n430), .B(new_n436), .C1(new_n482), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n439), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n331), .A2(new_n337), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  OR3_X1    g291(.A1(new_n439), .A2(new_n492), .A3(new_n488), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n439), .B2(new_n488), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n468), .B1(new_n487), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n445), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n499), .A2(KEYINPUT79), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(KEYINPUT79), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT34), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n322), .A2(new_n417), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n407), .B(new_n318), .C1(new_n321), .C2(new_n306), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G227gat), .A2(G233gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(KEYINPUT64), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n509), .A2(KEYINPUT34), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n511), .B1(new_n504), .B2(new_n505), .ZN(new_n512));
  OAI21_X1  g311(.A(KEYINPUT77), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n506), .A2(new_n510), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT77), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n504), .A2(new_n505), .B1(G227gat), .B2(G233gat), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n515), .B(new_n516), .C1(new_n503), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT33), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(KEYINPUT32), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G43gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(G71gat), .B(G99gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n523), .A2(new_n524), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT33), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n521), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT76), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT76), .A4(new_n529), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n514), .B1(new_n513), .B2(new_n518), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n520), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI221_X4 g337(.A(new_n514), .B1(new_n513), .B2(new_n518), .C1(new_n534), .C2(new_n535), .ZN(new_n539));
  OAI211_X1 g338(.A(new_n501), .B(new_n502), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n489), .A2(new_n490), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n433), .A2(new_n429), .A3(new_n434), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n438), .ZN(new_n543));
  INV_X1    g342(.A(new_n494), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n439), .A2(new_n492), .A3(new_n488), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n467), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n513), .A2(new_n518), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT78), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n549), .A2(new_n519), .A3(new_n534), .A4(new_n535), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT78), .A3(new_n548), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT36), .A4(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n540), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n498), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n552), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n468), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT35), .B1(new_n557), .B2(new_n546), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n467), .B1(new_n550), .B2(new_n552), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT35), .B1(new_n437), .B2(new_n438), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n495), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n248), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(G85gat), .A2(G92gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  INV_X1    g365(.A(G85gat), .ZN(new_n567));
  INV_X1    g366(.A(G92gat), .ZN(new_n568));
  AOI22_X1  g367(.A1(KEYINPUT8), .A2(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G99gat), .B(G106gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT101), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n229), .A2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G232gat), .A2(G233gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n228), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n575), .A2(KEYINPUT41), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n581), .B(KEYINPUT100), .Z(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(KEYINPUT102), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(KEYINPUT102), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n579), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G57gat), .B(G64gat), .Z(new_n589));
  INV_X1    g388(.A(KEYINPUT9), .ZN(new_n590));
  INV_X1    g389(.A(G71gat), .ZN(new_n591));
  INV_X1    g390(.A(G78gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(KEYINPUT99), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G71gat), .B(G78gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G127gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n207), .B1(new_n597), .B2(new_n598), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G155gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n604), .B(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n588), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n572), .B(new_n596), .Z(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n572), .A2(new_n596), .A3(KEYINPUT10), .ZN(new_n615));
  AOI22_X1  g414(.A1(new_n614), .A2(new_n615), .B1(G230gat), .B2(G233gat), .ZN(new_n616));
  INV_X1    g415(.A(G230gat), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n612), .A2(new_n617), .A3(new_n250), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT103), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n619), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n625), .A2(KEYINPUT104), .A3(new_n627), .ZN(new_n628));
  OR3_X1    g427(.A1(new_n619), .A2(KEYINPUT104), .A3(new_n626), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n611), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g431(.A1(new_n563), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n543), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G1gat), .ZN(G1324gat));
  INV_X1    g435(.A(new_n495), .ZN(new_n637));
  AND2_X1   g436(.A1(new_n563), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(new_n632), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT105), .Z(new_n640));
  XOR2_X1   g439(.A(KEYINPUT16), .B(G8gat), .Z(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT42), .ZN(new_n642));
  OAI22_X1  g441(.A1(new_n640), .A2(new_n206), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(KEYINPUT42), .B1(new_n640), .B2(new_n641), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT106), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(G1325gat));
  AOI21_X1  g448(.A(G15gat), .B1(new_n633), .B2(new_n556), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n540), .A2(new_n553), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(G15gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n652), .B(KEYINPUT107), .Z(new_n653));
  AOI21_X1  g452(.A(new_n650), .B1(new_n633), .B2(new_n653), .ZN(G1326gat));
  NAND2_X1  g453(.A1(new_n633), .A2(new_n467), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT43), .B(G22gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT108), .B(KEYINPUT109), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(G1327gat));
  AOI21_X1  g458(.A(new_n341), .B1(KEYINPUT37), .B2(new_n351), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n443), .B1(new_n660), .B2(new_n440), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n353), .A2(KEYINPUT95), .A3(new_n441), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n496), .B1(new_n663), .B2(new_n339), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n540), .A2(new_n547), .A3(new_n553), .ZN(new_n665));
  AND4_X1   g464(.A1(new_n468), .A2(new_n556), .A3(new_n495), .A4(new_n560), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT35), .ZN(new_n667));
  INV_X1    g466(.A(new_n546), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n667), .B1(new_n559), .B2(new_n668), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n664), .A2(new_n665), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n588), .ZN(new_n671));
  INV_X1    g470(.A(new_n609), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(new_n631), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n247), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n675), .A2(new_n217), .A3(new_n634), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT45), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT112), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n588), .B(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT111), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n558), .A2(new_n682), .A3(new_n561), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT111), .B1(new_n666), .B2(new_n669), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n681), .B1(new_n685), .B2(new_n555), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687));
  INV_X1    g486(.A(new_n588), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n555), .B2(new_n562), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n689), .B2(new_n680), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n671), .A2(KEYINPUT110), .A3(KEYINPUT44), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n686), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n692), .A2(new_n543), .A3(new_n674), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n677), .B1(new_n693), .B2(new_n217), .ZN(G1328gat));
  NOR2_X1   g493(.A1(new_n692), .A2(new_n674), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n218), .B1(new_n695), .B2(new_n637), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n638), .A2(new_n218), .A3(new_n588), .A4(new_n673), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT46), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n696), .A2(new_n698), .ZN(G1329gat));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n651), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(G43gat), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(KEYINPUT113), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n673), .A2(new_n588), .ZN(new_n703));
  INV_X1    g502(.A(new_n556), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n703), .A2(G43gat), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n563), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT114), .Z(new_n707));
  OR2_X1    g506(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n701), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n701), .A2(new_n706), .A3(new_n708), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n702), .A2(new_n709), .B1(new_n710), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n467), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n468), .A2(G50gat), .ZN(new_n713));
  AOI22_X1  g512(.A1(new_n712), .A2(G50gat), .B1(new_n675), .B2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g514(.A1(new_n685), .A2(new_n555), .ZN(new_n716));
  AND4_X1   g515(.A1(new_n248), .A2(new_n716), .A3(new_n610), .A4(new_n631), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n634), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT115), .B(G57gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n637), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  NAND3_X1  g523(.A1(new_n717), .A2(new_n591), .A3(new_n556), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n717), .A2(new_n651), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n591), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g527(.A1(new_n717), .A2(new_n467), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G78gat), .ZN(G1335gat));
  INV_X1    g529(.A(KEYINPUT116), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n247), .A2(new_n672), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n631), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(new_n692), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n681), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT110), .B1(new_n671), .B2(KEYINPUT44), .ZN(new_n737));
  AOI211_X1 g536(.A(new_n687), .B(new_n680), .C1(new_n670), .C2(new_n588), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n733), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(KEYINPUT116), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n734), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n543), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n716), .A2(new_n588), .A3(new_n732), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT51), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n631), .A2(new_n567), .A3(new_n634), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT117), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n745), .B2(new_n747), .ZN(G1336gat));
  OR4_X1    g547(.A1(G92gat), .A2(new_n745), .A3(new_n495), .A4(new_n630), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n739), .A2(new_n740), .ZN(new_n751));
  OAI21_X1  g550(.A(G92gat), .B1(new_n751), .B2(new_n495), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G92gat), .B1(new_n742), .B2(new_n495), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n749), .A2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(new_n750), .ZN(G1337gat));
  INV_X1    g555(.A(new_n651), .ZN(new_n757));
  OAI21_X1  g556(.A(G99gat), .B1(new_n742), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n704), .A2(new_n630), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OR2_X1    g559(.A1(new_n760), .A2(G99gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n758), .B1(new_n745), .B2(new_n761), .ZN(G1338gat));
  OR3_X1    g561(.A1(new_n468), .A2(G106gat), .A3(new_n630), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n766));
  OAI21_X1  g565(.A(G106gat), .B1(new_n751), .B2(new_n468), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n734), .A2(new_n467), .A3(new_n741), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n765), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT118), .B1(new_n771), .B2(KEYINPUT53), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n764), .B1(new_n769), .B2(G106gat), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774));
  NOR3_X1   g573(.A1(new_n773), .A2(new_n774), .A3(new_n766), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n768), .B1(new_n772), .B2(new_n775), .ZN(G1339gat));
  NOR3_X1   g575(.A1(new_n611), .A2(new_n247), .A3(new_n631), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n626), .B1(new_n616), .B2(new_n778), .ZN(new_n779));
  OR2_X1    g578(.A1(new_n616), .A2(new_n778), .ZN(new_n780));
  AND4_X1   g579(.A1(G230gat), .A2(new_n614), .A3(G233gat), .A4(new_n615), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT119), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n627), .A3(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n230), .A2(new_n231), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n235), .A2(new_n236), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n242), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT120), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n246), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n248), .A2(new_n787), .B1(new_n630), .B2(new_n794), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n588), .B(KEYINPUT112), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n787), .A2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n679), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n777), .B1(new_n800), .B2(new_n609), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(new_n543), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n495), .A3(new_n559), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(new_n248), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(new_n378), .ZN(G1340gat));
  NOR2_X1   g604(.A1(new_n803), .A2(new_n630), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(new_n376), .ZN(G1341gat));
  NOR2_X1   g606(.A1(new_n803), .A2(new_n609), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT121), .B(G127gat), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n808), .B(new_n809), .ZN(G1342gat));
  NOR2_X1   g609(.A1(new_n803), .A2(new_n688), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n381), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n387), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n812), .B1(KEYINPUT56), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(KEYINPUT56), .B2(new_n813), .ZN(G1343gat));
  NOR2_X1   g614(.A1(new_n651), .A2(new_n468), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n248), .A2(G141gat), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n802), .A2(new_n495), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n651), .A2(new_n543), .A3(new_n637), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n801), .B2(new_n468), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n468), .A2(new_n821), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n795), .A2(new_n688), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n672), .B1(new_n824), .B2(new_n799), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(new_n777), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n820), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n361), .B1(new_n827), .B2(new_n247), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT122), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n818), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI211_X1 g629(.A(KEYINPUT122), .B(new_n361), .C1(new_n827), .C2(new_n247), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT58), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT58), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n835), .A2(KEYINPUT123), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT123), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n828), .A2(new_n837), .A3(new_n834), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n832), .B1(new_n836), .B2(new_n838), .ZN(G1344gat));
  AND3_X1   g638(.A1(new_n802), .A2(new_n495), .A3(new_n816), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n367), .A2(new_n369), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(new_n841), .A3(new_n631), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843));
  INV_X1    g642(.A(new_n824), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n787), .A2(new_n688), .A3(new_n794), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n609), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n777), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n468), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n467), .A2(KEYINPUT57), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n848), .A2(KEYINPUT57), .B1(new_n801), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n631), .A3(new_n819), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n843), .B1(new_n851), .B2(G148gat), .ZN(new_n852));
  AOI211_X1 g651(.A(KEYINPUT59), .B(new_n841), .C1(new_n827), .C2(new_n631), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(G1345gat));
  AND2_X1   g653(.A1(new_n840), .A2(new_n672), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(G155gat), .B1(new_n855), .B2(new_n856), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n609), .A2(new_n354), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n857), .A2(new_n858), .B1(new_n827), .B2(new_n859), .ZN(G1346gat));
  NAND2_X1  g659(.A1(new_n827), .A2(new_n679), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n355), .B1(new_n861), .B2(KEYINPUT125), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(KEYINPUT125), .B2(new_n861), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n355), .A3(new_n588), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1347gat));
  NOR2_X1   g664(.A1(new_n801), .A2(new_n634), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n801), .A2(KEYINPUT126), .A3(new_n634), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n637), .B(new_n559), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(new_n248), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n495), .A2(new_n467), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n866), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n704), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n248), .A2(new_n254), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n871), .A2(new_n254), .B1(new_n874), .B2(new_n875), .ZN(G1348gat));
  NOR3_X1   g675(.A1(new_n873), .A2(new_n253), .A3(new_n760), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n870), .A2(new_n630), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n266), .ZN(G1349gat));
  NAND2_X1  g678(.A1(new_n874), .A2(new_n672), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(G183gat), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n672), .A2(new_n280), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n881), .B1(new_n870), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT60), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT60), .ZN(new_n885));
  OAI211_X1 g684(.A(new_n881), .B(new_n885), .C1(new_n870), .C2(new_n882), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(G1350gat));
  INV_X1    g686(.A(KEYINPUT61), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n874), .A2(new_n588), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n888), .B1(new_n889), .B2(G190gat), .ZN(new_n890));
  AOI211_X1 g689(.A(KEYINPUT61), .B(new_n259), .C1(new_n874), .C2(new_n588), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n679), .A2(new_n259), .ZN(new_n892));
  OAI22_X1  g691(.A1(new_n890), .A2(new_n891), .B1(new_n870), .B2(new_n892), .ZN(G1351gat));
  NOR3_X1   g692(.A1(new_n651), .A2(new_n634), .A3(new_n495), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n850), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(G197gat), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(new_n248), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n868), .A2(new_n869), .ZN(new_n898));
  AND2_X1   g697(.A1(new_n898), .A2(new_n637), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n247), .A3(new_n816), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n897), .B1(new_n900), .B2(new_n896), .ZN(G1352gat));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n630), .A2(G204gat), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n899), .A2(new_n902), .A3(new_n816), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n850), .A2(new_n631), .A3(new_n894), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(G204gat), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n898), .A2(new_n637), .A3(new_n816), .ZN(new_n907));
  INV_X1    g706(.A(new_n903), .ZN(new_n908));
  OAI21_X1  g707(.A(KEYINPUT62), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n904), .A2(new_n906), .A3(new_n909), .ZN(G1353gat));
  NAND3_X1  g709(.A1(new_n850), .A2(new_n672), .A3(new_n894), .ZN(new_n911));
  AND4_X1   g710(.A1(KEYINPUT127), .A2(new_n911), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n912));
  OAI21_X1  g711(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n911), .A2(new_n914), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n609), .A2(G211gat), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n912), .A2(new_n915), .B1(new_n907), .B2(new_n916), .ZN(G1354gat));
  OAI21_X1  g716(.A(G218gat), .B1(new_n895), .B2(new_n688), .ZN(new_n918));
  OR2_X1    g717(.A1(new_n796), .A2(G218gat), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n907), .B2(new_n919), .ZN(G1355gat));
endmodule


