//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(new_n207), .A2(new_n208), .B1(new_n210), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n214), .B1(new_n208), .B2(new_n207), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n205), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT64), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n215), .B(new_n224), .C1(KEYINPUT1), .C2(new_n222), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XOR2_X1   g0029(.A(G250), .B(G257), .Z(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XOR2_X1   g0033(.A(G68), .B(G77), .Z(new_n234));
  XNOR2_X1  g0034(.A(G50), .B(G58), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  INV_X1    g0040(.A(KEYINPUT66), .ZN(new_n241));
  INV_X1    g0041(.A(G33), .ZN(new_n242));
  OAI21_X1  g0042(.A(new_n241), .B1(new_n205), .B2(new_n242), .ZN(new_n243));
  NAND4_X1  g0043(.A1(KEYINPUT66), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G1), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n245), .A2(G13), .A3(G20), .ZN(new_n246));
  NAND4_X1  g0046(.A1(new_n243), .A2(new_n211), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT69), .ZN(new_n248));
  OAI21_X1  g0048(.A(new_n248), .B1(new_n212), .B2(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n245), .A2(KEYINPUT69), .A3(G20), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G20), .A2(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n212), .A2(G33), .ZN(new_n257));
  XNOR2_X1  g0057(.A(KEYINPUT15), .B(G87), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n253), .B1(new_n254), .B2(new_n256), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n243), .A2(new_n211), .A3(new_n244), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n246), .ZN(new_n262));
  INV_X1    g0062(.A(G77), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n252), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G238), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT3), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n242), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1698), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G232), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  INV_X1    g0077(.A(G107), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT70), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G107), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n271), .B(new_n276), .C1(new_n277), .C2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT65), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT65), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G41), .ZN(new_n289));
  INV_X1    g0089(.A(G45), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G274), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G1), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n211), .ZN(new_n295));
  NAND2_X1  g0095(.A1(G33), .A2(G41), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n245), .B1(G41), .B2(G45), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n294), .B1(G244), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n285), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n265), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n270), .A2(G223), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n275), .A2(G222), .B1(new_n268), .B2(G77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n284), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n294), .B1(G226), .B2(new_n299), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G169), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(G58), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT67), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n254), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT68), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n257), .B(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n326));
  INV_X1    g0126(.A(G150), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n325), .B(new_n326), .C1(new_n327), .C2(new_n256), .ZN(new_n328));
  INV_X1    g0128(.A(G50), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n328), .A2(new_n260), .B1(new_n329), .B2(new_n262), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n251), .A2(G50), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G169), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n302), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n301), .A2(new_n316), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n265), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n308), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n330), .A2(KEYINPUT9), .A3(new_n331), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n314), .A2(G200), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n339), .B(new_n340), .C1(new_n303), .C2(new_n314), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT9), .B1(new_n330), .B2(new_n331), .ZN(new_n342));
  NOR3_X1   g0142(.A1(new_n341), .A2(KEYINPUT10), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT10), .B1(new_n341), .B2(new_n342), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT17), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n254), .A2(new_n321), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n249), .A2(new_n250), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n348), .A2(KEYINPUT75), .A3(new_n349), .A4(new_n319), .ZN(new_n350));
  INV_X1    g0150(.A(new_n247), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT75), .B1(new_n322), .B2(new_n349), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n352), .A2(new_n353), .B1(new_n246), .B2(new_n322), .ZN(new_n354));
  INV_X1    g0154(.A(G68), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n273), .A2(new_n212), .A3(new_n274), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n274), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n355), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n318), .A2(new_n355), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n361), .B2(new_n201), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n255), .A2(G159), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT16), .B1(new_n360), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(KEYINPUT7), .B1(new_n268), .B2(new_n212), .ZN(new_n366));
  INV_X1    g0166(.A(new_n359), .ZN(new_n367));
  OAI21_X1  g0167(.A(G68), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT16), .ZN(new_n369));
  INV_X1    g0169(.A(new_n364), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n354), .B1(new_n372), .B2(new_n260), .ZN(new_n373));
  OAI211_X1 g0173(.A(G223), .B(new_n269), .C1(new_n266), .C2(new_n267), .ZN(new_n374));
  OAI211_X1 g0174(.A(G226), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n375));
  INV_X1    g0175(.A(G87), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n374), .B(new_n375), .C1(new_n242), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n284), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n291), .A2(new_n293), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n297), .A2(G232), .A3(new_n298), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(new_n382), .A3(new_n303), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n284), .B2(new_n377), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(G200), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n347), .B1(new_n373), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n369), .B1(new_n368), .B2(new_n370), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n360), .A2(KEYINPUT16), .A3(new_n364), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n260), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n354), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n389), .A2(new_n385), .A3(new_n347), .A4(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT76), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n373), .A2(KEYINPUT76), .A3(new_n347), .A4(new_n385), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n386), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n384), .A2(G179), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n334), .B2(new_n384), .ZN(new_n397));
  INV_X1    g0197(.A(new_n260), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n398), .B1(new_n365), .B2(new_n371), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n397), .B1(new_n399), .B2(new_n354), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT18), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n397), .B(new_n402), .C1(new_n399), .C2(new_n354), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  OAI211_X1 g0206(.A(G232), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n407));
  OAI211_X1 g0207(.A(G226), .B(new_n269), .C1(new_n266), .C2(new_n267), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT71), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT71), .B1(new_n275), .B2(G226), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n284), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n294), .B1(G238), .B2(new_n299), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT13), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G169), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT14), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n412), .A2(KEYINPUT72), .A3(new_n413), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT72), .B1(new_n412), .B2(new_n413), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT13), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(G179), .A3(new_n416), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT14), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n419), .A2(new_n426), .A3(G169), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n421), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n324), .A2(G77), .ZN(new_n429));
  AOI22_X1  g0229(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n355), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n398), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT11), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n251), .A2(G68), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(KEYINPUT11), .ZN(new_n434));
  INV_X1    g0234(.A(G13), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G1), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(G20), .A3(new_n355), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT12), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n432), .A2(new_n433), .A3(new_n434), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n428), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n346), .A2(new_n405), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n439), .B1(new_n419), .B2(G200), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT73), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n303), .B1(new_n414), .B2(new_n415), .ZN(new_n444));
  AND3_X1   g0244(.A1(new_n424), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n443), .B1(new_n424), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT74), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT74), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n442), .B(new_n449), .C1(new_n445), .C2(new_n446), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT24), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n212), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT22), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n277), .A2(new_n456), .A3(new_n212), .A4(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT83), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT23), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n460), .A2(new_n278), .A3(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(G20), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n279), .B2(new_n281), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n458), .A2(new_n459), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n459), .B1(new_n458), .B2(new_n465), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n453), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(G20), .B1(new_n273), .B2(new_n274), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n456), .B1(new_n469), .B2(G87), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n454), .A2(KEYINPUT22), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n465), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n458), .A2(new_n459), .A3(new_n465), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n473), .A2(KEYINPUT24), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n468), .A2(new_n475), .A3(new_n260), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n262), .A2(new_n278), .ZN(new_n477));
  XNOR2_X1  g0277(.A(new_n477), .B(KEYINPUT25), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n242), .A2(G1), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n247), .A2(new_n278), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(G250), .B(new_n269), .C1(new_n266), .C2(new_n267), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G294), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n284), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n287), .A2(new_n289), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT79), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n286), .A3(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n245), .A2(G45), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n286), .A2(KEYINPUT5), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(KEYINPUT79), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n292), .B1(new_n295), .B2(new_n296), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n489), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT79), .B1(new_n488), .B2(G41), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n290), .A2(G1), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT5), .B1(new_n287), .B2(new_n289), .ZN(new_n500));
  OAI211_X1 g0300(.A(G264), .B(new_n297), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n486), .A2(new_n496), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n305), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(G190), .B2(new_n502), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n476), .A2(new_n481), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n486), .A2(G179), .A3(new_n496), .A4(new_n501), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n502), .A2(G169), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n502), .A2(KEYINPUT84), .A3(G169), .ZN(new_n511));
  AOI221_X4 g0311(.A(new_n506), .B1(new_n510), .B2(new_n511), .C1(new_n476), .C2(new_n481), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n476), .A2(new_n481), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT85), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(G257), .B(new_n297), .C1(new_n499), .C2(new_n500), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n517), .A2(new_n496), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(G1698), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(G244), .C1(new_n267), .C2(new_n266), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  INV_X1    g0322(.A(G244), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n523), .B1(new_n273), .B2(new_n274), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n521), .B(new_n522), .C1(new_n524), .C2(KEYINPUT4), .ZN(new_n525));
  OAI21_X1  g0325(.A(G250), .B1(new_n266), .B2(new_n267), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n269), .B1(new_n526), .B2(KEYINPUT4), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n284), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n518), .A2(KEYINPUT80), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT80), .B1(new_n518), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g0330(.A(G190), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g0331(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n532));
  NAND2_X1  g0332(.A1(KEYINPUT77), .A2(KEYINPUT6), .ZN(new_n533));
  INV_X1    g0333(.A(G97), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n532), .B(new_n533), .C1(new_n534), .C2(G107), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  XNOR2_X1  g0336(.A(G97), .B(G107), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(G20), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n255), .A2(G77), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n282), .B1(new_n358), .B2(new_n359), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n260), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n247), .A2(new_n479), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n262), .A2(new_n534), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n528), .A2(KEYINPUT78), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT78), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n549), .B(new_n284), .C1(new_n525), .C2(new_n527), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n518), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G200), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n531), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n518), .A2(new_n528), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT80), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n518), .A2(new_n528), .A3(KEYINPUT80), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n334), .A3(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n548), .A2(new_n316), .A3(new_n518), .A4(new_n550), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n546), .ZN(new_n560));
  NOR2_X1   g0360(.A1(G87), .A2(G97), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n279), .A2(new_n281), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n212), .B1(new_n406), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n277), .A2(new_n212), .A3(G68), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n563), .B1(new_n406), .B2(G20), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n260), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n543), .A2(G87), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n258), .A2(new_n262), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n492), .A2(G250), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n293), .A2(G45), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n284), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(G238), .B(new_n269), .C1(new_n266), .C2(new_n267), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n577));
  NAND2_X1  g0377(.A1(G33), .A2(G116), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI211_X1 g0379(.A(new_n303), .B(new_n575), .C1(new_n284), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n284), .ZN(new_n582));
  INV_X1    g0382(.A(new_n575), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G200), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(G179), .A3(new_n583), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n575), .B1(new_n579), .B2(new_n284), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n334), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n543), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n569), .B(new_n571), .C1(new_n258), .C2(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n581), .A2(new_n585), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n553), .A2(new_n560), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT20), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n242), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(G20), .B1(new_n594), .B2(new_n522), .ZN(new_n595));
  INV_X1    g0395(.A(G116), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n212), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n398), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n260), .B(KEYINPUT20), .C1(new_n595), .C2(new_n597), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n246), .A2(G116), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n543), .B2(G116), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n268), .A2(G303), .ZN(new_n606));
  OAI211_X1 g0406(.A(G264), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n607));
  OAI211_X1 g0407(.A(G257), .B(new_n269), .C1(new_n266), .C2(new_n267), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT81), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT81), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n606), .A2(new_n611), .A3(new_n607), .A4(new_n608), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n284), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(G270), .B(new_n297), .C1(new_n499), .C2(new_n500), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n614), .A2(new_n496), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(G190), .ZN(new_n617));
  AOI21_X1  g0417(.A(G200), .B1(new_n613), .B2(new_n615), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n605), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(KEYINPUT82), .A2(KEYINPUT21), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n334), .B1(new_n601), .B2(new_n603), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n616), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n616), .A3(new_n621), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n604), .A2(G179), .A3(new_n613), .A4(new_n615), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n619), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n592), .A2(new_n627), .ZN(new_n628));
  AND4_X1   g0428(.A1(new_n452), .A2(new_n505), .A3(new_n516), .A4(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n345), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n343), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT90), .ZN(new_n632));
  INV_X1    g0432(.A(new_n404), .ZN(new_n633));
  INV_X1    g0433(.A(new_n337), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n439), .A2(new_n428), .B1(new_n447), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n395), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n632), .A2(new_n636), .B1(new_n332), .B2(new_n317), .ZN(new_n637));
  INV_X1    g0437(.A(new_n452), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n559), .A2(new_n546), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n639), .A2(new_n591), .A3(KEYINPUT26), .A4(new_n558), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT89), .ZN(new_n641));
  NOR3_X1   g0441(.A1(new_n529), .A2(new_n530), .A3(G169), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n559), .A2(new_n546), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT89), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(KEYINPUT26), .A4(new_n591), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n585), .A2(KEYINPUT86), .ZN(new_n648));
  OR3_X1    g0448(.A1(new_n587), .A2(KEYINPUT86), .A3(new_n305), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n581), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n588), .A2(new_n590), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n647), .B1(new_n560), .B2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n641), .A2(new_n646), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n651), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n656));
  INV_X1    g0456(.A(new_n481), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n473), .A2(new_n474), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n398), .B1(new_n658), .B2(new_n453), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(new_n475), .ZN(new_n660));
  INV_X1    g0460(.A(new_n514), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT87), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT87), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n513), .A2(new_n663), .A3(new_n514), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n656), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n650), .A2(new_n651), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n553), .A3(new_n560), .A4(new_n505), .ZN(new_n667));
  OAI21_X1  g0467(.A(KEYINPUT88), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n513), .A2(new_n663), .A3(new_n514), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n663), .B1(new_n513), .B2(new_n514), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT88), .ZN(new_n673));
  INV_X1    g0473(.A(new_n667), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n655), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n637), .B1(new_n638), .B2(new_n676), .ZN(G369));
  NAND2_X1  g0477(.A1(new_n436), .A2(new_n212), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n605), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n669), .B2(new_n619), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n686), .B1(new_n669), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n516), .A2(new_n505), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n513), .A2(new_n683), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n513), .A2(new_n514), .A3(new_n683), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n669), .A2(new_n683), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n690), .A2(new_n691), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n662), .A2(new_n664), .A3(new_n684), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n206), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n487), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G1), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n282), .A2(new_n596), .A3(new_n561), .ZN(new_n706));
  OAI22_X1  g0506(.A1(new_n705), .A2(new_n706), .B1(new_n209), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT94), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT93), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n581), .A2(new_n585), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n651), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n710), .B(new_n647), .C1(new_n560), .C2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n666), .A2(new_n644), .A3(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n639), .A2(new_n591), .A3(new_n558), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n710), .B1(new_n716), .B2(new_n647), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n709), .B(new_n651), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n515), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n513), .A2(KEYINPUT85), .A3(new_n514), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n674), .B1(new_n721), .B2(new_n656), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n647), .B1(new_n560), .B2(new_n712), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT93), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n713), .A3(new_n714), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n709), .B1(new_n726), .B2(new_n651), .ZN(new_n727));
  OAI211_X1 g0527(.A(KEYINPUT29), .B(new_n684), .C1(new_n723), .C2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n676), .A2(new_n683), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n728), .B1(new_n729), .B2(KEYINPUT29), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n616), .A2(new_n316), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n587), .A2(new_n501), .A3(new_n486), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n732), .C1(new_n530), .C2(new_n529), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AND4_X1   g0536(.A1(new_n316), .A2(new_n616), .A3(new_n502), .A4(new_n584), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n733), .A2(new_n734), .B1(new_n551), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n684), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n628), .A2(new_n516), .A3(new_n505), .A4(new_n684), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(new_n740), .B2(KEYINPUT31), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n683), .A2(KEYINPUT31), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT92), .ZN(new_n744));
  OR2_X1    g0544(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n735), .B1(new_n738), .B2(new_n744), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n741), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G330), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n730), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n708), .B1(new_n750), .B2(G1), .ZN(G364));
  NOR2_X1   g0551(.A1(new_n435), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n705), .B1(G45), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n687), .A2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT95), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n756), .B1(new_n755), .B2(new_n754), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n689), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT96), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n211), .B1(G20), .B2(new_n334), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n316), .A2(new_n305), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n212), .A2(G190), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n268), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n212), .A2(new_n303), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G179), .A3(new_n305), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n763), .A2(G179), .A3(new_n305), .ZN(new_n769));
  INV_X1    g0569(.A(G311), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n767), .A2(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G190), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n765), .B(new_n771), .C1(G294), .C2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n305), .A2(G179), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n763), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G283), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n766), .A2(new_n762), .ZN(new_n780));
  INV_X1    g0580(.A(G326), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n766), .A2(new_n776), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n763), .A2(new_n772), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n779), .B(new_n784), .C1(G329), .C2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n775), .A2(new_n787), .A3(KEYINPUT100), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n329), .A2(new_n780), .B1(new_n769), .B2(new_n263), .ZN(new_n789));
  INV_X1    g0589(.A(new_n767), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(G58), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n785), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(KEYINPUT99), .B(KEYINPUT32), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n774), .A2(G97), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n277), .B1(new_n764), .B2(new_n355), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n782), .A2(new_n376), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n777), .A2(new_n278), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n797), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n791), .A2(new_n795), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT100), .B1(new_n775), .B2(new_n787), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n760), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n753), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n277), .A2(new_n206), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT97), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n807), .A2(G355), .B1(new_n596), .B2(new_n702), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n702), .A2(new_n277), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n210), .A2(G45), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n236), .B2(G45), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n808), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G13), .A2(G33), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n212), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT98), .ZN(new_n816));
  INV_X1    g0616(.A(new_n760), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n805), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n804), .B(new_n820), .C1(new_n687), .C2(new_n816), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n759), .A2(new_n821), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT101), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G396));
  NAND2_X1  g0624(.A1(new_n634), .A2(new_n684), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n265), .A2(new_n683), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n337), .B1(new_n307), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  XNOR2_X1  g0629(.A(new_n729), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n749), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT102), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(KEYINPUT102), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n830), .A2(new_n749), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n832), .A2(new_n805), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n814), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n817), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n753), .B1(G77), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n767), .A2(new_n839), .B1(new_n769), .B2(new_n596), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n780), .A2(new_n783), .B1(new_n764), .B2(new_n778), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n777), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n277), .B1(new_n843), .B2(G87), .ZN(new_n844));
  INV_X1    g0644(.A(new_n782), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G107), .A2(new_n845), .B1(new_n786), .B2(G311), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n842), .A2(new_n796), .A3(new_n844), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n780), .ZN(new_n848));
  INV_X1    g0648(.A(new_n769), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G137), .A2(new_n848), .B1(new_n849), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n851), .B2(new_n767), .C1(new_n327), .C2(new_n764), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT34), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n277), .B1(new_n782), .B2(new_n329), .ZN(new_n855));
  INV_X1    g0655(.A(G132), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n777), .A2(new_n355), .B1(new_n785), .B2(new_n856), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n855), .B(new_n857), .C1(G58), .C2(new_n774), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n852), .A2(new_n853), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n847), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n838), .B1(new_n861), .B2(new_n760), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n829), .B2(new_n836), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n835), .A2(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n752), .A2(new_n245), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n728), .B(new_n452), .C1(new_n729), .C2(KEYINPUT29), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n637), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(KEYINPUT105), .ZN(new_n868));
  INV_X1    g0668(.A(new_n681), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n399), .B2(new_n354), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n395), .B2(new_n404), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n373), .A2(new_n385), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n873), .A2(new_n400), .A3(new_n870), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT37), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n873), .A2(new_n400), .A3(new_n876), .A4(new_n870), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n872), .A2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n878), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n439), .A2(new_n683), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n440), .A2(new_n447), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n428), .B1(new_n448), .B2(new_n450), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(new_n884), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n676), .A2(new_n683), .A3(new_n828), .ZN(new_n888));
  INV_X1    g0688(.A(new_n825), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n883), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n633), .A2(new_n869), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT39), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n881), .B2(new_n882), .ZN(new_n894));
  INV_X1    g0694(.A(new_n882), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT104), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n872), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(KEYINPUT104), .B(new_n871), .C1(new_n395), .C2(new_n404), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT103), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n878), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n875), .A2(KEYINPUT103), .A3(new_n877), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n897), .A2(new_n898), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n895), .B1(new_n902), .B2(new_n880), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n894), .B1(new_n903), .B2(new_n893), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n440), .A2(new_n683), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n890), .B(new_n892), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n868), .B(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n739), .A2(KEYINPUT31), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n741), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n910), .A2(new_n829), .A3(new_n883), .A4(new_n887), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n887), .B(new_n829), .C1(new_n741), .C2(new_n909), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n902), .A2(new_n880), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n915), .B2(new_n882), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n911), .A2(new_n912), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n910), .A2(new_n452), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n917), .B(new_n918), .Z(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n865), .B1(new_n908), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n908), .B2(new_n920), .ZN(new_n922));
  NOR3_X1   g0722(.A1(new_n209), .A2(new_n263), .A3(new_n361), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n355), .A2(G50), .ZN(new_n924));
  OAI211_X1 g0724(.A(G1), .B(new_n435), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n536), .A2(new_n537), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n926), .A2(new_n535), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n927), .A2(KEYINPUT35), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n927), .A2(KEYINPUT35), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n928), .A2(G116), .A3(new_n213), .A4(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT36), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n925), .A3(new_n931), .ZN(G367));
  OAI211_X1 g0732(.A(new_n553), .B(new_n560), .C1(new_n547), .C2(new_n684), .ZN(new_n933));
  OR3_X1    g0733(.A1(new_n697), .A2(KEYINPUT42), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT42), .B1(new_n697), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n560), .B1(new_n516), .B2(new_n933), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n684), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n572), .A2(new_n683), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n590), .B2(new_n588), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n652), .B2(new_n938), .ZN(new_n940));
  XNOR2_X1  g0740(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n934), .A2(new_n935), .A3(new_n937), .A4(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT107), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT107), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n942), .B1(KEYINPUT43), .B2(new_n940), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n944), .A2(new_n945), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n644), .A2(new_n683), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n933), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n695), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n949), .B(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n703), .B(KEYINPUT41), .Z(new_n955));
  INV_X1    g0755(.A(KEYINPUT111), .ZN(new_n956));
  XOR2_X1   g0756(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n957));
  INV_X1    g0757(.A(KEYINPUT110), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n699), .A2(new_n958), .A3(new_n952), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n699), .B2(new_n952), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(new_n957), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n963), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n697), .A2(new_n698), .A3(new_n951), .ZN(new_n966));
  XNOR2_X1  g0766(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n962), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n969), .A2(new_n689), .A3(new_n694), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n962), .A2(new_n965), .A3(new_n695), .A4(new_n968), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n697), .B1(new_n694), .B2(new_n696), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n689), .B(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(new_n750), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n956), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n970), .A2(new_n975), .A3(KEYINPUT111), .A4(new_n971), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n955), .B1(new_n979), .B2(new_n750), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n752), .A2(G45), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(G1), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(KEYINPUT112), .Z(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n954), .B1(new_n980), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n232), .A2(new_n810), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n819), .B1(new_n206), .B2(new_n258), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n767), .A2(new_n783), .B1(new_n764), .B2(new_n839), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n277), .B(new_n988), .C1(G317), .C2(new_n786), .ZN(new_n989));
  INV_X1    g0789(.A(new_n774), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(new_n282), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n845), .A2(G116), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n770), .A2(new_n780), .B1(new_n769), .B2(new_n778), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n777), .A2(new_n534), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n989), .A2(new_n991), .A3(new_n993), .A4(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(G137), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n777), .A2(new_n263), .B1(new_n785), .B2(new_n998), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n268), .B(new_n999), .C1(G58), .C2(new_n845), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n767), .A2(new_n327), .B1(new_n780), .B2(new_n851), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n329), .A2(new_n769), .B1(new_n764), .B2(new_n792), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1000), .B(new_n1003), .C1(new_n355), .C2(new_n990), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n997), .A2(new_n1004), .A3(KEYINPUT47), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n760), .ZN(new_n1006));
  AOI21_X1  g0806(.A(KEYINPUT47), .B1(new_n997), .B2(new_n1004), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n753), .B1(new_n986), .B2(new_n987), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT113), .Z(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n816), .B2(new_n940), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n985), .A2(new_n1010), .ZN(G387));
  NAND2_X1  g0811(.A1(new_n974), .A2(new_n984), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n694), .A2(new_n816), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n254), .A2(G50), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT50), .Z(new_n1015));
  OAI21_X1  g0815(.A(new_n290), .B1(new_n355), .B2(new_n263), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1015), .A2(new_n706), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n809), .B1(new_n229), .B2(new_n290), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n807), .A2(new_n706), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n206), .A2(G107), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n819), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G159), .A2(new_n848), .B1(new_n849), .B2(G68), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n329), .B2(new_n767), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n990), .A2(new_n258), .ZN(new_n1025));
  NOR4_X1   g0825(.A1(new_n1024), .A2(new_n268), .A3(new_n995), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n322), .A2(new_n763), .A3(new_n762), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n782), .A2(new_n263), .B1(new_n785), .B2(new_n327), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT114), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n277), .B1(new_n843), .B2(G116), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n990), .A2(new_n778), .B1(new_n782), .B2(new_n839), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n768), .A2(new_n780), .B1(new_n769), .B2(new_n783), .ZN(new_n1033));
  INV_X1    g0833(.A(G317), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n767), .A2(new_n1034), .B1(new_n764), .B2(new_n770), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1032), .B1(new_n1036), .B2(KEYINPUT48), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(KEYINPUT48), .B2(new_n1036), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1031), .B1(new_n781), .B2(new_n785), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n805), .B1(new_n1042), .B2(new_n760), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1022), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n976), .A2(new_n703), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n974), .A2(new_n750), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1012), .B1(new_n1013), .B2(new_n1044), .C1(new_n1045), .C2(new_n1046), .ZN(G393));
  AOI21_X1  g0847(.A(new_n704), .B1(new_n972), .B2(new_n976), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n979), .A2(new_n1048), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n767), .A2(new_n792), .B1(new_n780), .B2(new_n327), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1050), .B(KEYINPUT51), .Z(new_n1051));
  OAI22_X1  g0851(.A1(new_n782), .A2(new_n355), .B1(new_n785), .B2(new_n851), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n254), .A2(new_n769), .B1(new_n764), .B2(new_n329), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n277), .B1(new_n777), .B2(new_n376), .C1(new_n990), .C2(new_n263), .ZN(new_n1054));
  OR4_X1    g0854(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n767), .A2(new_n770), .B1(new_n780), .B2(new_n1034), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT52), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n839), .A2(new_n769), .B1(new_n782), .B2(new_n778), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n764), .A2(new_n783), .B1(new_n785), .B2(new_n768), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n277), .B(new_n799), .C1(G116), .C2(new_n774), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1057), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n817), .B1(new_n1055), .B2(new_n1062), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n239), .A2(new_n810), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n818), .B1(G97), .B2(new_n702), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n805), .B(new_n1063), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n951), .B2(new_n816), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n972), .B2(new_n983), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1049), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(G390));
  OAI211_X1 g0870(.A(G330), .B(new_n829), .C1(new_n741), .C2(new_n909), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n887), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n915), .A2(new_n893), .A3(new_n882), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n894), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1076), .B1(new_n1077), .B2(new_n906), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n915), .A2(new_n882), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n905), .B(KEYINPUT115), .Z(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n684), .B(new_n827), .C1(new_n723), .C2(new_n727), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n825), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n887), .A2(KEYINPUT116), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT116), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1085), .B(new_n885), .C1(new_n886), .C2(new_n884), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1081), .B1(new_n1083), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1073), .B1(new_n1078), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n910), .A2(G330), .A3(new_n452), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n866), .A2(new_n637), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n668), .A2(new_n675), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n655), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1094), .A2(new_n684), .A3(new_n829), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n825), .ZN(new_n1096));
  OAI211_X1 g0896(.A(G330), .B(new_n829), .C1(new_n741), .C2(new_n747), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1097), .A2(new_n1072), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n1098), .B2(new_n1073), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n748), .A2(G330), .A3(new_n829), .A4(new_n887), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1082), .A2(new_n825), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1071), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1091), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1072), .B1(new_n1095), .B2(new_n825), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n904), .B1(new_n1105), .B2(new_n905), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1083), .A2(new_n1087), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1081), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1106), .A2(new_n1109), .A3(new_n1100), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1089), .A2(new_n1104), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1089), .A2(new_n1104), .A3(new_n1110), .A4(KEYINPUT117), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1089), .A2(new_n1110), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1104), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n704), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1089), .A2(new_n1110), .A3(new_n984), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n753), .B1(new_n322), .B2(new_n837), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n769), .A2(new_n1122), .B1(new_n764), .B2(new_n998), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G159), .B2(new_n774), .ZN(new_n1124));
  XOR2_X1   g0924(.A(new_n1124), .B(KEYINPUT118), .Z(new_n1125));
  INV_X1    g0925(.A(G125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n782), .A2(new_n327), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT53), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n277), .B1(new_n1126), .B2(new_n785), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1128), .B2(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n848), .A2(G128), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n790), .A2(G132), .B1(new_n843), .B2(G50), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n990), .A2(new_n263), .B1(new_n767), .B2(new_n596), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT119), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n769), .A2(new_n534), .B1(new_n777), .B2(new_n355), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n1136), .A2(new_n277), .A3(new_n798), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n848), .A2(G283), .B1(new_n786), .B2(G294), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n1137), .B(new_n1138), .C1(new_n282), .C2(new_n764), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1125), .A2(new_n1133), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1121), .B1(new_n1140), .B2(new_n760), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n1076), .B2(new_n836), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1119), .A2(new_n1120), .A3(new_n1142), .ZN(G378));
  XOR2_X1   g0943(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1144));
  NAND2_X1  g0944(.A1(new_n332), .A2(new_n869), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n632), .A2(new_n333), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n632), .B2(new_n333), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1148), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1144), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1150), .A2(new_n1146), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1149), .A2(new_n1152), .A3(new_n814), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n753), .B1(G50), .B2(new_n837), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n998), .A2(new_n769), .B1(new_n764), .B2(new_n856), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT122), .Z(new_n1156));
  NOR2_X1   g0956(.A1(new_n990), .A2(new_n327), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n782), .A2(new_n1122), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n767), .A2(new_n1159), .B1(new_n780), .B2(new_n1126), .ZN(new_n1160));
  NOR4_X1   g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n242), .B(new_n286), .C1(new_n777), .C2(new_n792), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(G124), .B2(new_n786), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n268), .A2(new_n287), .A3(new_n289), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n777), .A2(new_n318), .B1(new_n785), .B2(new_n778), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1168), .B(new_n1169), .C1(G77), .C2(new_n845), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT121), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n258), .A2(new_n769), .B1(new_n764), .B2(new_n534), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n767), .A2(new_n278), .B1(new_n780), .B2(new_n596), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(G68), .C2(new_n774), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT58), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(KEYINPUT58), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1168), .B(new_n329), .C1(G33), .C2(G41), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT120), .Z(new_n1179));
  NAND4_X1  g0979(.A1(new_n1167), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1154), .B1(new_n1180), .B2(new_n760), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1153), .A2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT123), .ZN(new_n1183));
  NAND4_X1  g0983(.A1(new_n907), .A2(new_n1183), .A3(G330), .A4(new_n917), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n914), .A2(new_n916), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n883), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n912), .B1(new_n913), .B2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(G330), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT123), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n891), .B1(new_n1076), .B2(new_n905), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n890), .B(new_n1192), .C1(new_n1188), .C2(KEYINPUT123), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1184), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1191), .B1(new_n1184), .B2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1182), .B1(new_n1196), .B2(new_n983), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1091), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1115), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT57), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1091), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1196), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1197), .B1(new_n1205), .B2(new_n703), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(G375));
  OAI21_X1  g1007(.A(new_n753), .B1(G68), .B2(new_n837), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1087), .A2(new_n836), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n780), .A2(new_n856), .B1(new_n764), .B2(new_n1122), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n268), .B(new_n1210), .C1(G58), .C2(new_n843), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n790), .A2(G137), .B1(new_n845), .B2(G159), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n849), .A2(G150), .B1(new_n786), .B2(G128), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n774), .A2(G50), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n282), .A2(new_n769), .B1(new_n764), .B2(new_n596), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT124), .Z(new_n1217));
  OAI22_X1  g1017(.A1(new_n780), .A2(new_n839), .B1(new_n785), .B2(new_n783), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n767), .A2(new_n778), .B1(new_n782), .B2(new_n534), .ZN(new_n1219));
  OR4_X1    g1019(.A1(new_n1025), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n268), .B1(new_n777), .B2(new_n263), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT125), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1215), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1208), .B(new_n1209), .C1(new_n760), .C2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n984), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n955), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1117), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1225), .A2(new_n1198), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1226), .B1(new_n1228), .B2(new_n1229), .ZN(G381));
  INV_X1    g1030(.A(G378), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n985), .A2(new_n1069), .A3(new_n1010), .ZN(new_n1232));
  OR2_X1    g1032(.A1(G396), .A2(G393), .ZN(new_n1233));
  NOR4_X1   g1033(.A1(new_n1232), .A2(G384), .A3(G381), .A4(new_n1233), .ZN(new_n1234));
  AND2_X1   g1034(.A1(G375), .A2(KEYINPUT126), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G375), .A2(KEYINPUT126), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1231), .B(new_n1234), .C1(new_n1235), .C2(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n682), .A2(G213), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1231), .B(new_n1239), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(new_n1240), .A3(G213), .ZN(G409));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1229), .B(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1104), .A2(new_n704), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(KEYINPUT127), .A3(new_n1244), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1229), .A2(new_n1242), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1225), .A2(KEYINPUT60), .A3(new_n1198), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1244), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT127), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1245), .A2(new_n1250), .A3(new_n1226), .ZN(new_n1251));
  INV_X1    g1051(.A(G384), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1245), .A2(new_n1250), .A3(G384), .A4(new_n1226), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n704), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1257), .A2(new_n1231), .A3(new_n1197), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1197), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1199), .A2(new_n1227), .A3(new_n1201), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G378), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1238), .B(new_n1256), .C1(new_n1258), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT61), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1239), .A2(G2897), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1253), .A2(new_n1254), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1261), .B1(new_n1206), .B2(G378), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1268), .B1(new_n1269), .B2(new_n1239), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1200), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1203), .A2(new_n1196), .A3(KEYINPUT57), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n703), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(G378), .A3(new_n1259), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1261), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1238), .A4(new_n1256), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1263), .A2(new_n1264), .A3(new_n1270), .A4(new_n1278), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n823), .B(G393), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n985), .A2(new_n1010), .A3(new_n1069), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1069), .B1(new_n985), .B2(new_n1010), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1280), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1280), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1232), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1283), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1279), .A2(new_n1287), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1283), .A2(new_n1286), .A3(new_n1264), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1238), .A4(new_n1256), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT63), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1238), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1292), .B2(new_n1268), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1262), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1289), .B(new_n1290), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n1295), .ZN(G405));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1231), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1283), .A2(new_n1286), .A3(new_n1256), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1256), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1299));
  OAI211_X1 g1099(.A(new_n1274), .B(new_n1297), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1287), .A2(new_n1255), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1297), .A2(new_n1274), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1283), .A2(new_n1286), .A3(new_n1256), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(G402));
endmodule


