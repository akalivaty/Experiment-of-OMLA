

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U561 ( .A(KEYINPUT97), .ZN(n738) );
  INV_X1 U562 ( .A(KEYINPUT32), .ZN(n747) );
  NOR2_X1 U563 ( .A1(G2105), .A2(n548), .ZN(n904) );
  XOR2_X1 U564 ( .A(KEYINPUT95), .B(KEYINPUT30), .Z(n527) );
  NOR2_X1 U565 ( .A1(n983), .A2(n771), .ZN(n528) );
  XOR2_X1 U566 ( .A(n699), .B(KEYINPUT28), .Z(n529) );
  INV_X1 U567 ( .A(G168), .ZN(n730) );
  INV_X1 U568 ( .A(KEYINPUT31), .ZN(n734) );
  INV_X1 U569 ( .A(KEYINPUT89), .ZN(n725) );
  XNOR2_X1 U570 ( .A(n726), .B(n725), .ZN(n754) );
  OR2_X1 U571 ( .A1(n772), .A2(n528), .ZN(n806) );
  NOR2_X2 U572 ( .A1(G164), .A2(G1384), .ZN(n775) );
  NOR2_X1 U573 ( .A1(G651), .A2(n661), .ZN(n660) );
  NOR2_X1 U574 ( .A1(n598), .A2(n597), .ZN(n1003) );
  XOR2_X1 U575 ( .A(G543), .B(KEYINPUT0), .Z(n661) );
  NAND2_X1 U576 ( .A1(n660), .A2(G51), .ZN(n530) );
  XOR2_X1 U577 ( .A(KEYINPUT69), .B(n530), .Z(n533) );
  INV_X1 U578 ( .A(G651), .ZN(n537) );
  NOR2_X1 U579 ( .A1(G543), .A2(n537), .ZN(n531) );
  XOR2_X2 U580 ( .A(KEYINPUT1), .B(n531), .Z(n665) );
  NAND2_X1 U581 ( .A1(n665), .A2(G63), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U583 ( .A(KEYINPUT6), .B(n534), .ZN(n543) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT64), .ZN(n653) );
  NAND2_X1 U586 ( .A1(G89), .A2(n653), .ZN(n536) );
  XNOR2_X1 U587 ( .A(n536), .B(KEYINPUT4), .ZN(n539) );
  NOR2_X1 U588 ( .A1(n661), .A2(n537), .ZN(n652) );
  NAND2_X1 U589 ( .A1(G76), .A2(n652), .ZN(n538) );
  NAND2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U591 ( .A(KEYINPUT5), .B(n540), .Z(n541) );
  XNOR2_X1 U592 ( .A(KEYINPUT68), .B(n541), .ZN(n542) );
  NOR2_X1 U593 ( .A1(n543), .A2(n542), .ZN(n546) );
  XNOR2_X1 U594 ( .A(KEYINPUT71), .B(KEYINPUT7), .ZN(n544) );
  XNOR2_X1 U595 ( .A(n544), .B(KEYINPUT70), .ZN(n545) );
  XNOR2_X1 U596 ( .A(n546), .B(n545), .ZN(G168) );
  NOR2_X1 U597 ( .A1(G2104), .A2(G2105), .ZN(n547) );
  XOR2_X2 U598 ( .A(KEYINPUT17), .B(n547), .Z(n906) );
  AND2_X1 U599 ( .A1(G138), .A2(n906), .ZN(n555) );
  INV_X1 U600 ( .A(G2105), .ZN(n549) );
  INV_X1 U601 ( .A(G2104), .ZN(n548) );
  NAND2_X1 U602 ( .A1(G102), .A2(n904), .ZN(n553) );
  NOR2_X2 U603 ( .A1(n548), .A2(n549), .ZN(n898) );
  NAND2_X1 U604 ( .A1(G114), .A2(n898), .ZN(n551) );
  NOR2_X2 U605 ( .A1(G2104), .A2(n549), .ZN(n899) );
  NAND2_X1 U606 ( .A1(G126), .A2(n899), .ZN(n550) );
  AND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U609 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X2 U610 ( .A(n556), .B(KEYINPUT78), .ZN(G164) );
  NAND2_X1 U611 ( .A1(n906), .A2(G137), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G2104), .A2(G101), .ZN(n557) );
  OR2_X1 U613 ( .A1(G2105), .A2(n557), .ZN(n558) );
  XOR2_X1 U614 ( .A(KEYINPUT23), .B(n558), .Z(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G113), .A2(n898), .ZN(n562) );
  NAND2_X1 U617 ( .A1(G125), .A2(n899), .ZN(n561) );
  NAND2_X1 U618 ( .A1(n562), .A2(n561), .ZN(n563) );
  NOR2_X1 U619 ( .A1(n564), .A2(n563), .ZN(G160) );
  NAND2_X1 U620 ( .A1(n652), .A2(G72), .ZN(n566) );
  NAND2_X1 U621 ( .A1(G85), .A2(n653), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U623 ( .A1(G47), .A2(n660), .ZN(n568) );
  NAND2_X1 U624 ( .A1(G60), .A2(n665), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n569) );
  OR2_X1 U626 ( .A1(n570), .A2(n569), .ZN(G290) );
  XOR2_X1 U627 ( .A(G2443), .B(G2446), .Z(n572) );
  XNOR2_X1 U628 ( .A(G2427), .B(G2451), .ZN(n571) );
  XNOR2_X1 U629 ( .A(n572), .B(n571), .ZN(n578) );
  XOR2_X1 U630 ( .A(G2430), .B(G2454), .Z(n574) );
  XNOR2_X1 U631 ( .A(G1341), .B(G1348), .ZN(n573) );
  XNOR2_X1 U632 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U633 ( .A(G2435), .B(G2438), .Z(n575) );
  XNOR2_X1 U634 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U635 ( .A(n578), .B(n577), .Z(n579) );
  AND2_X1 U636 ( .A1(G14), .A2(n579), .ZN(G401) );
  NAND2_X1 U637 ( .A1(G52), .A2(n660), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G64), .A2(n665), .ZN(n580) );
  NAND2_X1 U639 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U640 ( .A1(n652), .A2(G77), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G90), .A2(n653), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n584), .Z(n585) );
  NOR2_X1 U644 ( .A1(n586), .A2(n585), .ZN(G171) );
  AND2_X1 U645 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U646 ( .A(G57), .ZN(G237) );
  INV_X1 U647 ( .A(G132), .ZN(G219) );
  INV_X1 U648 ( .A(G82), .ZN(G220) );
  NAND2_X1 U649 ( .A1(G7), .A2(G661), .ZN(n587) );
  XNOR2_X1 U650 ( .A(n587), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U651 ( .A(G223), .ZN(n842) );
  NAND2_X1 U652 ( .A1(n842), .A2(G567), .ZN(n588) );
  XOR2_X1 U653 ( .A(KEYINPUT11), .B(n588), .Z(G234) );
  NAND2_X1 U654 ( .A1(G81), .A2(n653), .ZN(n589) );
  XNOR2_X1 U655 ( .A(n589), .B(KEYINPUT12), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G68), .A2(n652), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n592), .B(KEYINPUT13), .ZN(n594) );
  NAND2_X1 U659 ( .A1(G43), .A2(n660), .ZN(n593) );
  NAND2_X1 U660 ( .A1(n594), .A2(n593), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G56), .A2(n665), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n595), .B(KEYINPUT14), .ZN(n596) );
  XNOR2_X1 U663 ( .A(n596), .B(KEYINPUT65), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n1003), .A2(G860), .ZN(G153) );
  XOR2_X1 U665 ( .A(G171), .B(KEYINPUT66), .Z(G301) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n608) );
  NAND2_X1 U667 ( .A1(n652), .A2(G79), .ZN(n600) );
  NAND2_X1 U668 ( .A1(G92), .A2(n653), .ZN(n599) );
  NAND2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U670 ( .A1(G54), .A2(n660), .ZN(n602) );
  NAND2_X1 U671 ( .A1(G66), .A2(n665), .ZN(n601) );
  NAND2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n606) );
  XNOR2_X1 U674 ( .A(KEYINPUT67), .B(KEYINPUT15), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n606), .B(n605), .ZN(n914) );
  INV_X1 U676 ( .A(n914), .ZN(n985) );
  INV_X1 U677 ( .A(G868), .ZN(n675) );
  NAND2_X1 U678 ( .A1(n985), .A2(n675), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(G284) );
  XOR2_X1 U680 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U681 ( .A1(G53), .A2(n660), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G65), .A2(n665), .ZN(n609) );
  NAND2_X1 U683 ( .A1(n610), .A2(n609), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n652), .A2(G78), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G91), .A2(n653), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n989) );
  INV_X1 U688 ( .A(n989), .ZN(G299) );
  NAND2_X1 U689 ( .A1(G868), .A2(G286), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G299), .A2(n675), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(G297) );
  INV_X1 U692 ( .A(G860), .ZN(n641) );
  NAND2_X1 U693 ( .A1(n641), .A2(G559), .ZN(n617) );
  NAND2_X1 U694 ( .A1(n617), .A2(n914), .ZN(n618) );
  XNOR2_X1 U695 ( .A(n618), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U696 ( .A1(n1003), .A2(n675), .ZN(n619) );
  XOR2_X1 U697 ( .A(KEYINPUT72), .B(n619), .Z(n622) );
  NAND2_X1 U698 ( .A1(G868), .A2(n914), .ZN(n620) );
  NOR2_X1 U699 ( .A1(G559), .A2(n620), .ZN(n621) );
  NOR2_X1 U700 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U701 ( .A1(n904), .A2(G99), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G135), .A2(n906), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G111), .A2(n898), .ZN(n623) );
  NAND2_X1 U704 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U705 ( .A1(n899), .A2(G123), .ZN(n625) );
  XOR2_X1 U706 ( .A(KEYINPUT18), .B(n625), .Z(n626) );
  NOR2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U709 ( .A(KEYINPUT73), .B(n630), .Z(n930) );
  XOR2_X1 U710 ( .A(G2096), .B(KEYINPUT74), .Z(n631) );
  XNOR2_X1 U711 ( .A(n930), .B(n631), .ZN(n633) );
  INV_X1 U712 ( .A(G2100), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G156) );
  NAND2_X1 U714 ( .A1(G55), .A2(n660), .ZN(n635) );
  NAND2_X1 U715 ( .A1(G67), .A2(n665), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n652), .A2(G80), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G93), .A2(n653), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n676) );
  NAND2_X1 U721 ( .A1(G559), .A2(n914), .ZN(n640) );
  XNOR2_X1 U722 ( .A(n640), .B(n1003), .ZN(n673) );
  NAND2_X1 U723 ( .A1(n641), .A2(n673), .ZN(n642) );
  XNOR2_X1 U724 ( .A(n642), .B(KEYINPUT75), .ZN(n643) );
  XNOR2_X1 U725 ( .A(n676), .B(n643), .ZN(G145) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(KEYINPUT76), .Z(n645) );
  NAND2_X1 U727 ( .A1(G73), .A2(n652), .ZN(n644) );
  XNOR2_X1 U728 ( .A(n645), .B(n644), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n660), .A2(G48), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G86), .A2(n653), .ZN(n646) );
  NAND2_X1 U731 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U732 ( .A1(n649), .A2(n648), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n665), .A2(G61), .ZN(n650) );
  NAND2_X1 U734 ( .A1(n651), .A2(n650), .ZN(G305) );
  NAND2_X1 U735 ( .A1(n652), .A2(G75), .ZN(n655) );
  NAND2_X1 U736 ( .A1(G88), .A2(n653), .ZN(n654) );
  NAND2_X1 U737 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U738 ( .A1(G50), .A2(n660), .ZN(n657) );
  NAND2_X1 U739 ( .A1(G62), .A2(n665), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U741 ( .A1(n659), .A2(n658), .ZN(G166) );
  NAND2_X1 U742 ( .A1(G49), .A2(n660), .ZN(n663) );
  NAND2_X1 U743 ( .A1(G87), .A2(n661), .ZN(n662) );
  NAND2_X1 U744 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U745 ( .A1(n665), .A2(n664), .ZN(n667) );
  NAND2_X1 U746 ( .A1(G651), .A2(G74), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(G288) );
  XNOR2_X1 U748 ( .A(G166), .B(KEYINPUT19), .ZN(n669) );
  XNOR2_X1 U749 ( .A(G290), .B(n989), .ZN(n668) );
  XNOR2_X1 U750 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U751 ( .A(n676), .B(n670), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n671), .B(G288), .ZN(n672) );
  XNOR2_X1 U753 ( .A(G305), .B(n672), .ZN(n918) );
  XNOR2_X1 U754 ( .A(n918), .B(n673), .ZN(n674) );
  NAND2_X1 U755 ( .A1(n674), .A2(G868), .ZN(n678) );
  NAND2_X1 U756 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U758 ( .A(KEYINPUT77), .B(n679), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2078), .A2(G2084), .ZN(n680) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n680), .Z(n681) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n681), .ZN(n682) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U763 ( .A1(n683), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U765 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U766 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U767 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G96), .A2(n686), .ZN(n846) );
  NAND2_X1 U769 ( .A1(n846), .A2(G2106), .ZN(n690) );
  NAND2_X1 U770 ( .A1(G69), .A2(G120), .ZN(n687) );
  NOR2_X1 U771 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U772 ( .A1(G108), .A2(n688), .ZN(n847) );
  NAND2_X1 U773 ( .A1(n847), .A2(G567), .ZN(n689) );
  NAND2_X1 U774 ( .A1(n690), .A2(n689), .ZN(n848) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n691) );
  NOR2_X1 U776 ( .A1(n848), .A2(n691), .ZN(n845) );
  NAND2_X1 U777 ( .A1(n845), .A2(G36), .ZN(G176) );
  XNOR2_X1 U778 ( .A(KEYINPUT79), .B(G166), .ZN(G303) );
  NAND2_X1 U779 ( .A1(G40), .A2(G160), .ZN(n693) );
  XNOR2_X1 U780 ( .A(n693), .B(KEYINPUT81), .ZN(n773) );
  NAND2_X2 U781 ( .A1(n775), .A2(n773), .ZN(n740) );
  NAND2_X1 U782 ( .A1(n740), .A2(G8), .ZN(n762) );
  INV_X1 U783 ( .A(KEYINPUT90), .ZN(n694) );
  XNOR2_X2 U784 ( .A(n740), .B(n694), .ZN(n718) );
  NAND2_X1 U785 ( .A1(n718), .A2(G2072), .ZN(n696) );
  XOR2_X1 U786 ( .A(KEYINPUT91), .B(KEYINPUT27), .Z(n695) );
  XNOR2_X1 U787 ( .A(n696), .B(n695), .ZN(n698) );
  INV_X1 U788 ( .A(G1956), .ZN(n1015) );
  NOR2_X1 U789 ( .A1(n718), .A2(n1015), .ZN(n697) );
  NOR2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n712) );
  NOR2_X1 U791 ( .A1(n989), .A2(n712), .ZN(n699) );
  XOR2_X1 U792 ( .A(G1996), .B(KEYINPUT92), .Z(n956) );
  NOR2_X1 U793 ( .A1(n956), .A2(n740), .ZN(n700) );
  XOR2_X1 U794 ( .A(KEYINPUT26), .B(n700), .Z(n701) );
  NAND2_X1 U795 ( .A1(n1003), .A2(n701), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G1341), .A2(n740), .ZN(n702) );
  XNOR2_X1 U797 ( .A(KEYINPUT93), .B(n702), .ZN(n703) );
  NOR2_X1 U798 ( .A1(n704), .A2(n703), .ZN(n709) );
  NAND2_X1 U799 ( .A1(n914), .A2(n709), .ZN(n708) );
  NAND2_X1 U800 ( .A1(G2067), .A2(n718), .ZN(n706) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n740), .ZN(n705) );
  NAND2_X1 U802 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n711) );
  OR2_X1 U804 ( .A1(n914), .A2(n709), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n989), .A2(n712), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n529), .A2(n715), .ZN(n717) );
  XOR2_X1 U809 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n716) );
  XNOR2_X1 U810 ( .A(n717), .B(n716), .ZN(n722) );
  XNOR2_X1 U811 ( .A(KEYINPUT25), .B(G2078), .ZN(n957) );
  NAND2_X1 U812 ( .A1(n718), .A2(n957), .ZN(n720) );
  INV_X1 U813 ( .A(G1961), .ZN(n1010) );
  NAND2_X1 U814 ( .A1(n1010), .A2(n740), .ZN(n719) );
  NAND2_X1 U815 ( .A1(n720), .A2(n719), .ZN(n723) );
  NAND2_X1 U816 ( .A1(n723), .A2(G171), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n737) );
  NOR2_X1 U818 ( .A1(G171), .A2(n723), .ZN(n724) );
  XNOR2_X1 U819 ( .A(n724), .B(KEYINPUT96), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G1966), .A2(n762), .ZN(n726) );
  NOR2_X1 U821 ( .A1(G2084), .A2(n740), .ZN(n727) );
  XOR2_X1 U822 ( .A(KEYINPUT88), .B(n727), .Z(n749) );
  NAND2_X1 U823 ( .A1(n749), .A2(G8), .ZN(n728) );
  NOR2_X1 U824 ( .A1(n754), .A2(n728), .ZN(n729) );
  XNOR2_X1 U825 ( .A(n729), .B(n527), .ZN(n731) );
  AND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n735) );
  XNOR2_X1 U828 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n752) );
  NAND2_X1 U830 ( .A1(n752), .A2(G286), .ZN(n739) );
  XNOR2_X1 U831 ( .A(n739), .B(n738), .ZN(n745) );
  NOR2_X1 U832 ( .A1(G1971), .A2(n762), .ZN(n742) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U835 ( .A1(G303), .A2(n743), .ZN(n744) );
  NAND2_X1 U836 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n746), .A2(G8), .ZN(n748) );
  XNOR2_X1 U838 ( .A(n748), .B(n747), .ZN(n756) );
  INV_X1 U839 ( .A(n749), .ZN(n750) );
  NAND2_X1 U840 ( .A1(G8), .A2(n750), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n807) );
  INV_X1 U844 ( .A(n807), .ZN(n760) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U846 ( .A1(G8), .A2(n757), .ZN(n758) );
  XOR2_X1 U847 ( .A(KEYINPUT101), .B(n758), .Z(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U849 ( .A1(n762), .A2(n761), .ZN(n766) );
  INV_X1 U850 ( .A(n762), .ZN(n814) );
  NOR2_X1 U851 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XNOR2_X1 U852 ( .A(n763), .B(KEYINPUT24), .ZN(n764) );
  NAND2_X1 U853 ( .A1(n814), .A2(n764), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n772) );
  XNOR2_X1 U855 ( .A(G1981), .B(G305), .ZN(n983) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n769) );
  NOR2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n991) );
  NAND2_X1 U858 ( .A1(n814), .A2(n991), .ZN(n767) );
  NOR2_X1 U859 ( .A1(n769), .A2(n767), .ZN(n768) );
  XOR2_X1 U860 ( .A(n768), .B(KEYINPUT100), .Z(n813) );
  INV_X1 U861 ( .A(n813), .ZN(n770) );
  OR2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  INV_X1 U863 ( .A(n773), .ZN(n774) );
  NOR2_X1 U864 ( .A1(n775), .A2(n774), .ZN(n837) );
  XNOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  XNOR2_X1 U866 ( .A(KEYINPUT83), .B(KEYINPUT36), .ZN(n786) );
  NAND2_X1 U867 ( .A1(G116), .A2(n898), .ZN(n777) );
  NAND2_X1 U868 ( .A1(G128), .A2(n899), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U870 ( .A(KEYINPUT35), .B(n778), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G140), .A2(n906), .ZN(n780) );
  NAND2_X1 U872 ( .A1(G104), .A2(n904), .ZN(n779) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n782) );
  XOR2_X1 U874 ( .A(KEYINPUT82), .B(KEYINPUT34), .Z(n781) );
  XNOR2_X1 U875 ( .A(n782), .B(n781), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U877 ( .A(n786), .B(n785), .ZN(n887) );
  NOR2_X1 U878 ( .A1(n835), .A2(n887), .ZN(n944) );
  NAND2_X1 U879 ( .A1(n837), .A2(n944), .ZN(n833) );
  XOR2_X1 U880 ( .A(KEYINPUT38), .B(KEYINPUT87), .Z(n788) );
  NAND2_X1 U881 ( .A1(G105), .A2(n904), .ZN(n787) );
  XNOR2_X1 U882 ( .A(n788), .B(n787), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G141), .A2(n906), .ZN(n790) );
  NAND2_X1 U884 ( .A1(G129), .A2(n899), .ZN(n789) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n898), .A2(G117), .ZN(n791) );
  XOR2_X1 U887 ( .A(KEYINPUT86), .B(n791), .Z(n792) );
  NOR2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n889) );
  NAND2_X1 U890 ( .A1(n889), .A2(G1996), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G107), .A2(n898), .ZN(n797) );
  NAND2_X1 U892 ( .A1(G119), .A2(n899), .ZN(n796) );
  NAND2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U894 ( .A(KEYINPUT84), .B(n798), .ZN(n801) );
  NAND2_X1 U895 ( .A1(G131), .A2(n906), .ZN(n799) );
  XNOR2_X1 U896 ( .A(KEYINPUT85), .B(n799), .ZN(n800) );
  NOR2_X1 U897 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U898 ( .A1(n904), .A2(G95), .ZN(n802) );
  NAND2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n886) );
  NAND2_X1 U900 ( .A1(n886), .A2(G1991), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n929) );
  NAND2_X1 U902 ( .A1(n929), .A2(n837), .ZN(n827) );
  AND2_X1 U903 ( .A1(n833), .A2(n827), .ZN(n817) );
  NAND2_X1 U904 ( .A1(n806), .A2(n817), .ZN(n822) );
  NOR2_X1 U905 ( .A1(n991), .A2(n807), .ZN(n810) );
  NOR2_X1 U906 ( .A1(G1971), .A2(G303), .ZN(n808) );
  XOR2_X1 U907 ( .A(KEYINPUT98), .B(n808), .Z(n809) );
  NAND2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U909 ( .A1(G1976), .A2(G288), .ZN(n993) );
  NAND2_X1 U910 ( .A1(n811), .A2(n993), .ZN(n812) );
  XNOR2_X1 U911 ( .A(n812), .B(KEYINPUT99), .ZN(n820) );
  AND2_X1 U912 ( .A1(n814), .A2(n813), .ZN(n816) );
  INV_X1 U913 ( .A(n983), .ZN(n815) );
  AND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n818) );
  AND2_X1 U915 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT102), .ZN(n826) );
  XNOR2_X1 U919 ( .A(G1986), .B(KEYINPUT80), .ZN(n824) );
  XNOR2_X1 U920 ( .A(n824), .B(G290), .ZN(n995) );
  NAND2_X1 U921 ( .A1(n995), .A2(n837), .ZN(n825) );
  NAND2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n840) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n889), .ZN(n937) );
  INV_X1 U924 ( .A(n827), .ZN(n830) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U926 ( .A1(G1991), .A2(n886), .ZN(n933) );
  NOR2_X1 U927 ( .A1(n828), .A2(n933), .ZN(n829) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U929 ( .A1(n937), .A2(n831), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n832), .B(KEYINPUT39), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n835), .A2(n887), .ZN(n941) );
  NAND2_X1 U933 ( .A1(n836), .A2(n941), .ZN(n838) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n841), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n842), .ZN(G217) );
  AND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U939 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U940 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U943 ( .A(G120), .ZN(G236) );
  INV_X1 U944 ( .A(G96), .ZN(G221) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  NOR2_X1 U946 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  INV_X1 U948 ( .A(n848), .ZN(G319) );
  XOR2_X1 U949 ( .A(KEYINPUT104), .B(G1976), .Z(n850) );
  XNOR2_X1 U950 ( .A(G1961), .B(G1956), .ZN(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n851), .B(KEYINPUT41), .Z(n853) );
  XNOR2_X1 U953 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U955 ( .A(G1981), .B(G1971), .Z(n855) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1966), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U958 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT105), .B(G2474), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(G229) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2090), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2084), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n862), .B(G2100), .Z(n864) );
  XNOR2_X1 U965 ( .A(G2078), .B(G2072), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U967 ( .A(G2096), .B(KEYINPUT43), .Z(n866) );
  XNOR2_X1 U968 ( .A(G2678), .B(KEYINPUT103), .ZN(n865) );
  XNOR2_X1 U969 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U970 ( .A(n868), .B(n867), .Z(G227) );
  NAND2_X1 U971 ( .A1(G124), .A2(n899), .ZN(n869) );
  XNOR2_X1 U972 ( .A(n869), .B(KEYINPUT106), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G112), .A2(n898), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G136), .A2(n906), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G100), .A2(n904), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U980 ( .A1(G118), .A2(n898), .ZN(n878) );
  NAND2_X1 U981 ( .A1(G130), .A2(n899), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n885) );
  XNOR2_X1 U983 ( .A(KEYINPUT108), .B(KEYINPUT45), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n906), .A2(G142), .ZN(n881) );
  NAND2_X1 U985 ( .A1(n904), .A2(G106), .ZN(n879) );
  XOR2_X1 U986 ( .A(KEYINPUT107), .B(n879), .Z(n880) );
  NAND2_X1 U987 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U988 ( .A(n883), .B(n882), .Z(n884) );
  NOR2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n897) );
  XOR2_X1 U990 ( .A(n887), .B(n886), .Z(n888) );
  XNOR2_X1 U991 ( .A(n930), .B(n888), .ZN(n893) );
  XNOR2_X1 U992 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n891) );
  XNOR2_X1 U993 ( .A(n889), .B(KEYINPUT109), .ZN(n890) );
  XNOR2_X1 U994 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U995 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U996 ( .A(G160), .B(G162), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n912) );
  XNOR2_X1 U999 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(G115), .A2(n898), .ZN(n901) );
  NAND2_X1 U1001 ( .A1(G127), .A2(n899), .ZN(n900) );
  NAND2_X1 U1002 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U1003 ( .A(n903), .B(n902), .ZN(n910) );
  NAND2_X1 U1004 ( .A1(n904), .A2(G103), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n905), .B(KEYINPUT110), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n906), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n946) );
  XNOR2_X1 U1009 ( .A(G164), .B(n946), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n913), .ZN(G395) );
  XOR2_X1 U1012 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n916) );
  XNOR2_X1 U1013 ( .A(G171), .B(n914), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(n917), .B(G286), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(n920), .B(n1003), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G37), .A2(n921), .ZN(G397) );
  NOR2_X1 U1019 ( .A1(G229), .A2(G227), .ZN(n922) );
  XOR2_X1 U1020 ( .A(KEYINPUT49), .B(n922), .Z(n923) );
  NAND2_X1 U1021 ( .A1(G319), .A2(n923), .ZN(n924) );
  NOR2_X1 U1022 ( .A1(G401), .A2(n924), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT114), .B(n925), .ZN(n927) );
  NOR2_X1 U1024 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT115), .B(n928), .Z(G225) );
  INV_X1 U1027 ( .A(G225), .ZN(G308) );
  INV_X1 U1028 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1029 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1043) );
  XNOR2_X1 U1030 ( .A(KEYINPUT52), .B(KEYINPUT117), .ZN(n953) );
  INV_X1 U1031 ( .A(n929), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G160), .B(G2084), .ZN(n931) );
  NAND2_X1 U1033 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1035 ( .A1(n935), .A2(n934), .ZN(n940) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(n938), .B(KEYINPUT51), .ZN(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n942) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(KEYINPUT116), .B(n945), .ZN(n951) );
  XOR2_X1 U1043 ( .A(G2072), .B(n946), .Z(n948) );
  XOR2_X1 U1044 ( .A(G164), .B(G2078), .Z(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(KEYINPUT50), .B(n949), .ZN(n950) );
  NAND2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n953), .B(n952), .ZN(n954) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n978) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n978), .ZN(n955) );
  NAND2_X1 U1051 ( .A1(n955), .A2(G29), .ZN(n1041) );
  XOR2_X1 U1052 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n969) );
  XOR2_X1 U1053 ( .A(n956), .B(G32), .Z(n959) );
  XOR2_X1 U1054 ( .A(n957), .B(G27), .Z(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(G1991), .B(G25), .ZN(n961) );
  XNOR2_X1 U1057 ( .A(G33), .B(G2072), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(G28), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(KEYINPUT118), .B(G2067), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(G26), .B(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(n969), .B(n968), .ZN(n976) );
  XOR2_X1 U1065 ( .A(KEYINPUT120), .B(G34), .Z(n971) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(n971), .B(n970), .ZN(n972) );
  XNOR2_X1 U1068 ( .A(G2084), .B(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G2090), .B(G35), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n978), .B(n977), .ZN(n980) );
  INV_X1 U1073 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1075 ( .A1(G11), .A2(n981), .ZN(n1039) );
  XNOR2_X1 U1076 ( .A(G16), .B(KEYINPUT56), .ZN(n1009) );
  XOR2_X1 U1077 ( .A(G168), .B(G1966), .Z(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n984), .Z(n1007) );
  XOR2_X1 U1080 ( .A(G171), .B(G1961), .Z(n987) );
  XNOR2_X1 U1081 ( .A(n985), .B(G1348), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1083 ( .A(KEYINPUT122), .B(n988), .ZN(n1002) );
  XNOR2_X1 U1084 ( .A(n1015), .B(n989), .ZN(n990) );
  XNOR2_X1 U1085 ( .A(n990), .B(KEYINPUT123), .ZN(n997) );
  INV_X1 U1086 ( .A(n991), .ZN(n992) );
  NAND2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G1971), .B(G303), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(KEYINPUT124), .B(n998), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(n1003), .B(G1341), .Z(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1037) );
  INV_X1 U1098 ( .A(G16), .ZN(n1035) );
  XNOR2_X1 U1099 ( .A(G5), .B(n1010), .ZN(n1025) );
  XOR2_X1 U1100 ( .A(G1341), .B(G19), .Z(n1011) );
  XNOR2_X1 U1101 ( .A(KEYINPUT125), .B(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G6), .B(G1981), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT126), .B(n1014), .ZN(n1017) );
  XNOR2_X1 U1105 ( .A(n1015), .B(G20), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(KEYINPUT59), .B(G1348), .Z(n1018) );
  XNOR2_X1 U1108 ( .A(G4), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1110 ( .A(KEYINPUT60), .B(n1021), .Z(n1023) );
  XNOR2_X1 U1111 ( .A(G1966), .B(G21), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1113 ( .A1(n1025), .A2(n1024), .ZN(n1032) );
  XNOR2_X1 U1114 ( .A(G1971), .B(G22), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(G23), .B(G1976), .ZN(n1026) );
  NOR2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(G1986), .B(G24), .Z(n1028) );
  NAND2_X1 U1118 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1119 ( .A(KEYINPUT58), .B(n1030), .ZN(n1031) );
  NOR2_X1 U1120 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1121 ( .A(KEYINPUT61), .B(n1033), .ZN(n1034) );
  NAND2_X1 U1122 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1123 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  NOR2_X1 U1124 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  NAND2_X1 U1125 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XNOR2_X1 U1126 ( .A(n1043), .B(n1042), .ZN(G311) );
  INV_X1 U1127 ( .A(G311), .ZN(G150) );
endmodule

