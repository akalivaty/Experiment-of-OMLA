//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n206));
  AND2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  XOR2_X1   g0009(.A(KEYINPUT66), .B(G77), .Z(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  OAI221_X1 g0012(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT65), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n204), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  NOR2_X1   g0017(.A1(new_n204), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AND2_X1   g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(G58), .A2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n224), .A2(G50), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n217), .B(new_n220), .C1(new_n222), .C2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n230), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND2_X1  g0047(.A1(G1), .A2(G13), .ZN(new_n248));
  OAI21_X1  g0048(.A(KEYINPUT68), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n221), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n246), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G238), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G97), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n232), .A2(G1698), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(G226), .B2(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n255), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n247), .A2(new_n248), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n247), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n250), .B1(new_n221), .B2(new_n251), .ZN(new_n267));
  OAI211_X1 g0067(.A(G274), .B(new_n246), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(new_n249), .B2(new_n252), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT69), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(new_n272), .A3(new_n246), .ZN(new_n273));
  AND3_X1   g0073(.A1(new_n269), .A2(KEYINPUT75), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT75), .B1(new_n269), .B2(new_n273), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n254), .B(new_n265), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(KEYINPUT13), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT75), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n268), .A2(KEYINPUT69), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n271), .B2(new_n246), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n278), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n269), .A2(KEYINPUT75), .A3(new_n273), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n283), .A2(new_n284), .A3(new_n254), .A4(new_n265), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n277), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G169), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n286), .A2(new_n289), .A3(G169), .ZN(new_n290));
  INV_X1    g0090(.A(G179), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n288), .B(new_n290), .C1(new_n291), .C2(new_n286), .ZN(new_n292));
  NAND3_X1  g0092(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n248), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n260), .A2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G77), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G50), .ZN(new_n301));
  INV_X1    g0101(.A(G20), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n300), .A2(new_n301), .B1(new_n302), .B2(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n294), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT11), .ZN(new_n305));
  INV_X1    g0105(.A(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OR3_X1    g0110(.A1(new_n310), .A2(KEYINPUT12), .A3(G68), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT12), .B1(new_n310), .B2(G68), .ZN(new_n312));
  INV_X1    g0112(.A(new_n307), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n313), .A2(new_n294), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n311), .A2(new_n312), .B1(G68), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n305), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n292), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n286), .A2(G200), .ZN(new_n318));
  INV_X1    g0118(.A(new_n316), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n286), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n269), .A2(new_n273), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT3), .B(G33), .ZN(new_n323));
  NAND2_X1  g0123(.A1(G238), .A2(G1698), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n323), .B(new_n324), .C1(new_n232), .C2(G1698), .ZN(new_n325));
  OAI211_X1 g0125(.A(new_n325), .B(new_n264), .C1(G107), .C2(new_n323), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n253), .A2(G244), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n291), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n314), .A2(G77), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT73), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT8), .B(G58), .ZN(new_n333));
  OAI22_X1  g0133(.A1(new_n211), .A2(new_n302), .B1(new_n300), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT15), .B(G87), .Z(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n296), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n294), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n332), .B(new_n338), .C1(new_n210), .C2(new_n310), .ZN(new_n339));
  INV_X1    g0139(.A(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n328), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n330), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n317), .A2(new_n321), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G1698), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G222), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G223), .A2(G1698), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n323), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n347), .B(new_n264), .C1(new_n210), .C2(new_n323), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n253), .A2(G226), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n322), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n350), .A2(new_n320), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(G200), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT10), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OR3_X1    g0155(.A1(new_n313), .A2(KEYINPUT71), .A3(new_n301), .ZN(new_n356));
  INV_X1    g0156(.A(new_n294), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT71), .B1(new_n313), .B2(new_n301), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n310), .A4(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n224), .B2(G50), .ZN(new_n360));
  INV_X1    g0160(.A(G150), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n300), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT70), .ZN(new_n363));
  XNOR2_X1  g0163(.A(new_n333), .B(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n362), .B1(new_n364), .B2(new_n295), .ZN(new_n365));
  OAI221_X1 g0165(.A(new_n359), .B1(G50), .B2(new_n310), .C1(new_n365), .C2(new_n357), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT9), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n367), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n368), .A2(new_n352), .A3(new_n351), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n368), .A2(new_n369), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n353), .C1(new_n354), .C2(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n350), .A2(new_n340), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n374), .A2(new_n366), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT72), .B1(new_n350), .B2(G179), .ZN(new_n376));
  OR3_X1    g0176(.A1(new_n350), .A2(KEYINPUT72), .A3(G179), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n371), .A2(new_n373), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT76), .B1(new_n258), .B2(G33), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n260), .A3(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n302), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(KEYINPUT77), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n384), .B2(G20), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n387), .A2(G68), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G58), .ZN(new_n392));
  INV_X1    g0192(.A(G68), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(new_n223), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n299), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n391), .A2(KEYINPUT16), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(new_n396), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n388), .B1(new_n323), .B2(G20), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n258), .A2(G33), .ZN(new_n401));
  OAI211_X1 g0201(.A(KEYINPUT7), .B(new_n302), .C1(new_n380), .C2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n393), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n398), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n397), .A2(new_n404), .A3(new_n294), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT78), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n333), .B(KEYINPUT70), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n407), .A2(new_n314), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n364), .A2(new_n309), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n310), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n411), .B(KEYINPUT78), .C1(new_n407), .C2(new_n314), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n405), .A2(new_n413), .ZN(new_n414));
  OR2_X1    g0214(.A1(G223), .A2(G1698), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n344), .A2(G226), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n384), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(G33), .A2(G87), .ZN(new_n418));
  XOR2_X1   g0218(.A(new_n418), .B(KEYINPUT79), .Z(new_n419));
  OAI21_X1  g0219(.A(new_n264), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n253), .A2(G232), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n322), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT80), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n269), .A2(new_n273), .B1(G232), .B2(new_n253), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT80), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n425), .A3(new_n420), .ZN(new_n426));
  AOI21_X1  g0226(.A(G200), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n422), .A2(G190), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n414), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n414), .B(KEYINPUT17), .C1(new_n427), .C2(new_n428), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n422), .A2(G179), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n423), .A2(new_n426), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n433), .B1(new_n434), .B2(new_n340), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n405), .A2(new_n413), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT18), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n424), .A2(new_n425), .A3(new_n420), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n425), .B1(new_n424), .B2(new_n420), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n340), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n433), .ZN(new_n441));
  AND4_X1   g0241(.A1(KEYINPUT18), .A2(new_n440), .A3(new_n436), .A4(new_n441), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n431), .B(new_n432), .C1(new_n437), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n339), .B1(new_n329), .B2(G190), .ZN(new_n445));
  INV_X1    g0245(.A(G200), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(new_n329), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n379), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n343), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n381), .A2(new_n383), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT22), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n452), .A2(new_n208), .A3(G20), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n451), .A2(new_n259), .A3(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n259), .A2(new_n261), .A3(new_n302), .A4(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(new_n452), .ZN(new_n456));
  INV_X1    g0256(.A(G107), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n302), .A2(G33), .A3(G116), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n454), .A2(new_n456), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT24), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n384), .A2(new_n453), .B1(new_n455), .B2(new_n452), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT24), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n464), .A2(new_n465), .A3(new_n460), .A4(new_n461), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n294), .ZN(new_n468));
  AOI211_X1 g0268(.A(new_n294), .B(new_n309), .C1(new_n306), .C2(G33), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G107), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n309), .A2(new_n457), .ZN(new_n471));
  XOR2_X1   g0271(.A(new_n471), .B(KEYINPUT25), .Z(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n209), .A2(new_n344), .ZN(new_n474));
  INV_X1    g0274(.A(G257), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G1698), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n384), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n264), .ZN(new_n480));
  AND2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  NOR2_X1   g0281(.A1(KEYINPUT5), .A2(G41), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n306), .B(G45), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n271), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n249), .A2(new_n252), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(G264), .A3(new_n483), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n480), .A2(G179), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n264), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n477), .B2(new_n478), .ZN(new_n490));
  INV_X1    g0290(.A(new_n485), .ZN(new_n491));
  INV_X1    g0291(.A(new_n487), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n488), .B(KEYINPUT91), .C1(new_n493), .C2(new_n340), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT91), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n495), .A3(G179), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n473), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n490), .A2(new_n492), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n485), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G200), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n467), .A2(new_n294), .B1(G107), .B2(new_n469), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n493), .A2(G190), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(new_n472), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT92), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT92), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n497), .A2(new_n506), .A3(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n475), .A2(new_n344), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n384), .B(new_n509), .C1(G264), .C2(new_n344), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT88), .B(G303), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n262), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n264), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n486), .A2(G270), .A3(new_n483), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n485), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n291), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(G20), .ZN(new_n522));
  AOI21_X1  g0322(.A(G20), .B1(G33), .B2(G283), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n260), .A2(G97), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT89), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT89), .B1(new_n523), .B2(new_n524), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n294), .B(new_n522), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  INV_X1    g0330(.A(G97), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n530), .B(new_n302), .C1(G33), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT89), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n523), .A2(new_n524), .A3(KEYINPUT89), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(KEYINPUT20), .A3(new_n294), .A4(new_n522), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n309), .A2(new_n521), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n469), .A2(G116), .ZN(new_n540));
  AND4_X1   g0340(.A1(KEYINPUT90), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n529), .A2(new_n537), .B1(new_n469), .B2(G116), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT90), .B1(new_n542), .B2(new_n539), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n520), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n517), .B1(new_n264), .B2(new_n514), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n340), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n541), .B2(new_n543), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT21), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(KEYINPUT21), .B(new_n546), .C1(new_n541), .C2(new_n543), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n519), .A2(new_n320), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n545), .A2(new_n446), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n541), .A2(new_n543), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AND4_X1   g0355(.A1(new_n544), .A2(new_n549), .A3(new_n550), .A4(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n393), .A2(G20), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n451), .A2(new_n259), .A3(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n208), .A2(new_n531), .A3(new_n457), .ZN(new_n561));
  AND2_X1   g0361(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n562));
  NOR2_X1   g0362(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n563));
  NOR3_X1   g0363(.A1(new_n562), .A2(new_n563), .A3(new_n255), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n561), .B1(new_n564), .B2(G20), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n296), .A2(new_n531), .B1(new_n562), .B2(new_n563), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n384), .A2(KEYINPUT86), .A3(new_n557), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n294), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n336), .A2(new_n309), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n469), .A2(new_n335), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n306), .A2(G45), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n209), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n486), .B(new_n574), .C1(G274), .C2(new_n573), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G238), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n212), .B2(G1698), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n384), .A2(new_n577), .B1(G33), .B2(G116), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n575), .B1(new_n578), .B2(new_n489), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n340), .ZN(new_n580));
  INV_X1    g0380(.A(new_n579), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n291), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n572), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n568), .A2(new_n294), .B1(new_n309), .B2(new_n336), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n575), .B(G190), .C1(new_n489), .C2(new_n578), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n469), .A2(G87), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n579), .A2(G200), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT87), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n583), .A2(KEYINPUT87), .A3(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n310), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n469), .B2(G97), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n400), .A2(new_n402), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n597), .B2(G107), .ZN(new_n598));
  AOI211_X1 g0398(.A(KEYINPUT81), .B(new_n457), .C1(new_n400), .C2(new_n402), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT6), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n600), .A2(new_n531), .A3(G107), .ZN(new_n601));
  XNOR2_X1  g0401(.A(G97), .B(G107), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n302), .B1(new_n297), .B2(new_n300), .ZN(new_n604));
  NOR3_X1   g0404(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n595), .B1(new_n605), .B2(new_n357), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT82), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT4), .B1(new_n384), .B2(G244), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT4), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n609), .A2(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n610), .A2(new_n259), .A3(new_n261), .A4(G244), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n530), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n259), .A2(new_n261), .A3(G250), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n344), .B1(new_n613), .B2(KEYINPUT4), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n608), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n607), .B1(new_n615), .B2(new_n489), .ZN(new_n616));
  OAI211_X1 g0416(.A(G257), .B(new_n483), .C1(new_n266), .C2(new_n267), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT83), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT83), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n486), .A2(new_n619), .A3(G257), .A4(new_n483), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n618), .A2(new_n485), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n451), .A2(G244), .A3(new_n259), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n609), .ZN(new_n623));
  INV_X1    g0423(.A(new_n614), .ZN(new_n624));
  INV_X1    g0424(.A(new_n612), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(KEYINPUT82), .A3(new_n264), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n616), .A2(new_n291), .A3(new_n621), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n264), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n340), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n606), .A2(new_n628), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT84), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n323), .A2(new_n388), .A3(G20), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT7), .B1(new_n262), .B2(new_n302), .ZN(new_n636));
  OAI21_X1  g0436(.A(G107), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT81), .ZN(new_n638));
  INV_X1    g0438(.A(new_n604), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n597), .A2(new_n596), .A3(G107), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n638), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(new_n294), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n642), .A2(new_n595), .B1(new_n630), .B2(new_n340), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(KEYINPUT84), .A3(new_n628), .ZN(new_n644));
  INV_X1    g0444(.A(new_n606), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n616), .A2(new_n621), .A3(new_n627), .ZN(new_n646));
  INV_X1    g0446(.A(new_n630), .ZN(new_n647));
  AOI22_X1  g0447(.A1(G200), .A2(new_n646), .B1(new_n647), .B2(G190), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n634), .A2(new_n644), .B1(new_n645), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n508), .A2(new_n556), .A3(new_n593), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n450), .A2(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n378), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n437), .A2(new_n442), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n342), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n292), .A2(new_n316), .B1(new_n321), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n431), .A2(new_n432), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n371), .A2(new_n373), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT93), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT84), .B1(new_n643), .B2(new_n628), .ZN(new_n663));
  AND4_X1   g0463(.A1(KEYINPUT84), .A2(new_n606), .A3(new_n628), .A4(new_n631), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n662), .B1(new_n665), .B2(new_n593), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n589), .A2(new_n632), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n583), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n661), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n503), .A2(new_n583), .A3(new_n588), .ZN(new_n670));
  INV_X1    g0470(.A(new_n497), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n549), .A2(new_n544), .A3(new_n550), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n649), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n592), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT87), .B1(new_n583), .B2(new_n588), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n634), .B(new_n644), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(new_n583), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n589), .A2(new_n632), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n678), .B1(new_n679), .B2(new_n662), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(KEYINPUT93), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n669), .A2(new_n673), .A3(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n660), .B1(new_n450), .B2(new_n683), .ZN(G369));
  INV_X1    g0484(.A(KEYINPUT94), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n308), .A2(G20), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(new_n221), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT27), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n685), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G213), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  OAI211_X1 g0492(.A(KEYINPUT94), .B(KEYINPUT27), .C1(new_n687), .C2(new_n221), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n554), .A2(new_n697), .ZN(new_n698));
  MUX2_X1   g0498(.A(new_n556), .B(new_n672), .S(new_n698), .Z(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n508), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n697), .B1(new_n501), .B2(new_n472), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n702), .A2(new_n703), .B1(new_n497), .B2(new_n697), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n671), .A2(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n672), .A2(new_n697), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n508), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n705), .A2(new_n706), .A3(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n218), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n561), .A2(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n225), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n665), .A2(new_n662), .A3(new_n593), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n667), .A2(KEYINPUT26), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n673), .A2(new_n718), .A3(new_n583), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n697), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n682), .A2(new_n697), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(KEYINPUT29), .ZN(new_n724));
  AND4_X1   g0524(.A1(new_n498), .A2(new_n520), .A3(new_n647), .A4(new_n581), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT30), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n545), .A2(new_n581), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n646), .A2(new_n728), .A3(new_n291), .A4(new_n499), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n696), .ZN(new_n731));
  OAI211_X1 g0531(.A(KEYINPUT31), .B(new_n731), .C1(new_n650), .C2(new_n696), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n731), .A2(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n724), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n717), .B1(new_n737), .B2(G1), .ZN(G364));
  OR2_X1    g0538(.A1(new_n699), .A2(G330), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n306), .B1(new_n686), .B2(G45), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n712), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n739), .A2(new_n700), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n320), .A2(G20), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n446), .A2(G179), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G283), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n302), .A2(new_n320), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n747), .ZN(new_n753));
  INV_X1    g0553(.A(G303), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n291), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  OAI221_X1 g0557(.A(new_n262), .B1(new_n753), .B2(new_n754), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n291), .A2(new_n446), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n746), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n746), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n752), .A2(new_n755), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(G329), .B1(new_n768), .B2(G322), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n751), .A2(new_n763), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n302), .B1(new_n764), .B2(G190), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G326), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n759), .A2(new_n752), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n770), .B1(new_n771), .B2(new_n775), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n749), .A2(new_n457), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(G68), .B2(new_n761), .ZN(new_n780));
  INV_X1    g0580(.A(new_n753), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G87), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n775), .A2(new_n531), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n211), .A2(new_n756), .B1(new_n301), .B2(new_n777), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(G58), .B2(new_n768), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(new_n785), .B2(KEYINPUT96), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n766), .A2(G159), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT32), .Z(new_n788));
  NAND4_X1  g0588(.A1(new_n780), .A2(new_n782), .A3(new_n786), .A4(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n323), .B1(new_n785), .B2(KEYINPUT96), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n778), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n248), .B1(G20), .B2(new_n340), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G13), .A2(G33), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(G20), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n793), .B1(new_n699), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n218), .A2(G355), .A3(new_n323), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n711), .A2(new_n384), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G45), .B2(new_n225), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n239), .A2(new_n245), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n799), .B1(G116), .B2(new_n218), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(new_n792), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n743), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT95), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n744), .B1(new_n798), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT99), .ZN(G396));
  NOR2_X1   g0608(.A1(new_n342), .A2(new_n696), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n339), .A2(new_n696), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n447), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n809), .B1(new_n811), .B2(new_n342), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n723), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n682), .A2(new_n697), .A3(new_n812), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(new_n736), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n743), .ZN(new_n818));
  INV_X1    g0618(.A(new_n792), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n262), .B1(new_n777), .B2(new_n754), .C1(new_n521), .C2(new_n756), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n749), .A2(new_n208), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n783), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n771), .B2(new_n767), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(G311), .C2(new_n766), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n457), .B2(new_n753), .C1(new_n825), .C2(new_n760), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n761), .A2(G150), .B1(new_n768), .B2(G143), .ZN(new_n827));
  INV_X1    g0627(.A(new_n777), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G137), .ZN(new_n829));
  INV_X1    g0629(.A(G159), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n827), .B(new_n829), .C1(new_n830), .C2(new_n756), .ZN(new_n831));
  XOR2_X1   g0631(.A(KEYINPUT100), .B(KEYINPUT34), .Z(new_n832));
  XNOR2_X1  g0632(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n384), .B1(new_n301), .B2(new_n753), .C1(new_n775), .C2(new_n392), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(G68), .B2(new_n750), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n833), .B(new_n835), .C1(new_n836), .C2(new_n765), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n819), .B1(new_n826), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n792), .A2(new_n794), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n743), .B(new_n838), .C1(new_n297), .C2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n795), .B2(new_n812), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n818), .A2(new_n841), .ZN(G384));
  NOR2_X1   g0642(.A1(new_n319), .A2(new_n697), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n289), .B1(new_n286), .B2(G169), .ZN(new_n845));
  AOI211_X1 g0645(.A(KEYINPUT14), .B(new_n340), .C1(new_n277), .C2(new_n285), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n286), .A2(new_n291), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n321), .B(new_n844), .C1(new_n848), .C2(new_n319), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT102), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n848), .B2(new_n844), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n292), .A2(KEYINPUT102), .A3(new_n843), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n397), .A2(new_n294), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n391), .B2(new_n396), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n854), .A2(new_n855), .B1(new_n409), .B2(new_n408), .ZN(new_n856));
  INV_X1    g0656(.A(new_n694), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n443), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n440), .A2(new_n436), .A3(new_n441), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n436), .A2(new_n857), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n429), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n440), .A2(new_n856), .A3(new_n441), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n429), .A2(new_n865), .A3(new_n858), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n864), .B1(new_n866), .B2(new_n862), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT38), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n809), .B(KEYINPUT101), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI221_X4 g0673(.A(new_n853), .B1(new_n870), .B2(new_n871), .C1(new_n815), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n654), .A2(new_n857), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT103), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n860), .A2(KEYINPUT38), .A3(new_n867), .ZN(new_n877));
  AOI21_X1  g0677(.A(KEYINPUT38), .B1(new_n860), .B2(new_n867), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT39), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT39), .ZN(new_n881));
  INV_X1    g0681(.A(new_n863), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n443), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n429), .A2(new_n861), .A3(new_n863), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n864), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n881), .B1(new_n877), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n880), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n317), .A2(new_n696), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n815), .A2(new_n873), .ZN(new_n893));
  INV_X1    g0693(.A(new_n879), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT103), .ZN(new_n897));
  INV_X1    g0697(.A(new_n875), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n876), .A2(new_n892), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n724), .A2(new_n449), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n660), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n895), .A2(new_n732), .A3(new_n733), .A4(new_n812), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n877), .B2(new_n887), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n443), .A2(new_n882), .B1(new_n885), .B2(new_n864), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n871), .B(KEYINPUT104), .C1(KEYINPUT38), .C2(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n905), .A2(KEYINPUT40), .A3(new_n907), .A4(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT40), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n904), .B2(new_n879), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n734), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n449), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n916), .A2(new_n735), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n903), .B(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n306), .B2(new_n686), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT35), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n222), .B1(new_n603), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n921), .B(G116), .C1(new_n920), .C2(new_n603), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT36), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n225), .A2(new_n394), .ZN(new_n924));
  OAI22_X1  g0724(.A1(new_n924), .A2(new_n211), .B1(G50), .B2(new_n393), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(G1), .A3(new_n308), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n923), .A3(new_n926), .ZN(G367));
  OAI21_X1  g0727(.A(new_n649), .B1(new_n645), .B2(new_n697), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n643), .A2(new_n628), .A3(new_n696), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n705), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n584), .A2(new_n586), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n696), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n583), .A3(new_n588), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n583), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT105), .Z(new_n938));
  NAND3_X1  g0738(.A1(new_n708), .A2(new_n508), .A3(new_n649), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT42), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n665), .B1(new_n930), .B2(new_n671), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n941), .A2(new_n696), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n938), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n932), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n932), .B1(new_n943), .B2(new_n945), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n944), .A2(KEYINPUT106), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n712), .B(KEYINPUT41), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n709), .A2(new_n706), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n931), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT44), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n955), .A2(new_n931), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n705), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n704), .A2(new_n708), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(KEYINPUT107), .B2(new_n709), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(KEYINPUT107), .B2(new_n709), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n701), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n737), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n954), .B1(new_n968), .B2(new_n737), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n952), .B1(new_n969), .B2(new_n741), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n230), .A2(new_n711), .A3(new_n384), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n804), .B1(new_n218), .B2(new_n336), .ZN(new_n972));
  INV_X1    g0772(.A(G143), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n760), .A2(new_n830), .B1(new_n777), .B2(new_n973), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n323), .B1(new_n392), .B2(new_n753), .C1(new_n211), .C2(new_n748), .ZN(new_n975));
  INV_X1    g0775(.A(new_n756), .ZN(new_n976));
  AOI211_X1 g0776(.A(new_n974), .B(new_n975), .C1(G50), .C2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n775), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(G68), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n768), .A2(G150), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n766), .A2(G137), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n977), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n976), .A2(G283), .B1(new_n761), .B2(G294), .ZN(new_n983));
  INV_X1    g0783(.A(G317), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n531), .B2(new_n748), .C1(new_n984), .C2(new_n765), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n512), .B2(new_n768), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n781), .A2(G116), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT46), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n384), .B1(new_n828), .B2(G311), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n775), .A2(new_n457), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n982), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n992), .B(KEYINPUT47), .Z(new_n993));
  OAI221_X1 g0793(.A(new_n742), .B1(new_n971), .B2(new_n972), .C1(new_n993), .C2(new_n819), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT108), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n797), .B2(new_n936), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n970), .A2(new_n996), .ZN(G387));
  OR2_X1    g0797(.A1(new_n966), .A2(new_n737), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n998), .A2(new_n712), .A3(new_n967), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n235), .A2(G45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT109), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n333), .A2(G50), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT110), .Z(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  AOI21_X1  g0804(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n714), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n800), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n218), .A2(new_n323), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1007), .B1(G107), .B2(new_n218), .C1(new_n714), .C2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n804), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n742), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n704), .A2(new_n797), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n384), .B1(new_n407), .B2(new_n760), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n978), .A2(new_n335), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(G159), .A2(new_n828), .B1(new_n781), .B2(new_n210), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1014), .B(new_n1015), .C1(new_n393), .C2(new_n756), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(G150), .C2(new_n766), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n301), .B2(new_n767), .C1(new_n531), .C2(new_n749), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n761), .A2(G311), .B1(new_n768), .B2(G317), .ZN(new_n1019));
  INV_X1    g0819(.A(G322), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n777), .C1(new_n511), .C2(new_n756), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT48), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n825), .B2(new_n775), .C1(new_n771), .C2(new_n753), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n385), .B1(new_n748), .B2(new_n521), .C1(new_n776), .C2(new_n765), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1018), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1011), .B(new_n1012), .C1(new_n792), .C2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n966), .B2(new_n741), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n999), .A2(new_n1029), .ZN(G393));
  NAND2_X1  g0830(.A1(new_n962), .A2(new_n967), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n968), .A2(new_n712), .A3(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n962), .A2(new_n740), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n978), .A2(G116), .B1(new_n512), .B2(new_n761), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT113), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n771), .C2(new_n756), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT114), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n777), .A2(new_n984), .B1(new_n767), .B2(new_n757), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT52), .Z(new_n1041));
  OAI21_X1  g0841(.A(new_n262), .B1(new_n753), .B2(new_n825), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1041), .A2(new_n779), .A3(new_n1042), .ZN(new_n1043));
  OAI211_X1 g0843(.A(new_n1039), .B(new_n1043), .C1(new_n1020), .C2(new_n765), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(G150), .A2(new_n828), .B1(new_n768), .B2(G159), .ZN(new_n1045));
  AND2_X1   g0845(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(KEYINPUT51), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n753), .A2(new_n393), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1046), .A2(new_n821), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n978), .A2(G77), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n766), .A2(G143), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n384), .B1(new_n756), .B2(new_n333), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(G50), .B2(new_n761), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n819), .B1(new_n1044), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n804), .B1(new_n218), .B2(new_n531), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n800), .B2(new_n242), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1055), .A2(new_n743), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n931), .A2(new_n796), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT112), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1033), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1032), .A2(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(G390));
  NAND2_X1  g0865(.A1(new_n893), .A2(new_n895), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n891), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(KEYINPUT116), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT116), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n853), .B1(new_n815), .B2(new_n873), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1069), .B1(new_n1070), .B2(new_n891), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1068), .A2(new_n889), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n720), .A2(new_n697), .A3(new_n812), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n873), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n891), .B1(new_n1074), .B2(new_n895), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n907), .A3(new_n909), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1072), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n732), .A2(new_n733), .A3(G330), .A4(new_n812), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n853), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n1078), .A2(new_n853), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1072), .A2(new_n1076), .A3(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n741), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n890), .A2(new_n795), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1050), .B1(new_n393), .B2(new_n749), .C1(new_n771), .C2(new_n765), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n777), .A2(new_n825), .ZN(new_n1087));
  NOR2_X1   g0887(.A1(new_n767), .A2(new_n521), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n976), .A2(G97), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n761), .A2(G107), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1089), .A2(new_n1090), .A3(new_n262), .A4(new_n782), .ZN(new_n1091));
  NOR4_X1   g0891(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n323), .B1(new_n748), .B2(new_n301), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT117), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1093), .A2(new_n1094), .B1(G137), .B2(new_n761), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT54), .B(G143), .Z(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .C1(new_n756), .C2(new_n1097), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n753), .A2(KEYINPUT53), .A3(new_n361), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n765), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G128), .A2(new_n828), .B1(new_n768), .B2(G132), .ZN(new_n1102));
  OAI21_X1  g0902(.A(KEYINPUT53), .B1(new_n753), .B2(new_n361), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n775), .C2(new_n830), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n792), .B1(new_n1092), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n407), .A2(new_n839), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n742), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1084), .B1(new_n1085), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1078), .A2(new_n853), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1081), .A2(new_n873), .A3(new_n1073), .A4(new_n1110), .ZN(new_n1111));
  AND2_X1   g0911(.A1(new_n1078), .A2(new_n853), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n893), .B1(new_n1112), .B2(new_n1079), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n914), .A2(G330), .A3(new_n449), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n901), .A2(new_n660), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1083), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1080), .A2(new_n1119), .A3(new_n1082), .ZN(new_n1121));
  AND2_X1   g0921(.A1(new_n1121), .A2(new_n712), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1109), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(G378));
  NAND2_X1  g0924(.A1(new_n1121), .A2(new_n1117), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n907), .A2(KEYINPUT40), .A3(new_n909), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n912), .B(G330), .C1(new_n1126), .C2(new_n904), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n379), .B(new_n1128), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n366), .A2(new_n857), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1129), .B(new_n1130), .Z(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n910), .A2(new_n1131), .A3(G330), .A4(new_n912), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI211_X1 g0935(.A(KEYINPUT103), .B(new_n875), .C1(new_n1070), .C2(new_n894), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n897), .B1(new_n896), .B2(new_n898), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1135), .A2(new_n892), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n900), .A2(new_n1134), .A3(new_n1133), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT121), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1139), .A2(new_n1140), .A3(KEYINPUT121), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1125), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT57), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1139), .A2(KEYINPUT123), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1139), .A2(new_n1140), .A3(KEYINPUT123), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1125), .A2(KEYINPUT57), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n712), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1143), .A2(new_n741), .A3(new_n1144), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n777), .A2(new_n521), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n761), .A2(G97), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n976), .A2(new_n335), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n979), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1156), .B(new_n244), .C1(new_n392), .C2(new_n748), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(G107), .C2(new_n768), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n384), .B1(new_n781), .B2(new_n210), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n825), .C2(new_n765), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G41), .B1(new_n384), .B2(G33), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n775), .A2(new_n361), .B1(new_n1100), .B2(new_n777), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n768), .A2(G128), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n753), .C2(new_n1097), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G137), .B2(new_n976), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n836), .B2(new_n760), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(G41), .B1(new_n766), .B2(G124), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n1171), .B(new_n260), .C1(new_n830), .C2(new_n748), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1161), .B1(G50), .B2(new_n1162), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT120), .Z(new_n1174));
  AOI21_X1  g0974(.A(new_n743), .B1(new_n1174), .B2(new_n792), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n839), .A2(new_n301), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n1175), .B(new_n1176), .C1(new_n795), .C2(new_n1132), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT122), .B1(new_n1152), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1152), .A2(KEYINPUT122), .A3(new_n1177), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1151), .B1(new_n1178), .B2(new_n1180), .ZN(G375));
  NAND3_X1  g0981(.A1(new_n1116), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1118), .A2(new_n953), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n853), .A2(new_n794), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1014), .B1(new_n521), .B2(new_n760), .C1(new_n825), .C2(new_n767), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G77), .B2(new_n750), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n754), .B2(new_n765), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n323), .B(new_n1187), .C1(G97), .C2(new_n781), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n457), .B2(new_n756), .C1(new_n771), .C2(new_n777), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n775), .A2(new_n301), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n976), .A2(G150), .B1(new_n781), .B2(G159), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n392), .B2(new_n748), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(G137), .C2(new_n768), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n766), .A2(G128), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n761), .A2(new_n1096), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n385), .B1(G132), .B2(new_n828), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n819), .B1(new_n1189), .B2(new_n1197), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n743), .B(new_n1198), .C1(new_n393), .C2(new_n839), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n1114), .A2(new_n741), .B1(new_n1184), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1183), .A2(new_n1200), .ZN(G381));
  NAND2_X1  g1001(.A1(new_n1152), .A2(new_n1177), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT122), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n713), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1204), .A2(new_n1179), .B1(new_n1205), .B2(new_n1150), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1123), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1063), .A2(new_n970), .A3(new_n996), .A4(new_n1064), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n1200), .A3(new_n1183), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1209), .A2(G396), .A3(G393), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1208), .A2(new_n1212), .ZN(G407));
  OAI21_X1  g1013(.A(new_n1208), .B1(new_n1212), .B2(new_n695), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(G213), .ZN(G409));
  NOR2_X1   g1015(.A1(new_n691), .A2(G343), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1145), .A2(new_n954), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1148), .A2(new_n741), .A3(new_n1149), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1123), .A2(new_n1218), .A3(new_n1177), .A4(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1217), .B(new_n1220), .C1(new_n1206), .C2(new_n1123), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT125), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT60), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1182), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(new_n1118), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(KEYINPUT124), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1116), .A2(new_n1111), .A3(new_n1113), .A4(KEYINPUT60), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n712), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT124), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1224), .A2(new_n1230), .A3(new_n1118), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1229), .A3(new_n1231), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1232), .A2(G384), .A3(new_n1200), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1232), .B2(new_n1200), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1222), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1224), .A2(new_n1230), .A3(new_n1118), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1230), .B1(new_n1224), .B2(new_n1118), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1228), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1200), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1210), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1232), .A2(G384), .A3(new_n1200), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(KEYINPUT125), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1235), .A2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT62), .B1(new_n1221), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1216), .A2(G2897), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1235), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G2897), .B(new_n1216), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT61), .B1(new_n1221), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1216), .B1(G375), .B2(G378), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1243), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1250), .A2(new_n1251), .A3(new_n1220), .A4(new_n1252), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1244), .A2(new_n1249), .A3(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G390), .A2(G387), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1255), .A2(new_n1209), .A3(KEYINPUT126), .ZN(new_n1256));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1255), .A2(new_n1209), .A3(KEYINPUT126), .A4(new_n1257), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1254), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT63), .B1(new_n1221), .B2(new_n1243), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT63), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1250), .A2(new_n1265), .A3(new_n1220), .A4(new_n1252), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1261), .A3(new_n1249), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1263), .A2(new_n1268), .ZN(G405));
  NAND2_X1  g1069(.A1(G375), .A2(G378), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n1207), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1222), .A2(KEYINPUT127), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1270), .B(new_n1207), .C1(KEYINPUT127), .C2(new_n1243), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1274), .A2(new_n1261), .A3(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1261), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1276), .A2(new_n1277), .ZN(G402));
endmodule


