//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  NAND2_X1  g035(.A1(new_n455), .A2(G2106), .ZN(new_n461));
  INV_X1    g036(.A(G567), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  AND2_X1   g040(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n467));
  OAI211_X1 g042(.A(KEYINPUT69), .B(G2104), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT68), .A2(KEYINPUT3), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n476), .B1(KEYINPUT3), .B2(new_n470), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n468), .B(new_n469), .C1(new_n475), .C2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G137), .ZN(new_n480));
  NAND2_X1  g055(.A1(G113), .A2(G2104), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n472), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G125), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n470), .A2(G2105), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n486), .A2(G2105), .B1(G101), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G160));
  NAND2_X1  g065(.A1(new_n479), .A2(G136), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n468), .B(G2105), .C1(new_n475), .C2(new_n477), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  MUX2_X1   g069(.A(G100), .B(G112), .S(G2105), .Z(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2104), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n491), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR4_X1   g074(.A1(new_n484), .A2(KEYINPUT4), .A3(new_n499), .A4(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n478), .B2(new_n499), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(new_n466), .B2(new_n467), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n482), .A2(KEYINPUT69), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n506), .A2(G138), .A3(new_n469), .A4(new_n468), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n500), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  MUX2_X1   g084(.A(G102), .B(G114), .S(G2105), .Z(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G2104), .ZN(new_n511));
  INV_X1    g086(.A(G126), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n492), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT70), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  OAI211_X1 g090(.A(new_n515), .B(new_n511), .C1(new_n492), .C2(new_n512), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n509), .A2(new_n517), .ZN(G164));
  OAI21_X1  g093(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT73), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(KEYINPUT72), .A2(KEYINPUT73), .A3(KEYINPUT5), .A4(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT6), .B(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(G88), .B1(G50), .B2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G166));
  NAND2_X1  g111(.A1(new_n526), .A2(G89), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n528), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n539));
  XOR2_X1   g114(.A(KEYINPUT75), .B(KEYINPUT7), .Z(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n540), .B(new_n541), .ZN(new_n542));
  AND4_X1   g117(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n531), .ZN(new_n545));
  INV_X1    g120(.A(G90), .ZN(new_n546));
  INV_X1    g121(.A(G52), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n525), .A2(new_n546), .B1(new_n527), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AND2_X1   g124(.A1(new_n523), .A2(G56), .ZN(new_n550));
  AND2_X1   g125(.A1(G68), .A2(G543), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n526), .A2(G81), .B1(G43), .B2(new_n528), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g134(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G36), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n528), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n523), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n531), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n526), .A2(G91), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  INV_X1    g146(.A(G168), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  NAND2_X1  g148(.A1(new_n526), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n528), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G288));
  AOI22_X1  g152(.A1(new_n526), .A2(G86), .B1(G48), .B2(new_n528), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n523), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n531), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n526), .A2(G85), .B1(G47), .B2(new_n528), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n531), .B2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n526), .A2(G92), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT10), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n586), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n523), .A2(G66), .ZN(new_n589));
  NAND2_X1  g164(.A1(G79), .A2(G543), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n531), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(G54), .B2(new_n528), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(KEYINPUT78), .ZN(new_n595));
  AND3_X1   g170(.A1(new_n588), .A2(KEYINPUT78), .A3(new_n592), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G284));
  XNOR2_X1  g173(.A(G284), .B(KEYINPUT79), .ZN(G321));
  OR2_X1    g174(.A1(G299), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G168), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT80), .ZN(G297));
  INV_X1    g178(.A(new_n602), .ZN(G280));
  XOR2_X1   g179(.A(KEYINPUT81), .B(G559), .Z(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(G860), .B2(new_n605), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT82), .Z(G148));
  NAND2_X1  g182(.A1(new_n597), .A2(new_n605), .ZN(new_n608));
  MUX2_X1   g183(.A(new_n556), .B(new_n608), .S(G868), .Z(G323));
  XNOR2_X1  g184(.A(KEYINPUT83), .B(KEYINPUT11), .ZN(new_n610));
  XNOR2_X1  g185(.A(G323), .B(new_n610), .ZN(G282));
  NAND2_X1  g186(.A1(new_n479), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n493), .A2(G123), .ZN(new_n613));
  AND2_X1   g188(.A1(G111), .A2(G2105), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G99), .B2(new_n469), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n470), .C2(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n469), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(G156));
  XOR2_X1   g198(.A(KEYINPUT15), .B(G2435), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2427), .ZN(new_n626));
  INV_X1    g201(.A(G2430), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n628), .A2(KEYINPUT14), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT85), .ZN(new_n631));
  XNOR2_X1  g206(.A(G1341), .B(G1348), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n633), .A2(new_n638), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n639), .A2(G14), .A3(new_n640), .ZN(G401));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  NOR2_X1   g218(.A1(G2072), .A2(G2078), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n642), .B(new_n643), .C1(new_n444), .C2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n444), .A2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT17), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n643), .B(KEYINPUT86), .ZN(new_n649));
  AND2_X1   g224(.A1(new_n649), .A2(new_n642), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n642), .B1(new_n649), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT87), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n649), .B2(new_n648), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(KEYINPUT87), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(G2096), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(G227));
  XNOR2_X1  g233(.A(G1956), .B(G2474), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n660), .A2(new_n661), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n668), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n664), .A3(new_n662), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n665), .B2(new_n667), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT90), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n676), .B(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NOR2_X1   g256(.A1(G168), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n681), .B2(G21), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT103), .B(G1966), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(G29), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n686), .A2(KEYINPUT91), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(KEYINPUT91), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n616), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT31), .B(G11), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT104), .B(G28), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(new_n686), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n692), .B1(new_n694), .B2(new_n696), .C1(new_n683), .C2(new_n684), .ZN(new_n697));
  NOR2_X1   g272(.A1(G171), .A2(new_n681), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G5), .B2(new_n681), .ZN(new_n699));
  INV_X1    g274(.A(G1961), .ZN(new_n700));
  INV_X1    g275(.A(G2084), .ZN(new_n701));
  NOR2_X1   g276(.A1(KEYINPUT24), .A2(G34), .ZN(new_n702));
  AND2_X1   g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n690), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(new_n489), .B2(new_n686), .ZN(new_n705));
  OAI22_X1  g280(.A1(new_n699), .A2(new_n700), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  NOR3_X1   g281(.A1(new_n691), .A2(new_n697), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n690), .A2(G26), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n479), .A2(G140), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n493), .A2(G128), .ZN(new_n711));
  MUX2_X1   g286(.A(G104), .B(G116), .S(G2105), .Z(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G2104), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n709), .B1(new_n715), .B2(new_n686), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G2067), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n681), .A2(G20), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT23), .Z(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G299), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1956), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(G2067), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n707), .A2(new_n717), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n705), .A2(new_n701), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT105), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n699), .A2(new_n700), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n686), .A2(G32), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT100), .B(KEYINPUT26), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT101), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  AND3_X1   g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n493), .A2(G129), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n730), .A2(new_n732), .B1(G105), .B2(new_n487), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(G141), .B2(new_n479), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT102), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n727), .B1(new_n743), .B2(new_n686), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n725), .B(new_n726), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G115), .A2(G2104), .ZN(new_n750));
  INV_X1    g325(.A(G127), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n484), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT98), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n469), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n753), .B2(new_n752), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n479), .A2(G139), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n487), .A2(G103), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT25), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT99), .Z(new_n760));
  MUX2_X1   g335(.A(G33), .B(new_n760), .S(G29), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(new_n442), .ZN(new_n762));
  NOR2_X1   g337(.A1(G4), .A2(G16), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n597), .B2(G16), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT96), .B(G1348), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n766), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n749), .A2(new_n762), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n744), .A2(new_n746), .ZN(new_n770));
  INV_X1    g345(.A(G2090), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n689), .A2(G35), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n689), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT29), .Z(new_n774));
  AOI21_X1  g349(.A(new_n770), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n681), .A2(G19), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT97), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n557), .B2(new_n681), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1341), .Z(new_n779));
  OAI211_X1 g354(.A(new_n775), .B(new_n779), .C1(new_n771), .C2(new_n774), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n690), .A2(G27), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT107), .Z(new_n782));
  INV_X1    g357(.A(G164), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n689), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT108), .B(G2078), .Z(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n747), .B2(new_n748), .ZN(new_n788));
  OR4_X1    g363(.A1(new_n723), .A2(new_n769), .A3(new_n780), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n681), .A2(G22), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n681), .ZN(new_n791));
  XNOR2_X1  g366(.A(KEYINPUT95), .B(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G6), .A2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G305), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n681), .A2(G23), .ZN(new_n799));
  INV_X1    g374(.A(G288), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n681), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT33), .B(G1976), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n793), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n690), .A2(G25), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT92), .ZN(new_n808));
  MUX2_X1   g383(.A(G95), .B(G107), .S(G2105), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(G2104), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT93), .Z(new_n811));
  NAND2_X1  g386(.A1(new_n493), .A2(G119), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n479), .A2(G131), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT94), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n808), .B1(new_n815), .B2(new_n689), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G24), .B(G290), .S(G16), .Z(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(G1986), .Z(new_n821));
  NAND4_X1  g396(.A1(new_n805), .A2(new_n806), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT36), .Z(new_n823));
  NOR2_X1   g398(.A1(new_n789), .A2(new_n823), .ZN(G311));
  INV_X1    g399(.A(G311), .ZN(G150));
  AOI22_X1  g400(.A1(new_n526), .A2(G93), .B1(G55), .B2(new_n528), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n531), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  INV_X1    g406(.A(new_n829), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n554), .A2(new_n555), .A3(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n832), .B1(new_n554), .B2(new_n555), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT38), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n597), .A2(G559), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n837), .B(new_n838), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n840), .B2(KEYINPUT39), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n831), .B1(new_n841), .B2(new_n843), .ZN(G145));
  NOR2_X1   g419(.A1(new_n743), .A2(new_n715), .ZN(new_n845));
  MUX2_X1   g420(.A(G106), .B(G118), .S(G2105), .Z(new_n846));
  AOI22_X1  g421(.A1(new_n493), .A2(G130), .B1(G2104), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G142), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n478), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(new_n620), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n814), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n742), .A2(new_n714), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n845), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n845), .B2(new_n852), .ZN(new_n854));
  INV_X1    g429(.A(new_n500), .ZN(new_n855));
  AND3_X1   g430(.A1(new_n507), .A2(KEYINPUT71), .A3(KEYINPUT4), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT71), .B1(new_n507), .B2(KEYINPUT4), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n513), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n760), .B(new_n860), .Z(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n853), .A2(new_n854), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G160), .B(new_n497), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n865), .B(new_n616), .Z(new_n866));
  AOI21_X1  g441(.A(new_n862), .B1(new_n853), .B2(new_n854), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n864), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n866), .B1(new_n864), .B2(new_n867), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g447(.A1(new_n829), .A2(G868), .ZN(new_n873));
  XNOR2_X1  g448(.A(G166), .B(new_n795), .ZN(new_n874));
  XNOR2_X1  g449(.A(G290), .B(G288), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n835), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(new_n833), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n608), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n593), .A2(G299), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n593), .A2(G299), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n885), .A2(KEYINPUT41), .A3(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n882), .A2(new_n883), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n879), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n888), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n876), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(new_n876), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n873), .B1(new_n899), .B2(G868), .ZN(G295));
  AOI21_X1  g475(.A(new_n873), .B1(new_n899), .B2(G868), .ZN(G331));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n902));
  NOR2_X1   g477(.A1(G171), .A2(KEYINPUT109), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(G171), .A2(KEYINPUT109), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT110), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n906), .A3(G168), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n906), .B1(new_n905), .B2(G168), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n909), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(new_n903), .A3(new_n907), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n836), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n878), .A2(new_n912), .A3(new_n910), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n887), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT113), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n890), .A3(new_n915), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n876), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(KEYINPUT111), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n914), .A2(new_n915), .A3(new_n922), .A4(new_n890), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n914), .A2(new_n915), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(new_n884), .A3(new_n886), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n876), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n869), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n920), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n916), .B1(new_n921), .B2(new_n923), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n930), .A2(new_n876), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n930), .B2(new_n876), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n902), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT112), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n930), .A2(new_n876), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n936), .B(KEYINPUT43), .C1(new_n928), .C2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n926), .A2(KEYINPUT113), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n916), .A2(new_n917), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n919), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n897), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n933), .A3(new_n932), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n931), .A2(new_n932), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n936), .B1(new_n945), .B2(KEYINPUT43), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n935), .B1(new_n947), .B2(new_n902), .ZN(G397));
  AOI21_X1  g523(.A(G1384), .B1(new_n858), .B2(new_n859), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n480), .A2(G40), .A3(new_n488), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  XNOR2_X1  g526(.A(KEYINPUT114), .B(KEYINPUT45), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n742), .A2(G1996), .ZN(new_n956));
  INV_X1    g531(.A(G2067), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n714), .B(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n955), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1996), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT115), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n743), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(new_n814), .B(new_n817), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n963), .B1(new_n955), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(G290), .B(G1986), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n965), .B1(new_n954), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(new_n950), .C1(new_n509), .C2(new_n513), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n969), .A2(G2067), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n509), .B2(new_n517), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n951), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT117), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT50), .ZN(new_n974));
  AND4_X1   g549(.A1(new_n973), .A2(new_n860), .A3(new_n974), .A4(new_n968), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n973), .B1(new_n949), .B2(new_n974), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n972), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n970), .B1(new_n977), .B2(new_n765), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(G299), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(G299), .B2(new_n983), .ZN(new_n984));
  OAI211_X1 g559(.A(KEYINPUT45), .B(new_n968), .C1(new_n509), .C2(new_n513), .ZN(new_n985));
  INV_X1    g560(.A(new_n517), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n986), .B2(new_n858), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n950), .C1(new_n987), .C2(new_n953), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT56), .B(G2072), .Z(new_n989));
  NAND2_X1  g564(.A1(new_n971), .A2(new_n974), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n949), .A2(KEYINPUT50), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n951), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI221_X1 g567(.A(new_n984), .B1(new_n988), .B2(new_n989), .C1(new_n992), .C2(G1956), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n979), .A2(new_n597), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n984), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n992), .A2(G1956), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n988), .A2(new_n989), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(KEYINPUT58), .B(G1341), .Z(new_n1000));
  NAND2_X1  g575(.A1(new_n969), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(new_n988), .B2(G1996), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n557), .ZN(new_n1003));
  NAND2_X1  g578(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n998), .A2(KEYINPUT61), .A3(new_n993), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT61), .B1(new_n998), .B2(new_n993), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n597), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT60), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n979), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n978), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1011), .B(new_n1012), .C1(KEYINPUT60), .C2(new_n978), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n999), .B1(new_n1008), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT124), .ZN(new_n1015));
  XOR2_X1   g590(.A(KEYINPUT121), .B(G1961), .Z(new_n1016));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n971), .A2(new_n952), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1018), .A2(new_n443), .A3(new_n950), .A4(new_n985), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n977), .A2(new_n1016), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n949), .A2(new_n953), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT122), .B1(new_n1021), .B2(new_n951), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT122), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1023), .B(new_n950), .C1(new_n949), .C2(new_n953), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1017), .A2(G2078), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1022), .A2(new_n985), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1020), .A2(KEYINPUT123), .A3(G301), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1020), .A2(G301), .A3(new_n1026), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n950), .B1(new_n949), .B2(KEYINPUT45), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n971), .A2(new_n952), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1025), .ZN(new_n1034));
  AOI21_X1  g609(.A(G301), .B1(new_n1020), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1030), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1020), .A2(G171), .A3(new_n1026), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n977), .A2(new_n1016), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1019), .A2(new_n1017), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n1034), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1028), .B1(new_n1041), .B2(G301), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n1029), .A2(new_n1037), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n534), .A2(G8), .A3(new_n535), .ZN(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT55), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT116), .B(G1971), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n992), .A2(new_n771), .B1(new_n988), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n988), .A2(new_n1046), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n977), .B2(G2090), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1045), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(G8), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT118), .B1(new_n969), .B2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n969), .A2(KEYINPUT118), .A3(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n800), .A2(G1976), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT52), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1056), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1058), .B(new_n1062), .C1(new_n1063), .C2(new_n1054), .ZN(new_n1064));
  INV_X1    g639(.A(G1981), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n795), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G305), .A2(G1981), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1066), .A2(KEYINPUT49), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT49), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1063), .B2(new_n1054), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1064), .A2(new_n1071), .ZN(new_n1072));
  AND4_X1   g647(.A1(new_n1049), .A2(new_n1053), .A3(new_n1060), .A4(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n701), .B(new_n972), .C1(new_n975), .C2(new_n976), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n684), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(G168), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT51), .ZN(new_n1078));
  AOI21_X1  g653(.A(G168), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  OAI211_X1 g655(.A(G8), .B(new_n1076), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1073), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1015), .B1(new_n1043), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1042), .A2(new_n1038), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1036), .B1(new_n1041), .B2(G171), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n1020), .A2(G301), .A3(new_n1026), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1053), .A2(new_n1049), .A3(new_n1072), .A4(new_n1060), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(KEYINPUT124), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1014), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1072), .A2(new_n1060), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G288), .A2(G1976), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1071), .A2(new_n1096), .B1(new_n1065), .B2(new_n795), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1057), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1095), .A2(new_n1053), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT63), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1101), .A2(G8), .A3(G168), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1091), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1095), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(new_n1100), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1051), .A2(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1045), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1053), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1099), .B1(new_n1103), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1078), .A2(new_n1081), .A3(new_n1110), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1073), .A2(new_n1111), .A3(KEYINPUT125), .A4(new_n1035), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1082), .A2(KEYINPUT62), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1035), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1091), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT125), .B1(new_n1116), .B2(new_n1111), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1109), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n967), .B1(new_n1094), .B2(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n815), .A2(new_n818), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n963), .A2(new_n1120), .B1(new_n957), .B2(new_n715), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1121), .A2(new_n955), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n955), .B1(new_n743), .B2(new_n958), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n962), .B2(KEYINPUT46), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(KEYINPUT46), .B2(new_n962), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n965), .A2(KEYINPUT127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n955), .A2(G1986), .A3(G290), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n1129), .B(KEYINPUT48), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n965), .A2(KEYINPUT127), .ZN(new_n1132));
  AOI211_X1 g707(.A(new_n1122), .B(new_n1127), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1119), .A2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g709(.A1(G401), .A2(G229), .A3(new_n464), .A4(G227), .ZN(new_n1136));
  OAI211_X1 g710(.A(new_n871), .B(new_n1136), .C1(new_n944), .C2(new_n946), .ZN(G225));
  INV_X1    g711(.A(G225), .ZN(G308));
endmodule


