//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g033(.A1(new_n458), .A2(KEYINPUT65), .B1(G567), .B2(new_n454), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n459), .B1(KEYINPUT65), .B2(new_n458), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G125), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT67), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n472), .A2(KEYINPUT3), .A3(new_n473), .ZN(new_n477));
  INV_X1    g052(.A(G2105), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n477), .A2(G137), .A3(new_n478), .A4(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND3_X1  g056(.A1(new_n477), .A2(new_n478), .A3(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n477), .A2(G2105), .A3(new_n464), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n478), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  AND2_X1   g065(.A1(new_n478), .A2(G138), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n477), .A2(new_n464), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n494), .A2(new_n478), .A3(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n467), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n477), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n478), .ZN(new_n501));
  AND2_X1   g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AND2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI22_X1  g096(.A1(new_n518), .A2(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT68), .B(G88), .Z(new_n523));
  OAI22_X1  g098(.A1(new_n516), .A2(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n512), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT7), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT70), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n529), .A2(new_n530), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT69), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G51), .ZN(new_n536));
  AND4_X1   g111(.A1(new_n531), .A2(new_n532), .A3(new_n534), .A4(new_n536), .ZN(G168));
  AOI22_X1  g112(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n511), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n516), .A2(new_n540), .B1(new_n522), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  AOI22_X1  g118(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n511), .ZN(new_n545));
  INV_X1    g120(.A(new_n522), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n546), .A2(G81), .B1(G43), .B2(new_n535), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT71), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n535), .A2(new_n555), .A3(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n522), .A2(KEYINPUT73), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n515), .A2(new_n509), .A3(new_n559), .ZN(new_n560));
  AND2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G91), .ZN(new_n562));
  INV_X1    g137(.A(G78), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n563), .A2(new_n506), .A3(KEYINPUT74), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT74), .B1(new_n563), .B2(new_n506), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n519), .A2(new_n518), .ZN(new_n567));
  OAI211_X1 g142(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n557), .A2(new_n562), .A3(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g146(.A(G171), .B(new_n571), .ZN(G301));
  NAND4_X1  g147(.A1(new_n532), .A2(new_n531), .A3(new_n534), .A4(new_n536), .ZN(G286));
  INV_X1    g148(.A(G166), .ZN(G303));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n511), .B1(new_n567), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(G49), .B2(new_n535), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n558), .A2(G87), .A3(new_n560), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G288));
  AND3_X1   g154(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(KEYINPUT76), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(G61), .B1(new_n519), .B2(new_n518), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(G48), .B2(new_n535), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n558), .A2(G86), .A3(new_n560), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n546), .A2(G85), .B1(G47), .B2(new_n535), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OAI22_X1  g166(.A1(new_n589), .A2(new_n590), .B1(new_n511), .B2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n561), .A2(G92), .ZN(new_n593));
  XNOR2_X1  g168(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n594), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n567), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n535), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  MUX2_X1   g177(.A(G301), .B(new_n601), .S(new_n602), .Z(G321));
  XNOR2_X1  g178(.A(G321), .B(KEYINPUT79), .ZN(G284));
  NAND2_X1  g179(.A1(G299), .A2(new_n602), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G168), .B2(new_n602), .ZN(G297));
  OAI21_X1  g181(.A(new_n605), .B1(G168), .B2(new_n602), .ZN(G280));
  INV_X1    g182(.A(new_n601), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT80), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(new_n602), .ZN(new_n613));
  AOI21_X1  g188(.A(new_n613), .B1(new_n602), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g190(.A1(new_n474), .A2(new_n464), .A3(new_n466), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n483), .A2(G135), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT82), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n478), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AOI22_X1  g200(.A1(new_n485), .A2(G123), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n620), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XOR2_X1   g205(.A(KEYINPUT15), .B(G2435), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2438), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT84), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n641), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n661), .A2(new_n666), .A3(new_n664), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n666), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n669));
  AOI211_X1 g244(.A(new_n665), .B(new_n667), .C1(new_n668), .C2(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n668), .B2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NOR2_X1   g253(.A1(G166), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n678), .B2(G22), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G1971), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(G1971), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n678), .A2(G6), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G305), .B2(G16), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT32), .B(G1981), .Z(new_n686));
  OAI211_X1 g261(.A(new_n682), .B(new_n683), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n688), .A2(new_n678), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n678), .B2(G23), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT33), .B(G1976), .Z(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n685), .A2(new_n686), .ZN(new_n694));
  AND2_X1   g269(.A1(new_n690), .A2(new_n692), .ZN(new_n695));
  NOR4_X1   g270(.A1(new_n687), .A2(new_n693), .A3(new_n694), .A4(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT34), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  MUX2_X1   g274(.A(G24), .B(G290), .S(G16), .Z(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(G1986), .Z(new_n701));
  NAND2_X1  g276(.A1(new_n483), .A2(G131), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n485), .A2(G119), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n478), .A2(G107), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n702), .B(new_n703), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G29), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT86), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT36), .ZN(new_n715));
  NAND2_X1  g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  INV_X1    g291(.A(G127), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n467), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(G2105), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n478), .A2(G103), .A3(G2104), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT25), .Z(new_n721));
  INV_X1    g296(.A(G139), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n721), .C1(new_n482), .C2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT89), .Z(new_n724));
  MUX2_X1   g299(.A(G33), .B(new_n724), .S(G29), .Z(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G2072), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G35), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G162), .B2(G29), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n736), .B2(KEYINPUT24), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT24), .B2(new_n736), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n480), .B2(new_n708), .ZN(new_n739));
  INV_X1    g314(.A(G2084), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n627), .A2(new_n708), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(KEYINPUT31), .B(G11), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n708), .B1(new_n743), .B2(G28), .ZN(new_n745));
  NOR2_X1   g320(.A1(G5), .A2(G16), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT92), .Z(new_n747));
  INV_X1    g322(.A(G171), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n678), .ZN(new_n749));
  INV_X1    g324(.A(G1961), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n742), .B1(new_n744), .B2(new_n745), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n741), .B(new_n751), .C1(new_n740), .C2(new_n739), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G19), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n548), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n750), .B2(new_n749), .ZN(new_n756));
  INV_X1    g331(.A(G1966), .ZN(new_n757));
  NOR2_X1   g332(.A1(G168), .A2(new_n678), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n678), .B2(G21), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n752), .B(new_n756), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n731), .A2(new_n732), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n678), .A2(G20), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT95), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT23), .ZN(new_n764));
  AND3_X1   g339(.A1(new_n557), .A2(new_n562), .A3(new_n569), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n678), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n759), .A2(new_n757), .B1(new_n766), .B2(G1956), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G1956), .B2(new_n766), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n760), .A2(new_n761), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n678), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n608), .B2(new_n678), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT87), .B(G1348), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n708), .A2(G32), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n483), .A2(G141), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT91), .ZN(new_n776));
  NAND3_X1  g351(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT26), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n474), .A2(G105), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G129), .B2(new_n485), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n708), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT27), .B(G1996), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n771), .A2(new_n773), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n708), .A2(G27), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G164), .B2(new_n708), .ZN(new_n788));
  INV_X1    g363(.A(G2078), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n786), .B(new_n790), .C1(new_n773), .C2(new_n771), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n483), .A2(G140), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n485), .A2(G128), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n478), .A2(G116), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G29), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n708), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT88), .B(G2067), .Z(new_n801));
  XOR2_X1   g376(.A(new_n800), .B(new_n801), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n725), .A2(G2072), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n784), .B2(new_n785), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n791), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n715), .A2(new_n735), .A3(new_n769), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n608), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n511), .ZN(new_n811));
  INV_X1    g386(.A(G55), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  OAI22_X1  g388(.A1(new_n516), .A2(new_n812), .B1(new_n522), .B2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n548), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n809), .B(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n819));
  INV_X1    g394(.A(G860), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(KEYINPUT39), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n815), .A2(new_n820), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT37), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  XNOR2_X1  g400(.A(new_n783), .B(new_n724), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n706), .B(new_n618), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n724), .B(new_n782), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(new_n827), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(G164), .B(new_n796), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n483), .A2(G142), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n485), .A2(G130), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n478), .A2(G118), .ZN(new_n836));
  OAI21_X1  g411(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n833), .B(new_n838), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n480), .B(new_n489), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n627), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n829), .A2(new_n839), .A3(new_n831), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n841), .B2(new_n844), .ZN(new_n848));
  OAI21_X1  g423(.A(KEYINPUT96), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n848), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n850), .A2(new_n851), .A3(new_n846), .A4(new_n845), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g429(.A(KEYINPUT103), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(new_n815), .B2(G868), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n601), .A2(G299), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n765), .A2(new_n595), .A3(new_n596), .A4(new_n600), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n859), .A2(KEYINPUT100), .A3(new_n860), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n859), .B2(KEYINPUT41), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT41), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT98), .A4(new_n867), .ZN(new_n868));
  AOI22_X1  g443(.A1(new_n863), .A2(new_n864), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n859), .B(KEYINPUT97), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n548), .B(new_n815), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n612), .B(new_n871), .ZN(new_n872));
  MUX2_X1   g447(.A(new_n869), .B(new_n870), .S(new_n872), .Z(new_n873));
  XOR2_X1   g448(.A(G288), .B(KEYINPUT101), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(G290), .ZN(new_n875));
  XNOR2_X1  g450(.A(G166), .B(G305), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT102), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n602), .B1(new_n873), .B2(new_n881), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n856), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(KEYINPUT103), .B2(new_n885), .ZN(G295));
  AOI21_X1  g461(.A(new_n884), .B1(KEYINPUT103), .B2(new_n885), .ZN(G331));
  NOR2_X1   g462(.A1(G301), .A2(G286), .ZN(new_n888));
  NAND2_X1  g463(.A1(G286), .A2(new_n748), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n871), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n892));
  XNOR2_X1  g467(.A(G171), .B(KEYINPUT75), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G168), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n817), .A3(new_n889), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(KEYINPUT104), .B(new_n871), .C1(new_n888), .C2(new_n890), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n859), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n891), .A2(new_n895), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n899), .B1(new_n869), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n880), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n863), .A2(new_n864), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n866), .A2(new_n868), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n880), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n898), .A2(KEYINPUT105), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n899), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(new_n910), .A3(new_n846), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT43), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n859), .A2(new_n867), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n896), .A2(new_n897), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(new_n870), .B2(new_n900), .ZN(new_n917));
  AOI21_X1  g492(.A(G37), .B1(new_n917), .B2(new_n880), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n910), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT106), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  AOI211_X1 g498(.A(new_n923), .B(KEYINPUT44), .C1(new_n912), .C2(new_n919), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n913), .B1(new_n910), .B2(new_n918), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n910), .A2(new_n913), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n846), .A3(new_n904), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT44), .ZN(new_n928));
  OAI22_X1  g503(.A1(new_n922), .A2(new_n924), .B1(new_n925), .B2(new_n928), .ZN(G397));
  INV_X1    g504(.A(G1384), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n496), .B1(new_n492), .B2(KEYINPUT4), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n499), .A2(new_n501), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT45), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n470), .A2(G40), .A3(new_n479), .A4(new_n475), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  OAI211_X1 g512(.A(KEYINPUT45), .B(new_n930), .C1(new_n931), .C2(new_n932), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g514(.A(KEYINPUT108), .B(G1971), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n936), .B1(new_n933), .B2(KEYINPUT50), .ZN(new_n942));
  NOR2_X1   g517(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n943), .B1(new_n931), .B2(new_n932), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n732), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(G8), .ZN(new_n947));
  XNOR2_X1  g522(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(G8), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n949), .B1(G166), .B2(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(G8), .B(new_n948), .C1(new_n512), .C2(new_n524), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n954), .B1(new_n503), .B2(new_n943), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n954), .B(new_n943), .C1(new_n931), .C2(new_n932), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n732), .B(new_n942), .C1(new_n955), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n950), .B1(new_n941), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n953), .A2(KEYINPUT111), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n961), .A3(new_n952), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n947), .A2(new_n953), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(G1384), .B1(new_n498), .B2(new_n502), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n937), .ZN(new_n966));
  INV_X1    g541(.A(G1976), .ZN(new_n967));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(G288), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n577), .A2(G1976), .A3(new_n578), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n966), .A2(new_n968), .A3(G8), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(G8), .B(new_n969), .C1(new_n933), .C2(new_n936), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT52), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT112), .B(G1981), .Z(new_n973));
  NAND3_X1  g548(.A1(new_n585), .A2(new_n586), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G61), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n507), .B2(new_n508), .ZN(new_n976));
  NAND2_X1  g551(.A1(G73), .A2(G543), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT76), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(KEYINPUT76), .A2(G73), .A3(G543), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(G651), .B1(new_n976), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n535), .A2(G48), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n515), .A2(new_n509), .A3(G86), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(G1981), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n974), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n950), .B1(new_n965), .B2(new_n937), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n989), .B1(new_n987), .B2(new_n988), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n970), .B(new_n972), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT115), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n987), .A2(new_n988), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT49), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n997), .A2(new_n991), .A3(new_n990), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n970), .A4(new_n972), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n964), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n944), .A2(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n956), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n942), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n750), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n936), .A2(KEYINPUT120), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n936), .B2(KEYINPUT120), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1007), .A2(new_n935), .A3(new_n1009), .A4(new_n938), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n939), .B2(G2078), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1006), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1013), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT121), .B1(new_n1013), .B2(G171), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1012), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT119), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1006), .B(new_n1019), .C1(new_n939), .C2(new_n1008), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n939), .A2(new_n1008), .ZN(new_n1021));
  AOI21_X1  g596(.A(G1961), .B1(new_n1004), .B2(new_n942), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT119), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1018), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G301), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1002), .B1(new_n1017), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n939), .A2(new_n757), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1004), .A2(new_n740), .A3(new_n942), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1027), .A2(new_n1028), .A3(G168), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  AOI21_X1  g605(.A(G168), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT51), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT118), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1029), .A2(new_n1034), .A3(G8), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1033), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT57), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n765), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n935), .A2(new_n937), .A3(new_n938), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1956), .B1(new_n942), .B2(new_n944), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n942), .A2(new_n944), .ZN(new_n1048));
  INV_X1    g623(.A(G1956), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(new_n1044), .A3(new_n1041), .A4(new_n1040), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT61), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n773), .B1(new_n1004), .B2(new_n942), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n966), .A2(G2067), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1052), .A2(new_n1053), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1056), .A2(new_n601), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n608), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1060));
  OAI21_X1  g635(.A(KEYINPUT60), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n1044), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1064), .A3(new_n1042), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1065), .A2(KEYINPUT61), .A3(new_n1051), .ZN(new_n1066));
  INV_X1    g641(.A(new_n966), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT58), .B(G1341), .ZN(new_n1068));
  OAI22_X1  g643(.A1(new_n939), .A2(G1996), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n548), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT59), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1069), .A2(new_n1072), .A3(new_n548), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1058), .A2(new_n1061), .A3(new_n1066), .A4(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1065), .B1(new_n601), .B2(new_n1056), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1051), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1024), .A2(G301), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1013), .A2(new_n893), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1016), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1026), .A2(new_n1038), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G286), .A2(new_n950), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n964), .A2(new_n1001), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n941), .A2(new_n958), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1089), .A2(G8), .A3(new_n963), .ZN(new_n1090));
  INV_X1    g665(.A(new_n953), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1089), .B2(G8), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1083), .A2(new_n1084), .A3(KEYINPUT63), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1090), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n1095));
  XNOR2_X1  g670(.A(new_n994), .B(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n998), .A2(new_n967), .A3(new_n688), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n974), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n991), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n994), .B(KEYINPUT114), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1090), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT116), .B1(new_n1098), .B2(new_n1105), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1086), .A2(new_n1087), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1104), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1082), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT122), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT122), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1082), .B(new_n1112), .C1(new_n1106), .C2(new_n1109), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1079), .A2(new_n1001), .A3(new_n964), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1038), .B2(KEYINPUT62), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1116), .A2(new_n1121), .A3(KEYINPUT62), .A4(new_n1117), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT124), .B(new_n1120), .C1(new_n1122), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1116), .A2(KEYINPUT62), .A3(new_n1117), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1123), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT124), .B1(new_n1129), .B2(new_n1120), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1111), .B(new_n1113), .C1(new_n1126), .C2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n935), .A2(new_n936), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n782), .B(G1996), .Z(new_n1134));
  XOR2_X1   g709(.A(new_n796), .B(G2067), .Z(new_n1135));
  AND2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n706), .B(new_n712), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1133), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g713(.A(G290), .B(G1986), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1132), .B2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1140), .B(KEYINPUT107), .Z(new_n1141));
  NAND2_X1  g716(.A1(new_n1131), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n796), .A2(G2067), .ZN(new_n1143));
  INV_X1    g718(.A(new_n712), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n706), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1136), .B2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1133), .A2(G1986), .A3(G290), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT125), .B(KEYINPUT48), .Z(new_n1148));
  XNOR2_X1  g723(.A(new_n1147), .B(new_n1148), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1133), .A2(new_n1146), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1133), .B1(new_n1135), .B2(new_n783), .ZN(new_n1151));
  OR3_X1    g726(.A1(new_n1133), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT46), .B1(new_n1133), .B2(G1996), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT47), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1150), .A2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n1156), .B(KEYINPUT126), .Z(new_n1157));
  NAND2_X1  g732(.A1(new_n1142), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  AOI22_X1  g733(.A1(new_n918), .A2(new_n926), .B1(new_n911), .B2(KEYINPUT43), .ZN(new_n1160));
  OR3_X1    g734(.A1(G401), .A2(new_n460), .A3(G227), .ZN(new_n1161));
  NOR2_X1   g735(.A1(G229), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n853), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g737(.A(KEYINPUT127), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1165));
  NAND4_X1  g739(.A1(new_n920), .A2(new_n1165), .A3(new_n853), .A4(new_n1162), .ZN(new_n1166));
  AND2_X1   g740(.A1(new_n1164), .A2(new_n1166), .ZN(G308));
  NAND3_X1  g741(.A1(new_n920), .A2(new_n853), .A3(new_n1162), .ZN(G225));
endmodule


