

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771;

  XNOR2_X1 U374 ( .A(KEYINPUT32), .B(n540), .ZN(n766) );
  INV_X1 U375 ( .A(n695), .ZN(n547) );
  INV_X1 U376 ( .A(n696), .ZN(n533) );
  XOR2_X1 U377 ( .A(n575), .B(n596), .Z(n679) );
  XNOR2_X1 U378 ( .A(n375), .B(G146), .ZN(n473) );
  INV_X1 U379 ( .A(G953), .ZN(n756) );
  XNOR2_X1 U380 ( .A(n531), .B(n530), .ZN(n768) );
  NOR2_X2 U381 ( .A1(n634), .A2(n742), .ZN(n636) );
  NOR2_X2 U382 ( .A1(n732), .A2(n742), .ZN(n733) );
  XNOR2_X2 U383 ( .A(n433), .B(n749), .ZN(n637) );
  XNOR2_X2 U384 ( .A(n427), .B(KEYINPUT45), .ZN(n743) );
  XNOR2_X2 U385 ( .A(n430), .B(n479), .ZN(n749) );
  XNOR2_X2 U386 ( .A(n473), .B(n459), .ZN(n725) );
  AND2_X2 U387 ( .A1(n547), .A2(n533), .ZN(n545) );
  INV_X1 U388 ( .A(n550), .ZN(n699) );
  NOR2_X1 U389 ( .A1(n720), .A2(G953), .ZN(n721) );
  AND2_X1 U390 ( .A1(n642), .A2(n641), .ZN(n644) );
  NOR2_X1 U391 ( .A1(n717), .A2(n716), .ZN(n719) );
  AND2_X1 U392 ( .A1(n677), .A2(n676), .ZN(n717) );
  AND2_X1 U393 ( .A1(n422), .A2(n423), .ZN(n421) );
  XNOR2_X1 U394 ( .A(n584), .B(KEYINPUT107), .ZN(n684) );
  XNOR2_X1 U395 ( .A(n416), .B(n415), .ZN(n480) );
  XNOR2_X1 U396 ( .A(G116), .B(KEYINPUT69), .ZN(n465) );
  XNOR2_X2 U397 ( .A(n585), .B(n586), .ZN(n707) );
  XNOR2_X2 U398 ( .A(n367), .B(KEYINPUT22), .ZN(n559) );
  NOR2_X2 U399 ( .A1(n549), .A2(n532), .ZN(n367) );
  XNOR2_X1 U400 ( .A(n489), .B(n436), .ZN(n574) );
  XOR2_X1 U401 ( .A(n456), .B(n513), .Z(n754) );
  XNOR2_X1 U402 ( .A(n475), .B(n356), .ZN(n550) );
  OR2_X1 U403 ( .A1(n631), .A2(G902), .ZN(n475) );
  XNOR2_X1 U404 ( .A(n614), .B(n369), .ZN(n392) );
  INV_X1 U405 ( .A(KEYINPUT66), .ZN(n369) );
  XNOR2_X1 U406 ( .A(KEYINPUT88), .B(KEYINPUT15), .ZN(n448) );
  NAND2_X1 U407 ( .A1(n460), .A2(G902), .ZN(n412) );
  XNOR2_X1 U408 ( .A(n398), .B(n396), .ZN(n521) );
  XNOR2_X1 U409 ( .A(KEYINPUT78), .B(KEYINPUT8), .ZN(n398) );
  NOR2_X1 U410 ( .A1(n397), .A2(G953), .ZN(n396) );
  INV_X1 U411 ( .A(G234), .ZN(n397) );
  NOR2_X1 U412 ( .A1(G953), .A2(G237), .ZN(n503) );
  XNOR2_X1 U413 ( .A(n526), .B(n455), .ZN(n375) );
  XNOR2_X1 U414 ( .A(KEYINPUT4), .B(G131), .ZN(n455) );
  XOR2_X1 U415 ( .A(G137), .B(G140), .Z(n456) );
  XNOR2_X1 U416 ( .A(n482), .B(n365), .ZN(n364) );
  INV_X1 U417 ( .A(KEYINPUT4), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n373), .B(G125), .ZN(n481) );
  INV_X1 U419 ( .A(G146), .ZN(n373) );
  INV_X1 U420 ( .A(KEYINPUT68), .ZN(n463) );
  XNOR2_X1 U421 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n441) );
  XNOR2_X1 U422 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U423 ( .A(G128), .B(KEYINPUT94), .ZN(n440) );
  XNOR2_X1 U424 ( .A(KEYINPUT93), .B(KEYINPUT73), .ZN(n439) );
  XNOR2_X1 U425 ( .A(G119), .B(G110), .ZN(n437) );
  XNOR2_X1 U426 ( .A(n481), .B(n372), .ZN(n513) );
  INV_X1 U427 ( .A(KEYINPUT10), .ZN(n372) );
  INV_X1 U428 ( .A(n456), .ZN(n414) );
  XNOR2_X1 U429 ( .A(G104), .B(G107), .ZN(n415) );
  XNOR2_X1 U430 ( .A(n417), .B(G110), .ZN(n416) );
  INV_X1 U431 ( .A(G101), .ZN(n417) );
  AND2_X1 U432 ( .A1(n609), .A2(n610), .ZN(n385) );
  NAND2_X1 U433 ( .A1(n384), .A2(KEYINPUT36), .ZN(n383) );
  INV_X1 U434 ( .A(n609), .ZN(n384) );
  NOR2_X1 U435 ( .A1(n739), .A2(G902), .ZN(n451) );
  XNOR2_X1 U436 ( .A(n550), .B(n476), .ZN(n604) );
  NOR2_X1 U437 ( .A1(n770), .A2(n394), .ZN(n393) );
  OR2_X1 U438 ( .A1(n769), .A2(KEYINPUT46), .ZN(n394) );
  NAND2_X1 U439 ( .A1(G234), .A2(G237), .ZN(n492) );
  INV_X1 U440 ( .A(KEYINPUT34), .ZN(n426) );
  INV_X1 U441 ( .A(G237), .ZN(n486) );
  NAND2_X1 U442 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U443 ( .A1(n410), .A2(n528), .ZN(n409) );
  INV_X1 U444 ( .A(KEYINPUT48), .ZN(n395) );
  XNOR2_X1 U445 ( .A(KEYINPUT3), .B(G119), .ZN(n464) );
  AND2_X1 U446 ( .A1(n743), .A2(n418), .ZN(n389) );
  AND2_X1 U447 ( .A1(n502), .A2(n426), .ZN(n425) );
  NOR2_X1 U448 ( .A1(n502), .A2(n426), .ZN(n424) );
  OR2_X1 U449 ( .A1(n409), .A2(KEYINPUT1), .ZN(n403) );
  XNOR2_X1 U450 ( .A(KEYINPUT5), .B(G137), .ZN(n469) );
  XNOR2_X1 U451 ( .A(n482), .B(G134), .ZN(n526) );
  XOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n507) );
  XNOR2_X1 U453 ( .A(G143), .B(G140), .ZN(n506) );
  XNOR2_X1 U454 ( .A(G113), .B(G131), .ZN(n510) );
  XOR2_X1 U455 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n505) );
  XNOR2_X1 U456 ( .A(n434), .B(n483), .ZN(n433) );
  XNOR2_X1 U457 ( .A(n358), .B(n364), .ZN(n434) );
  NOR2_X1 U458 ( .A1(n744), .A2(KEYINPUT2), .ZN(n366) );
  NOR2_X1 U459 ( .A1(n353), .A2(n675), .ZN(n677) );
  XNOR2_X1 U460 ( .A(n577), .B(n576), .ZN(n615) );
  XNOR2_X1 U461 ( .A(n480), .B(n431), .ZN(n430) );
  XNOR2_X1 U462 ( .A(n432), .B(G122), .ZN(n431) );
  INV_X1 U463 ( .A(KEYINPUT16), .ZN(n432) );
  XNOR2_X1 U464 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U465 ( .A(n438), .B(n437), .ZN(n446) );
  XNOR2_X1 U466 ( .A(n480), .B(n414), .ZN(n458) );
  NOR2_X1 U467 ( .A1(n756), .A2(G952), .ZN(n742) );
  XNOR2_X1 U468 ( .A(n578), .B(KEYINPUT40), .ZN(n770) );
  NOR2_X1 U469 ( .A1(n615), .A2(n660), .ZN(n578) );
  NAND2_X1 U470 ( .A1(n382), .A2(n381), .ZN(n667) );
  AND2_X1 U471 ( .A1(n380), .A2(n360), .ZN(n382) );
  INV_X1 U472 ( .A(KEYINPUT35), .ZN(n530) );
  NAND2_X1 U473 ( .A1(n420), .A2(KEYINPUT34), .ZN(n419) );
  AND2_X1 U474 ( .A1(n559), .A2(n371), .ZN(n540) );
  AND2_X1 U475 ( .A1(n355), .A2(n539), .ZN(n371) );
  XNOR2_X1 U476 ( .A(n536), .B(n535), .ZN(n374) );
  NOR2_X1 U477 ( .A1(n604), .A2(n390), .ZN(n557) );
  AND2_X1 U478 ( .A1(n770), .A2(KEYINPUT46), .ZN(n351) );
  XOR2_X1 U479 ( .A(n450), .B(KEYINPUT25), .Z(n352) );
  AND2_X1 U480 ( .A1(n673), .A2(KEYINPUT2), .ZN(n353) );
  AND2_X1 U481 ( .A1(n404), .A2(n402), .ZN(n354) );
  XNOR2_X1 U482 ( .A(KEYINPUT75), .B(n604), .ZN(n355) );
  XOR2_X1 U483 ( .A(n474), .B(KEYINPUT70), .Z(n356) );
  XOR2_X1 U484 ( .A(n597), .B(KEYINPUT74), .Z(n357) );
  XOR2_X1 U485 ( .A(n485), .B(n484), .Z(n358) );
  OR2_X1 U486 ( .A1(n580), .A2(n579), .ZN(n359) );
  AND2_X1 U487 ( .A1(n612), .A2(n383), .ZN(n360) );
  AND2_X1 U488 ( .A1(n392), .A2(n391), .ZN(n361) );
  AND2_X1 U489 ( .A1(n573), .A2(n679), .ZN(n362) );
  XNOR2_X1 U490 ( .A(n478), .B(KEYINPUT33), .ZN(n688) );
  AND2_X1 U491 ( .A1(n625), .A2(n629), .ZN(n363) );
  AND2_X1 U492 ( .A1(n544), .A2(KEYINPUT83), .ZN(n400) );
  NOR2_X2 U493 ( .A1(n650), .A2(n766), .ZN(n543) );
  NOR2_X1 U494 ( .A1(n400), .A2(n401), .ZN(n370) );
  NAND2_X1 U495 ( .A1(n428), .A2(n370), .ZN(n427) );
  XNOR2_X1 U496 ( .A(n366), .B(KEYINPUT79), .ZN(n676) );
  NAND2_X1 U497 ( .A1(n563), .A2(n562), .ZN(n401) );
  NAND2_X1 U498 ( .A1(n421), .A2(n419), .ZN(n531) );
  NOR2_X1 U499 ( .A1(n424), .A2(n357), .ZN(n423) );
  NAND2_X1 U500 ( .A1(n543), .A2(n768), .ZN(n541) );
  NAND2_X1 U501 ( .A1(n368), .A2(n595), .ZN(n603) );
  OR2_X1 U502 ( .A1(n594), .A2(KEYINPUT47), .ZN(n368) );
  NOR2_X2 U503 ( .A1(n589), .A2(n588), .ZN(n657) );
  XNOR2_X2 U504 ( .A(n608), .B(n491), .ZN(n589) );
  NAND2_X1 U505 ( .A1(n574), .A2(n678), .ZN(n608) );
  AND2_X2 U506 ( .A1(n376), .A2(n623), .ZN(n755) );
  XOR2_X1 U507 ( .A(n548), .B(KEYINPUT95), .Z(n565) );
  XNOR2_X1 U508 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U509 ( .A1(n361), .A2(n378), .ZN(n377) );
  XNOR2_X1 U510 ( .A(n377), .B(n395), .ZN(n376) );
  NOR2_X2 U511 ( .A1(n374), .A2(n691), .ZN(n650) );
  XNOR2_X1 U512 ( .A(n375), .B(n754), .ZN(n759) );
  NOR2_X1 U513 ( .A1(n393), .A2(n351), .ZN(n378) );
  NAND2_X1 U514 ( .A1(n379), .A2(KEYINPUT36), .ZN(n381) );
  INV_X1 U515 ( .A(n617), .ZN(n379) );
  NAND2_X1 U516 ( .A1(n617), .A2(n385), .ZN(n380) );
  NAND2_X1 U517 ( .A1(n613), .A2(n667), .ZN(n614) );
  NAND2_X1 U518 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X2 U519 ( .A(n386), .B(KEYINPUT64), .ZN(n738) );
  NAND2_X1 U520 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U521 ( .A1(n672), .A2(n363), .ZN(n387) );
  NAND2_X1 U522 ( .A1(n389), .A2(n755), .ZN(n388) );
  NAND2_X1 U523 ( .A1(n755), .A2(n743), .ZN(n672) );
  NOR2_X1 U524 ( .A1(n359), .A2(n691), .ZN(n605) );
  INV_X1 U525 ( .A(n691), .ZN(n390) );
  XNOR2_X2 U526 ( .A(n451), .B(n352), .ZN(n691) );
  NAND2_X1 U527 ( .A1(n769), .A2(KEYINPUT46), .ZN(n391) );
  NAND2_X1 U528 ( .A1(n399), .A2(n573), .ZN(n599) );
  NAND2_X1 U529 ( .A1(n399), .A2(n362), .ZN(n577) );
  XNOR2_X1 U530 ( .A(n565), .B(n564), .ZN(n399) );
  OR2_X1 U531 ( .A1(n725), .A2(n409), .ZN(n408) );
  INV_X1 U532 ( .A(n405), .ZN(n411) );
  OR2_X1 U533 ( .A1(n725), .A2(n403), .ZN(n402) );
  NAND2_X1 U534 ( .A1(n405), .A2(n461), .ZN(n404) );
  NAND2_X1 U535 ( .A1(n413), .A2(n412), .ZN(n405) );
  NAND2_X1 U536 ( .A1(n411), .A2(n408), .ZN(n582) );
  NAND2_X2 U537 ( .A1(n354), .A2(n406), .ZN(n696) );
  NAND2_X1 U538 ( .A1(n407), .A2(n411), .ZN(n406) );
  AND2_X1 U539 ( .A1(n408), .A2(KEYINPUT1), .ZN(n407) );
  INV_X1 U540 ( .A(n460), .ZN(n410) );
  NAND2_X1 U541 ( .A1(n725), .A2(n460), .ZN(n413) );
  AND2_X1 U542 ( .A1(n626), .A2(n629), .ZN(n418) );
  INV_X1 U543 ( .A(n688), .ZN(n420) );
  NAND2_X1 U544 ( .A1(n688), .A2(n425), .ZN(n422) );
  NAND2_X1 U545 ( .A1(n429), .A2(n542), .ZN(n428) );
  XNOR2_X1 U546 ( .A(n541), .B(KEYINPUT44), .ZN(n429) );
  NAND2_X1 U547 ( .A1(n637), .A2(n628), .ZN(n489) );
  XOR2_X1 U548 ( .A(n637), .B(n639), .Z(n435) );
  XOR2_X1 U549 ( .A(n488), .B(n487), .Z(n436) );
  INV_X1 U550 ( .A(KEYINPUT18), .ZN(n484) );
  INV_X1 U551 ( .A(KEYINPUT103), .ZN(n462) );
  XNOR2_X1 U552 ( .A(n545), .B(n462), .ZN(n477) );
  INV_X1 U553 ( .A(KEYINPUT106), .ZN(n564) );
  INV_X1 U554 ( .A(KEYINPUT120), .ZN(n718) );
  INV_X1 U555 ( .A(n742), .ZN(n641) );
  INV_X1 U556 ( .A(KEYINPUT63), .ZN(n635) );
  NAND2_X1 U557 ( .A1(G221), .A2(n521), .ZN(n438) );
  XOR2_X1 U558 ( .A(KEYINPUT77), .B(KEYINPUT92), .Z(n442) );
  XNOR2_X1 U559 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U560 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U561 ( .A(n447), .B(n754), .ZN(n739) );
  XNOR2_X2 U562 ( .A(n448), .B(G902), .ZN(n628) );
  NAND2_X1 U563 ( .A1(G234), .A2(n628), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n449), .B(KEYINPUT20), .ZN(n452) );
  AND2_X1 U565 ( .A1(G217), .A2(n452), .ZN(n450) );
  NAND2_X1 U566 ( .A1(G221), .A2(n452), .ZN(n454) );
  INV_X1 U567 ( .A(KEYINPUT21), .ZN(n453) );
  XNOR2_X1 U568 ( .A(n454), .B(n453), .ZN(n690) );
  XNOR2_X2 U569 ( .A(G143), .B(G128), .ZN(n482) );
  NAND2_X1 U570 ( .A1(G227), .A2(n756), .ZN(n457) );
  XNOR2_X1 U571 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U572 ( .A(KEYINPUT67), .B(G469), .Z(n460) );
  INV_X1 U573 ( .A(KEYINPUT1), .ZN(n461) );
  XNOR2_X1 U574 ( .A(n464), .B(n463), .ZN(n467) );
  XNOR2_X1 U575 ( .A(n465), .B(G113), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n467), .B(n466), .ZN(n479) );
  NAND2_X1 U577 ( .A1(n503), .A2(G210), .ZN(n468) );
  XNOR2_X1 U578 ( .A(n468), .B(G101), .ZN(n470) );
  XNOR2_X1 U579 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U580 ( .A(n479), .B(n471), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n473), .B(n472), .ZN(n631) );
  XNOR2_X1 U582 ( .A(G472), .B(KEYINPUT96), .ZN(n474) );
  XNOR2_X1 U583 ( .A(KEYINPUT100), .B(KEYINPUT6), .ZN(n476) );
  NAND2_X1 U584 ( .A1(n477), .A2(n604), .ZN(n478) );
  XOR2_X1 U585 ( .A(KEYINPUT72), .B(KEYINPUT19), .Z(n491) );
  XOR2_X1 U586 ( .A(n481), .B(KEYINPUT17), .Z(n483) );
  NAND2_X1 U587 ( .A1(G224), .A2(n756), .ZN(n485) );
  INV_X1 U588 ( .A(G902), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n528), .A2(n486), .ZN(n490) );
  NAND2_X1 U590 ( .A1(n490), .A2(G210), .ZN(n488) );
  INV_X1 U591 ( .A(KEYINPUT89), .ZN(n487) );
  NAND2_X1 U592 ( .A1(n490), .A2(G214), .ZN(n678) );
  XNOR2_X1 U593 ( .A(n492), .B(KEYINPUT14), .ZN(n494) );
  NAND2_X1 U594 ( .A1(G952), .A2(n494), .ZN(n493) );
  XNOR2_X1 U595 ( .A(KEYINPUT90), .B(n493), .ZN(n713) );
  NOR2_X1 U596 ( .A1(G953), .A2(n713), .ZN(n571) );
  INV_X1 U597 ( .A(n571), .ZN(n497) );
  NAND2_X1 U598 ( .A1(G902), .A2(n494), .ZN(n567) );
  INV_X1 U599 ( .A(n567), .ZN(n495) );
  NOR2_X1 U600 ( .A1(G898), .A2(n756), .ZN(n751) );
  NAND2_X1 U601 ( .A1(n495), .A2(n751), .ZN(n496) );
  NAND2_X1 U602 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U603 ( .A(KEYINPUT91), .B(n498), .ZN(n499) );
  NOR2_X2 U604 ( .A1(n589), .A2(n499), .ZN(n501) );
  XNOR2_X1 U605 ( .A(KEYINPUT85), .B(KEYINPUT0), .ZN(n500) );
  XNOR2_X2 U606 ( .A(n501), .B(n500), .ZN(n549) );
  INV_X1 U607 ( .A(n549), .ZN(n502) );
  NAND2_X1 U608 ( .A1(G214), .A2(n503), .ZN(n504) );
  XNOR2_X1 U609 ( .A(n505), .B(n504), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U611 ( .A(n509), .B(n508), .Z(n515) );
  XOR2_X1 U612 ( .A(G104), .B(G122), .Z(n511) );
  XNOR2_X1 U613 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n513), .B(n512), .ZN(n514) );
  XNOR2_X1 U615 ( .A(n515), .B(n514), .ZN(n729) );
  NOR2_X1 U616 ( .A1(G902), .A2(n729), .ZN(n516) );
  XOR2_X1 U617 ( .A(G475), .B(n516), .Z(n518) );
  INV_X1 U618 ( .A(KEYINPUT13), .ZN(n517) );
  XNOR2_X1 U619 ( .A(n518), .B(n517), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(G107), .Z(n520) );
  XNOR2_X1 U621 ( .A(G116), .B(G122), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n520), .B(n519), .ZN(n525) );
  XOR2_X1 U623 ( .A(KEYINPUT9), .B(KEYINPUT99), .Z(n523) );
  NAND2_X1 U624 ( .A1(G217), .A2(n521), .ZN(n522) );
  XNOR2_X1 U625 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U626 ( .A(n525), .B(n524), .ZN(n527) );
  XNOR2_X1 U627 ( .A(n526), .B(n527), .ZN(n734) );
  NAND2_X1 U628 ( .A1(n734), .A2(n528), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n529), .B(G478), .ZN(n553) );
  AND2_X1 U630 ( .A1(n554), .A2(n553), .ZN(n597) );
  NOR2_X1 U631 ( .A1(n553), .A2(n554), .ZN(n682) );
  NAND2_X1 U632 ( .A1(n682), .A2(n690), .ZN(n532) );
  NOR2_X1 U633 ( .A1(n533), .A2(n699), .ZN(n534) );
  NAND2_X1 U634 ( .A1(n559), .A2(n534), .ZN(n536) );
  INV_X1 U635 ( .A(KEYINPUT65), .ZN(n535) );
  INV_X1 U636 ( .A(KEYINPUT87), .ZN(n537) );
  XNOR2_X1 U637 ( .A(n696), .B(n537), .ZN(n611) );
  NOR2_X1 U638 ( .A1(n611), .A2(n691), .ZN(n538) );
  XNOR2_X1 U639 ( .A(n538), .B(KEYINPUT102), .ZN(n539) );
  INV_X1 U640 ( .A(KEYINPUT83), .ZN(n542) );
  NAND2_X1 U641 ( .A1(KEYINPUT44), .A2(n543), .ZN(n544) );
  NAND2_X1 U642 ( .A1(n545), .A2(n699), .ZN(n703) );
  NOR2_X1 U643 ( .A1(n549), .A2(n703), .ZN(n546) );
  XNOR2_X1 U644 ( .A(n546), .B(KEYINPUT31), .ZN(n662) );
  NAND2_X1 U645 ( .A1(n547), .A2(n582), .ZN(n548) );
  NOR2_X1 U646 ( .A1(n549), .A2(n565), .ZN(n551) );
  NAND2_X1 U647 ( .A1(n551), .A2(n550), .ZN(n646) );
  NAND2_X1 U648 ( .A1(n662), .A2(n646), .ZN(n556) );
  INV_X1 U649 ( .A(n554), .ZN(n552) );
  NAND2_X1 U650 ( .A1(n552), .A2(n553), .ZN(n663) );
  INV_X1 U651 ( .A(n553), .ZN(n555) );
  NAND2_X1 U652 ( .A1(n555), .A2(n554), .ZN(n660) );
  NAND2_X1 U653 ( .A1(n663), .A2(n660), .ZN(n683) );
  NAND2_X1 U654 ( .A1(n556), .A2(n683), .ZN(n561) );
  AND2_X1 U655 ( .A1(n557), .A2(n696), .ZN(n558) );
  AND2_X1 U656 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U657 ( .A(n560), .B(KEYINPUT101), .ZN(n764) );
  AND2_X1 U658 ( .A1(n561), .A2(n764), .ZN(n562) );
  NAND2_X1 U659 ( .A1(KEYINPUT83), .A2(n768), .ZN(n563) );
  NAND2_X1 U660 ( .A1(n699), .A2(n678), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n566), .B(KEYINPUT30), .ZN(n572) );
  NOR2_X1 U662 ( .A1(G900), .A2(n567), .ZN(n568) );
  NAND2_X1 U663 ( .A1(G953), .A2(n568), .ZN(n569) );
  XOR2_X1 U664 ( .A(KEYINPUT104), .B(n569), .Z(n570) );
  NOR2_X1 U665 ( .A1(n571), .A2(n570), .ZN(n580) );
  NOR2_X1 U666 ( .A1(n572), .A2(n580), .ZN(n573) );
  XNOR2_X1 U667 ( .A(KEYINPUT71), .B(KEYINPUT38), .ZN(n575) );
  INV_X1 U668 ( .A(n574), .ZN(n596) );
  INV_X1 U669 ( .A(KEYINPUT39), .ZN(n576) );
  INV_X1 U670 ( .A(n690), .ZN(n579) );
  NAND2_X1 U671 ( .A1(n605), .A2(n699), .ZN(n581) );
  XOR2_X1 U672 ( .A(n581), .B(KEYINPUT28), .Z(n583) );
  NAND2_X1 U673 ( .A1(n583), .A2(n582), .ZN(n588) );
  XOR2_X1 U674 ( .A(KEYINPUT108), .B(KEYINPUT41), .Z(n586) );
  NAND2_X1 U675 ( .A1(n678), .A2(n679), .ZN(n584) );
  NAND2_X1 U676 ( .A1(n684), .A2(n682), .ZN(n585) );
  NOR2_X1 U677 ( .A1(n588), .A2(n707), .ZN(n587) );
  XNOR2_X1 U678 ( .A(n587), .B(KEYINPUT42), .ZN(n769) );
  INV_X1 U679 ( .A(n683), .ZN(n590) );
  NAND2_X1 U680 ( .A1(KEYINPUT76), .A2(n590), .ZN(n591) );
  AND2_X1 U681 ( .A1(KEYINPUT47), .A2(n591), .ZN(n592) );
  NAND2_X1 U682 ( .A1(n657), .A2(n592), .ZN(n595) );
  NAND2_X1 U683 ( .A1(n657), .A2(n683), .ZN(n593) );
  NAND2_X1 U684 ( .A1(n593), .A2(KEYINPUT76), .ZN(n594) );
  INV_X1 U685 ( .A(n596), .ZN(n619) );
  NAND2_X1 U686 ( .A1(n619), .A2(n597), .ZN(n598) );
  NOR2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n656) );
  INV_X1 U688 ( .A(KEYINPUT76), .ZN(n600) );
  AND2_X1 U689 ( .A1(n683), .A2(n600), .ZN(n601) );
  NOR2_X1 U690 ( .A1(n656), .A2(n601), .ZN(n602) );
  AND2_X1 U691 ( .A1(n603), .A2(n602), .ZN(n613) );
  XNOR2_X1 U692 ( .A(n606), .B(KEYINPUT105), .ZN(n607) );
  INV_X1 U693 ( .A(n660), .ZN(n658) );
  AND2_X1 U694 ( .A1(n607), .A2(n658), .ZN(n617) );
  INV_X1 U695 ( .A(n608), .ZN(n609) );
  INV_X1 U696 ( .A(KEYINPUT36), .ZN(n610) );
  INV_X1 U697 ( .A(n611), .ZN(n612) );
  NOR2_X1 U698 ( .A1(n615), .A2(n663), .ZN(n669) );
  AND2_X1 U699 ( .A1(n696), .A2(n678), .ZN(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U701 ( .A(n618), .B(KEYINPUT43), .ZN(n621) );
  INV_X1 U702 ( .A(n619), .ZN(n620) );
  NAND2_X1 U703 ( .A1(n621), .A2(n620), .ZN(n671) );
  INV_X1 U704 ( .A(n671), .ZN(n622) );
  NOR2_X1 U705 ( .A1(n669), .A2(n622), .ZN(n623) );
  INV_X1 U706 ( .A(KEYINPUT81), .ZN(n627) );
  OR2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n624) );
  AND2_X1 U708 ( .A1(n624), .A2(KEYINPUT2), .ZN(n625) );
  NOR2_X1 U709 ( .A1(n628), .A2(KEYINPUT2), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n738), .A2(G472), .ZN(n633) );
  XNOR2_X1 U712 ( .A(KEYINPUT86), .B(KEYINPUT62), .ZN(n630) );
  XNOR2_X1 U713 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U714 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n636), .B(n635), .ZN(G57) );
  NAND2_X1 U716 ( .A1(n738), .A2(G210), .ZN(n640) );
  XNOR2_X1 U717 ( .A(KEYINPUT84), .B(KEYINPUT54), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n638), .B(KEYINPUT55), .ZN(n639) );
  XNOR2_X1 U719 ( .A(n640), .B(n435), .ZN(n642) );
  XNOR2_X1 U720 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n643) );
  XNOR2_X1 U721 ( .A(n644), .B(n643), .ZN(G51) );
  NOR2_X1 U722 ( .A1(n646), .A2(n660), .ZN(n645) );
  XOR2_X1 U723 ( .A(G104), .B(n645), .Z(G6) );
  NOR2_X1 U724 ( .A1(n646), .A2(n663), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U726 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U727 ( .A(G107), .B(n649), .ZN(G9) );
  XNOR2_X1 U728 ( .A(n650), .B(G110), .ZN(n651) );
  XNOR2_X1 U729 ( .A(n651), .B(KEYINPUT109), .ZN(G12) );
  XOR2_X1 U730 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n654) );
  INV_X1 U731 ( .A(n663), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n657), .A2(n652), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U734 ( .A(G128), .B(n655), .ZN(G30) );
  XOR2_X1 U735 ( .A(G143), .B(n656), .Z(G45) );
  NAND2_X1 U736 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U737 ( .A(G146), .B(n659), .ZN(G48) );
  NOR2_X1 U738 ( .A1(n660), .A2(n662), .ZN(n661) );
  XOR2_X1 U739 ( .A(G113), .B(n661), .Z(G15) );
  NOR2_X1 U740 ( .A1(n663), .A2(n662), .ZN(n665) );
  XNOR2_X1 U741 ( .A(G116), .B(KEYINPUT111), .ZN(n664) );
  XNOR2_X1 U742 ( .A(n665), .B(n664), .ZN(G18) );
  XOR2_X1 U743 ( .A(KEYINPUT112), .B(KEYINPUT37), .Z(n666) );
  XNOR2_X1 U744 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U745 ( .A(G125), .B(n668), .ZN(G27) );
  XOR2_X1 U746 ( .A(G134), .B(n669), .Z(G36) );
  XOR2_X1 U747 ( .A(G140), .B(KEYINPUT113), .Z(n670) );
  XNOR2_X1 U748 ( .A(n671), .B(n670), .ZN(G42) );
  INV_X1 U749 ( .A(n672), .ZN(n673) );
  NOR2_X1 U750 ( .A1(n755), .A2(KEYINPUT2), .ZN(n674) );
  XNOR2_X1 U751 ( .A(n674), .B(KEYINPUT80), .ZN(n675) );
  NOR2_X1 U752 ( .A1(n707), .A2(n420), .ZN(n715) );
  NOR2_X1 U753 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U754 ( .A(KEYINPUT118), .B(n680), .Z(n681) );
  NAND2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  NAND2_X1 U758 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U759 ( .A(KEYINPUT119), .B(n689), .ZN(n710) );
  XOR2_X1 U760 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n693) );
  OR2_X1 U761 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U762 ( .A(n693), .B(n692), .ZN(n694) );
  XOR2_X1 U763 ( .A(KEYINPUT114), .B(n694), .Z(n702) );
  XOR2_X1 U764 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n698) );
  NAND2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U766 ( .A(n698), .B(n697), .ZN(n700) );
  NOR2_X1 U767 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n704) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U770 ( .A(KEYINPUT51), .B(n705), .ZN(n706) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U772 ( .A(KEYINPUT117), .B(n708), .Z(n709) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U774 ( .A(n711), .B(KEYINPUT52), .ZN(n712) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  OR2_X1 U776 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U777 ( .A(KEYINPUT53), .B(n721), .ZN(G75) );
  BUF_X1 U778 ( .A(n738), .Z(n722) );
  NAND2_X1 U779 ( .A1(n722), .A2(G469), .ZN(n727) );
  XOR2_X1 U780 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n723) );
  XOR2_X1 U781 ( .A(n723), .B(KEYINPUT121), .Z(n724) );
  XNOR2_X1 U782 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U783 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U784 ( .A1(n742), .A2(n728), .ZN(G54) );
  NAND2_X1 U785 ( .A1(n738), .A2(G475), .ZN(n731) );
  XOR2_X1 U786 ( .A(n729), .B(KEYINPUT59), .Z(n730) );
  XNOR2_X1 U787 ( .A(n731), .B(n730), .ZN(n732) );
  XNOR2_X1 U788 ( .A(n733), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U789 ( .A1(n722), .A2(G478), .ZN(n736) );
  XOR2_X1 U790 ( .A(KEYINPUT122), .B(n734), .Z(n735) );
  XNOR2_X1 U791 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U792 ( .A1(n742), .A2(n737), .ZN(G63) );
  NAND2_X1 U793 ( .A1(n722), .A2(G217), .ZN(n740) );
  XNOR2_X1 U794 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U795 ( .A1(n742), .A2(n741), .ZN(G66) );
  BUF_X1 U796 ( .A(n743), .Z(n744) );
  NAND2_X1 U797 ( .A1(n756), .A2(n744), .ZN(n748) );
  NAND2_X1 U798 ( .A1(G953), .A2(G224), .ZN(n745) );
  XNOR2_X1 U799 ( .A(KEYINPUT61), .B(n745), .ZN(n746) );
  NAND2_X1 U800 ( .A1(n746), .A2(G898), .ZN(n747) );
  NAND2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n753) );
  XOR2_X1 U802 ( .A(n749), .B(KEYINPUT123), .Z(n750) );
  NOR2_X1 U803 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U804 ( .A(n753), .B(n752), .ZN(G69) );
  XNOR2_X1 U805 ( .A(n755), .B(n759), .ZN(n757) );
  NAND2_X1 U806 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U807 ( .A(n758), .B(KEYINPUT124), .ZN(n763) );
  XOR2_X1 U808 ( .A(n759), .B(G227), .Z(n760) );
  NAND2_X1 U809 ( .A1(n760), .A2(G900), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n761), .A2(G953), .ZN(n762) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(G72) );
  XNOR2_X1 U812 ( .A(G101), .B(n764), .ZN(G3) );
  XOR2_X1 U813 ( .A(G119), .B(KEYINPUT126), .Z(n765) );
  XNOR2_X1 U814 ( .A(n766), .B(n765), .ZN(G21) );
  XOR2_X1 U815 ( .A(G122), .B(KEYINPUT125), .Z(n767) );
  XNOR2_X1 U816 ( .A(n768), .B(n767), .ZN(G24) );
  XOR2_X1 U817 ( .A(n769), .B(G137), .Z(G39) );
  XNOR2_X1 U818 ( .A(G131), .B(KEYINPUT127), .ZN(n771) );
  XNOR2_X1 U819 ( .A(n771), .B(n770), .ZN(G33) );
endmodule

