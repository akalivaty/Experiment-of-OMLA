//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n189), .B(new_n191), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(G116), .B(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT5), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(new_n192), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n196), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT75), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G107), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(G107), .ZN(new_n205));
  INV_X1    g019(.A(G107), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT75), .A3(G104), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G101), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(new_n206), .A3(G104), .ZN(new_n212));
  INV_X1    g026(.A(G101), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n205), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n209), .A2(KEYINPUT77), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT77), .B1(new_n209), .B2(new_n214), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n201), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n210), .A2(new_n212), .A3(new_n205), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n189), .A2(new_n191), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT2), .B(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n213), .A2(KEYINPUT4), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n195), .A2(new_n223), .B1(new_n218), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n220), .A2(new_n225), .A3(KEYINPUT80), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT80), .B1(new_n220), .B2(new_n225), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n217), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT6), .ZN(new_n229));
  XNOR2_X1  g043(.A(G110), .B(G122), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n228), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n217), .B(new_n230), .C1(new_n226), .C2(new_n227), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT6), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n220), .A2(new_n225), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT80), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n225), .A3(KEYINPUT80), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n230), .B1(new_n239), .B2(new_n217), .ZN(new_n240));
  OAI211_X1 g054(.A(KEYINPUT81), .B(new_n232), .C1(new_n234), .C2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n228), .A2(new_n231), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT81), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT6), .A4(new_n233), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  XNOR2_X1  g060(.A(G143), .B(G146), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT0), .B(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT64), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n249), .A2(new_n251), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(KEYINPUT82), .A3(G125), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT82), .B1(new_n260), .B2(G125), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT83), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(G125), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n267), .A2(new_n268), .A3(new_n261), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n252), .A2(G143), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n256), .A2(new_n270), .B1(KEYINPUT1), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n247), .A2(new_n274), .A3(G128), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n264), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G224), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT84), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n264), .A2(new_n269), .A3(new_n280), .A4(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n245), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n280), .A2(KEYINPUT7), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n277), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n230), .B(KEYINPUT8), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n198), .A2(KEYINPUT85), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(new_n200), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n198), .A2(KEYINPUT85), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n195), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT77), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT75), .B1(new_n206), .B2(G104), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n206), .A2(G104), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n213), .B1(new_n298), .B2(new_n207), .ZN(new_n299));
  INV_X1    g113(.A(new_n214), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n295), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n209), .A2(KEYINPUT77), .A3(new_n214), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n299), .A2(new_n300), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n201), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n290), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n267), .A2(new_n261), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n276), .B(KEYINPUT86), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n287), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n306), .A2(new_n309), .A3(new_n233), .ZN(new_n310));
  AOI21_X1  g124(.A(G902), .B1(new_n289), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n285), .A2(new_n286), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n286), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n241), .A2(new_n244), .B1(new_n282), .B2(new_n283), .ZN(new_n314));
  INV_X1    g128(.A(G902), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n306), .A2(new_n309), .A3(new_n233), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(new_n288), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n313), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G478), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n320), .A2(KEYINPUT15), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n254), .A2(G128), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT13), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n270), .A2(G143), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n254), .A2(KEYINPUT13), .A3(G128), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AND2_X1   g142(.A1(new_n328), .A2(G134), .ZN(new_n329));
  INV_X1    g143(.A(G134), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n323), .A2(new_n326), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n190), .A2(G122), .ZN(new_n332));
  INV_X1    g146(.A(G122), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G116), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n334), .A3(new_n206), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n206), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n331), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT73), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(G217), .A3(new_n278), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT90), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n346), .B(KEYINPUT14), .C1(new_n333), .C2(G116), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n334), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n332), .B2(KEYINPUT14), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OR2_X1    g164(.A1(new_n332), .A2(KEYINPUT14), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT14), .B1(new_n333), .B2(G116), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT90), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT91), .A3(new_n334), .A4(new_n347), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n351), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(G107), .ZN(new_n356));
  INV_X1    g170(.A(new_n331), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n330), .B1(new_n323), .B2(new_n326), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n335), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n340), .B(new_n344), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n355), .B2(G107), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n343), .B1(new_n361), .B2(new_n339), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n322), .B1(new_n363), .B2(new_n315), .ZN(new_n364));
  AOI211_X1 g178(.A(G902), .B(new_n321), .C1(new_n360), .C2(new_n362), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G140), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G125), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n273), .A2(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT71), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n367), .A2(KEYINPUT71), .A3(G125), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT16), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n372), .A2(new_n252), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n252), .B1(new_n372), .B2(new_n374), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(G237), .A2(G953), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(G143), .A3(G214), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n378), .B2(G214), .ZN(new_n381));
  OAI21_X1  g195(.A(G131), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT88), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT17), .ZN(new_n385));
  INV_X1    g199(.A(G237), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(new_n278), .A3(G214), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n254), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n379), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT88), .A3(G131), .ZN(new_n390));
  INV_X1    g204(.A(G131), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n391), .A3(new_n379), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n384), .A2(new_n385), .A3(new_n390), .A4(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT88), .B1(new_n389), .B2(G131), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n383), .B(new_n391), .C1(new_n388), .C2(new_n379), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT17), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n377), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n370), .A2(new_n371), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT87), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n370), .A2(new_n371), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(G146), .A3(new_n401), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n368), .A2(new_n369), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n252), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(KEYINPUT18), .A2(G131), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n388), .A2(new_n379), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n389), .A2(KEYINPUT18), .A3(G131), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n203), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n397), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n397), .B2(new_n409), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n315), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(G475), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n407), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n404), .B2(new_n402), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n394), .A2(new_n395), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n376), .B1(new_n419), .B2(new_n392), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n399), .A2(KEYINPUT19), .A3(new_n401), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n403), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n252), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n418), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n412), .B1(new_n425), .B2(new_n411), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT20), .ZN(new_n427));
  NOR2_X1   g241(.A1(G475), .A2(G902), .ZN(new_n428));
  XOR2_X1   g242(.A(new_n428), .B(KEYINPUT89), .Z(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n426), .B2(new_n429), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n366), .B(new_n416), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n278), .A2(G952), .ZN(new_n434));
  INV_X1    g248(.A(G234), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n434), .B1(new_n435), .B2(new_n386), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI211_X1 g251(.A(new_n315), .B(new_n278), .C1(G234), .C2(G237), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G898), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n433), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G214), .B1(G237), .B2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n319), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n275), .A2(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n272), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n275), .A2(KEYINPUT76), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n304), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT10), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n272), .A2(new_n275), .ZN(new_n450));
  OAI211_X1 g264(.A(KEYINPUT10), .B(new_n450), .C1(new_n215), .C2(new_n216), .ZN(new_n451));
  INV_X1    g265(.A(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT65), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G137), .ZN(new_n455));
  AND2_X1   g269(.A1(KEYINPUT11), .A2(G134), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(KEYINPUT11), .A2(G134), .ZN(new_n458));
  NOR2_X1   g272(.A1(KEYINPUT11), .A2(G134), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n458), .B1(new_n459), .B2(G137), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n457), .A2(new_n391), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n391), .B1(new_n457), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n249), .A2(new_n251), .A3(new_n259), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n218), .A2(new_n224), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n220), .A3(new_n465), .ZN(new_n466));
  NAND4_X1  g280(.A1(new_n449), .A2(new_n451), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n278), .A2(G227), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n468), .B(KEYINPUT74), .ZN(new_n469));
  XNOR2_X1  g283(.A(G110), .B(G140), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n467), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT79), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n467), .A2(KEYINPUT79), .A3(new_n472), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n449), .A2(new_n451), .A3(new_n466), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n457), .A2(new_n460), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G131), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n457), .A2(new_n391), .A3(new_n460), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n475), .A2(new_n476), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n467), .ZN(new_n484));
  INV_X1    g298(.A(new_n450), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n301), .A2(new_n485), .A3(new_n302), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT78), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n301), .A2(new_n485), .A3(new_n488), .A4(new_n302), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n489), .A3(new_n447), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n481), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT12), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(KEYINPUT12), .A3(new_n481), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n484), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(G469), .B(new_n483), .C1(new_n495), .C2(new_n472), .ZN(new_n496));
  INV_X1    g310(.A(G469), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n473), .B1(new_n493), .B2(new_n494), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n472), .B1(new_n482), .B2(new_n467), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n497), .B(new_n315), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n497), .A2(new_n315), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G221), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n342), .B2(new_n315), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n187), .B1(new_n443), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n188), .B2(G128), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n270), .A2(KEYINPUT23), .A3(G119), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n510), .B(new_n511), .C1(G119), .C2(new_n270), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G110), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT24), .B(G110), .Z(new_n514));
  XNOR2_X1  g328(.A(G119), .B(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n377), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n376), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n512), .A2(G110), .B1(new_n515), .B2(new_n514), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n404), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G137), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n504), .A2(new_n435), .A3(G953), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  NAND3_X1  g338(.A1(new_n518), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n524), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n377), .A2(new_n517), .ZN(new_n527));
  INV_X1    g341(.A(new_n521), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n525), .A2(new_n529), .A3(new_n315), .ZN(new_n530));
  NOR2_X1   g344(.A1(KEYINPUT72), .A2(KEYINPUT25), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n525), .A2(new_n529), .A3(new_n315), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G217), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(G234), .B2(new_n315), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n525), .A2(new_n529), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(G902), .ZN(new_n539));
  AOI22_X1  g353(.A1(new_n535), .A2(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT28), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n464), .A2(new_n481), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n453), .A2(new_n455), .A3(new_n330), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n544), .B(G131), .C1(new_n330), .C2(new_n452), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n450), .A2(new_n480), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n195), .A2(new_n223), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n542), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n548), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n463), .A2(new_n260), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT66), .B1(new_n464), .B2(new_n481), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n551), .B(new_n546), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n547), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n555), .B1(new_n551), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n558));
  AOI21_X1  g372(.A(new_n550), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n378), .A2(G210), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT27), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n563), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n450), .A2(new_n480), .A3(new_n545), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n552), .B1(new_n463), .B2(new_n260), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n464), .A2(new_n481), .A3(KEYINPUT66), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AOI211_X1 g384(.A(KEYINPUT68), .B(new_n566), .C1(new_n570), .C2(new_n551), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT68), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n555), .B2(new_n563), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT30), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n547), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n548), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT67), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n546), .B1(new_n553), .B2(new_n554), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n575), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n570), .A2(KEYINPUT67), .A3(KEYINPUT30), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n577), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT31), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n574), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(new_n548), .B(new_n567), .C1(new_n568), .C2(new_n569), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT68), .B1(new_n585), .B2(new_n566), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n555), .A2(new_n572), .A3(new_n563), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n577), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n568), .A2(new_n569), .ZN(new_n590));
  AND4_X1   g404(.A1(KEYINPUT67), .A2(new_n590), .A3(KEYINPUT30), .A4(new_n546), .ZN(new_n591));
  AOI21_X1  g405(.A(KEYINPUT67), .B1(new_n570), .B2(KEYINPUT30), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT31), .B1(new_n588), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n565), .B1(new_n584), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(G472), .A2(G902), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT32), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n570), .A2(new_n551), .ZN(new_n600));
  OAI21_X1  g414(.A(KEYINPUT28), .B1(new_n600), .B2(new_n585), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n601), .A2(KEYINPUT29), .A3(new_n563), .A4(new_n549), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n563), .B1(new_n593), .B2(new_n555), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT29), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n551), .B1(new_n543), .B2(new_n546), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n570), .B2(new_n551), .ZN(new_n606));
  INV_X1    g420(.A(new_n558), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n549), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n604), .B1(new_n608), .B2(new_n566), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n315), .B(new_n602), .C1(new_n603), .C2(new_n609), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n595), .A2(new_n599), .B1(new_n610), .B2(G472), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n583), .B1(new_n574), .B2(new_n582), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n588), .A2(KEYINPUT31), .A3(new_n593), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n564), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n613), .B1(new_n616), .B2(new_n597), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n541), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n473), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n490), .A2(KEYINPUT12), .A3(new_n481), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT12), .B1(new_n490), .B2(new_n481), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n499), .ZN(new_n623));
  AOI21_X1  g437(.A(G902), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n501), .B1(new_n624), .B2(new_n497), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n505), .B1(new_n625), .B2(new_n496), .ZN(new_n626));
  INV_X1    g440(.A(new_n442), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n312), .B2(new_n318), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n626), .A2(KEYINPUT92), .A3(new_n628), .A4(new_n441), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n508), .A2(new_n618), .A3(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G101), .ZN(G3));
  OAI21_X1  g445(.A(G472), .B1(new_n616), .B2(G902), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n595), .A2(new_n596), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n635), .A2(new_n541), .A3(new_n507), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n320), .A2(G902), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n360), .A2(new_n638), .A3(new_n362), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n638), .B1(new_n360), .B2(new_n362), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT94), .ZN(new_n643));
  AOI21_X1  g457(.A(G478), .B1(new_n363), .B2(new_n315), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n637), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n363), .A2(KEYINPUT33), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(new_n639), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT94), .B1(new_n649), .B2(new_n644), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n426), .A2(new_n429), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT20), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n430), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n646), .A2(new_n650), .B1(new_n653), .B2(new_n416), .ZN(new_n654));
  INV_X1    g468(.A(new_n440), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n286), .B1(new_n285), .B2(new_n311), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n314), .A2(new_n317), .A3(new_n313), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n442), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(KEYINPUT93), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT93), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n628), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n656), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n636), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT34), .B(G104), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G6));
  OR2_X1    g480(.A1(new_n364), .A2(new_n365), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n667), .B(new_n416), .C1(new_n432), .C2(new_n431), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n655), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n660), .B2(new_n662), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n636), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT35), .B(G107), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G9));
  NAND2_X1  g488(.A1(new_n518), .A2(new_n521), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT95), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n527), .A2(new_n528), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT95), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n680), .B1(KEYINPUT36), .B2(new_n526), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n526), .A2(KEYINPUT36), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n676), .A2(new_n682), .A3(new_n679), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n539), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n535), .A2(new_n537), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n632), .A2(new_n633), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n508), .A2(new_n629), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  NAND2_X1  g504(.A1(new_n660), .A2(new_n662), .ZN(new_n691));
  INV_X1    g505(.A(new_n686), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n611), .B2(new_n617), .ZN(new_n693));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n438), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n436), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n668), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n691), .A2(new_n693), .A3(new_n626), .A4(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  INV_X1    g514(.A(KEYINPUT96), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n612), .B1(new_n595), .B2(new_n596), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n579), .A2(new_n548), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n563), .B1(new_n703), .B2(new_n555), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n588), .B2(new_n593), .ZN(new_n705));
  OAI21_X1  g519(.A(G472), .B1(new_n705), .B2(G902), .ZN(new_n706));
  INV_X1    g520(.A(new_n599), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n706), .B1(new_n616), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n701), .B1(new_n702), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n595), .A2(new_n599), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n617), .A2(new_n710), .A3(KEYINPUT96), .A4(new_n706), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n319), .B(KEYINPUT38), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n416), .B1(new_n431), .B2(new_n432), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n667), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n715), .A2(new_n686), .A3(new_n627), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n712), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(new_n696), .B(KEYINPUT39), .Z(new_n718));
  NOR2_X1   g532(.A1(new_n507), .A2(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n720), .A2(KEYINPUT40), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(KEYINPUT40), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n717), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT97), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  NOR3_X1   g539(.A1(new_n649), .A2(KEYINPUT94), .A3(new_n644), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n643), .B1(new_n642), .B2(new_n645), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n714), .B(new_n696), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT98), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n650), .A2(new_n646), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT98), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n730), .A2(new_n731), .A3(new_n714), .A4(new_n696), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n691), .A2(new_n693), .A3(new_n733), .A4(new_n626), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  INV_X1    g549(.A(KEYINPUT99), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n624), .A2(new_n497), .ZN(new_n737));
  AOI211_X1 g551(.A(G469), .B(G902), .C1(new_n622), .C2(new_n623), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n505), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n663), .A2(new_n736), .A3(new_n618), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n656), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n628), .A2(new_n661), .ZN(new_n742));
  AOI211_X1 g556(.A(KEYINPUT93), .B(new_n627), .C1(new_n312), .C2(new_n318), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n602), .A2(new_n315), .ZN(new_n745));
  INV_X1    g559(.A(new_n603), .ZN(new_n746));
  INV_X1    g560(.A(new_n609), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(G472), .ZN(new_n749));
  OAI22_X1  g563(.A1(new_n748), .A2(new_n749), .B1(new_n616), .B2(new_n707), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n540), .B(new_n739), .C1(new_n750), .C2(new_n702), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT99), .B1(new_n744), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n740), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND3_X1  g569(.A1(new_n671), .A2(new_n618), .A3(new_n739), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NAND4_X1  g571(.A1(new_n691), .A2(new_n693), .A3(new_n441), .A4(new_n739), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  INV_X1    g573(.A(KEYINPUT100), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n542), .B1(new_n703), .B2(new_n555), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n760), .B1(new_n761), .B2(new_n550), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n601), .A2(KEYINPUT100), .A3(new_n549), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(new_n566), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n584), .B2(new_n594), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n596), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n632), .A2(new_n766), .A3(new_n540), .ZN(new_n767));
  INV_X1    g581(.A(new_n715), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n622), .A2(new_n623), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n315), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(G469), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n506), .A3(new_n500), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n440), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n691), .A2(new_n767), .A3(new_n768), .A4(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G122), .ZN(G24));
  NAND2_X1  g589(.A1(new_n729), .A2(new_n732), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n632), .A2(new_n766), .A3(new_n686), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n772), .B1(new_n660), .B2(new_n662), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G125), .ZN(G27));
  NAND3_X1  g595(.A1(new_n312), .A2(new_n318), .A3(new_n442), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT102), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n501), .B(KEYINPUT101), .Z(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(new_n624), .B2(new_n497), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n505), .B1(new_n786), .B2(new_n496), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT102), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n312), .A2(new_n318), .A3(new_n788), .A4(new_n442), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n783), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(new_n618), .A3(new_n733), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT42), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT103), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n598), .B1(new_n616), .B2(new_n597), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n610), .A2(G472), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n710), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n496), .A2(new_n500), .A3(new_n784), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(KEYINPUT42), .A3(new_n506), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n797), .A2(new_n799), .A3(new_n540), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n783), .A2(new_n729), .A3(new_n732), .A4(new_n789), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n794), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n799), .A3(new_n540), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n801), .A3(KEYINPUT103), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n793), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G131), .ZN(G33));
  NAND3_X1  g621(.A1(new_n790), .A2(new_n618), .A3(new_n698), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G134), .ZN(G36));
  OAI21_X1  g623(.A(new_n483), .B1(new_n495), .B2(new_n472), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT45), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n813), .A3(new_n497), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n785), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT46), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n500), .B1(new_n815), .B2(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n506), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n718), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n783), .A2(new_n789), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n726), .A2(new_n727), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n823), .A2(KEYINPUT43), .A3(new_n714), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT43), .B1(new_n823), .B2(new_n714), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n635), .A3(new_n686), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n822), .B1(new_n828), .B2(KEYINPUT44), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n820), .B(new_n829), .C1(KEYINPUT44), .C2(new_n828), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  XNOR2_X1  g645(.A(KEYINPUT104), .B(KEYINPUT47), .ZN(new_n832));
  XOR2_X1   g646(.A(new_n819), .B(new_n832), .Z(new_n833));
  NAND4_X1  g647(.A1(new_n802), .A2(new_n611), .A3(new_n617), .A4(new_n541), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT105), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  NAND2_X1  g651(.A1(new_n826), .A2(new_n437), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT115), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n826), .A2(new_n840), .A3(new_n437), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n541), .B1(new_n611), .B2(new_n795), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n822), .A2(new_n772), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT48), .Z(new_n846));
  INV_X1    g660(.A(KEYINPUT118), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n842), .A2(new_n767), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(new_n779), .ZN(new_n849));
  INV_X1    g663(.A(new_n654), .ZN(new_n850));
  INV_X1    g664(.A(new_n712), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n541), .A2(new_n436), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n844), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n849), .B(new_n434), .C1(new_n850), .C2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n846), .B1(new_n847), .B2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n737), .A2(new_n738), .A3(new_n506), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n833), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n821), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT51), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n853), .A2(new_n714), .A3(new_n730), .ZN(new_n860));
  INV_X1    g674(.A(new_n777), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n842), .A2(new_n844), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n739), .A2(new_n627), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n865), .A2(new_n866), .A3(new_n713), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n848), .A2(KEYINPUT50), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT50), .B1(new_n848), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI221_X1 g684(.A(new_n855), .B1(new_n847), .B2(new_n854), .C1(new_n859), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT117), .ZN(new_n873));
  OR2_X1    g687(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n874), .B(new_n875), .C1(new_n857), .C2(new_n858), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n871), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n756), .A2(new_n758), .A3(new_n774), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n740), .B2(new_n752), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT114), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n715), .B1(new_n660), .B2(new_n662), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n798), .A2(new_n506), .ZN(new_n883));
  OR3_X1    g697(.A1(new_n686), .A2(KEYINPUT109), .A3(new_n697), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT109), .B1(new_n686), .B2(new_n697), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n712), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n887), .A2(new_n699), .A3(new_n780), .A4(new_n734), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT110), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n626), .B(new_n686), .C1(new_n750), .C2(new_n702), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n891), .B(new_n691), .C1(new_n698), .C2(new_n733), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT110), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n893), .A3(new_n780), .A4(new_n887), .ZN(new_n894));
  XNOR2_X1  g708(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n889), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n888), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n778), .A2(new_n790), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n433), .A2(new_n697), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n821), .A2(new_n693), .A3(new_n626), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n808), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n800), .A2(new_n794), .A3(new_n802), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT103), .B1(new_n804), .B2(new_n801), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n902), .B1(new_n905), .B2(new_n793), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n319), .A2(new_n442), .A3(new_n655), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n654), .A2(new_n669), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n634), .A3(new_n540), .A4(new_n626), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n630), .A2(new_n688), .A3(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n906), .A2(KEYINPUT53), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n881), .A2(new_n898), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT108), .ZN(new_n914));
  INV_X1    g728(.A(new_n902), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n806), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n751), .ZN(new_n917));
  INV_X1    g731(.A(new_n441), .ZN(new_n918));
  AOI211_X1 g732(.A(new_n692), .B(new_n918), .C1(new_n611), .C2(new_n617), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n917), .A2(new_n671), .B1(new_n919), .B2(new_n779), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n911), .A2(new_n753), .A3(new_n774), .A4(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n914), .B1(new_n916), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n906), .A2(new_n880), .A3(KEYINPUT108), .A4(new_n911), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n889), .A2(new_n897), .A3(new_n894), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n897), .B1(new_n889), .B2(new_n894), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT113), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT53), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n878), .B(new_n913), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n926), .A2(KEYINPUT53), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n898), .A2(new_n922), .A3(new_n923), .A4(new_n928), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n933), .A2(KEYINPUT54), .A3(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT112), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n933), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n877), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(G952), .B2(G953), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n540), .A2(new_n506), .A3(new_n442), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n942), .A2(new_n714), .A3(new_n823), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT49), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n737), .A2(new_n738), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT106), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n713), .B1(new_n944), .B2(new_n945), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n851), .A3(new_n948), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT107), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n941), .A2(new_n950), .ZN(G75));
  NOR2_X1   g765(.A1(new_n278), .A2(G952), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n926), .A2(new_n928), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(KEYINPUT113), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n955), .A2(new_n929), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n315), .B1(new_n956), .B2(new_n913), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(G210), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n245), .A2(new_n284), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n960), .A2(new_n314), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT55), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(KEYINPUT120), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(KEYINPUT120), .ZN(new_n964));
  XOR2_X1   g778(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n953), .B1(new_n959), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT56), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n958), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n967), .A2(new_n969), .ZN(G51));
  XOR2_X1   g784(.A(new_n784), .B(KEYINPUT57), .Z(new_n971));
  INV_X1    g785(.A(new_n932), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n878), .B1(new_n956), .B2(new_n913), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n769), .B(KEYINPUT121), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n814), .B(KEYINPUT122), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n957), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n952), .B1(new_n976), .B2(new_n978), .ZN(G54));
  NAND2_X1  g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT123), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n957), .A2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(new_n426), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n426), .B1(new_n957), .B2(new_n981), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n952), .A3(new_n985), .ZN(G60));
  NAND2_X1  g800(.A1(G478), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT59), .Z(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n939), .B2(new_n932), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n648), .A2(new_n639), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n953), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n648), .B2(new_n639), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n972), .B2(new_n973), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT124), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  OAI211_X1 g809(.A(KEYINPUT124), .B(new_n992), .C1(new_n972), .C2(new_n973), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n991), .B1(new_n995), .B2(new_n996), .ZN(G63));
  NAND2_X1  g811(.A1(new_n956), .A2(new_n913), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n681), .A2(new_n683), .ZN(new_n999));
  NAND2_X1  g813(.A1(G217), .A2(G902), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n1000), .B(KEYINPUT60), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n956), .B2(new_n913), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n1003), .B(new_n953), .C1(new_n538), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1004), .A2(new_n538), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n953), .A4(new_n1003), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(G66));
  XOR2_X1   g824(.A(new_n921), .B(KEYINPUT125), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n278), .ZN(new_n1012));
  INV_X1    g826(.A(G224), .ZN(new_n1013));
  OAI21_X1  g827(.A(G953), .B1(new_n439), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n241), .B(new_n244), .C1(G898), .C2(new_n278), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT126), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1015), .B(new_n1017), .ZN(G69));
  OAI21_X1  g832(.A(new_n576), .B1(new_n591), .B2(new_n592), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n421), .A2(new_n423), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(new_n1021));
  INV_X1    g835(.A(new_n908), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n821), .A2(new_n618), .A3(new_n719), .A4(new_n1022), .ZN(new_n1023));
  AND3_X1   g837(.A1(new_n836), .A2(new_n830), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n892), .A2(new_n780), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n724), .A2(new_n1026), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(KEYINPUT62), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1024), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1021), .B1(new_n1030), .B2(new_n278), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n1026), .A2(new_n808), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1032), .A2(new_n806), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n820), .A2(new_n882), .A3(new_n843), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1033), .A2(new_n836), .A3(new_n830), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1035), .A2(G953), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1021), .B1(new_n694), .B2(new_n278), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n1031), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n1040));
  XOR2_X1   g854(.A(new_n1039), .B(new_n1040), .Z(G72));
  NAND2_X1  g855(.A1(new_n593), .A2(new_n555), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1042), .A2(new_n563), .ZN(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  OAI21_X1  g859(.A(new_n1045), .B1(new_n1030), .B2(new_n1011), .ZN(new_n1046));
  OR2_X1    g860(.A1(new_n1046), .A2(KEYINPUT127), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1046), .A2(KEYINPUT127), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1043), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1045), .B1(new_n1035), .B2(new_n1011), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1042), .A2(new_n563), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n952), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n933), .A2(new_n934), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n588), .A2(new_n593), .ZN(new_n1054));
  INV_X1    g868(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1045), .B1(new_n1055), .B2(new_n603), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1052), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g871(.A1(new_n1049), .A2(new_n1057), .ZN(G57));
endmodule


