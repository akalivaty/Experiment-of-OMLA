//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n552, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n587, new_n588, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n632, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1198, new_n1199, new_n1200, new_n1201;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  OAI21_X1  g034(.A(KEYINPUT69), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(new_n462), .A3(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n465));
  AND3_X1   g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  AND2_X1   g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n465), .A2(new_n469), .A3(G125), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n465), .A2(new_n469), .A3(KEYINPUT68), .A4(G125), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n462), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n460), .B2(new_n463), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n458), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n480), .A2(new_n458), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT70), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n483), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n458), .A2(G102), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n480), .B2(G126), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n492), .B1(new_n495), .B2(new_n458), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n464), .A2(new_n458), .A3(new_n465), .A4(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n465), .A2(new_n469), .A3(G138), .A4(new_n458), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n496), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  OAI21_X1  g081(.A(KEYINPUT71), .B1(new_n506), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(new_n504), .A3(KEYINPUT5), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(G543), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n510), .A2(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n510), .A2(new_n520), .A3(G62), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n516), .B1(new_n522), .B2(G651), .ZN(G166));
  AND2_X1   g098(.A1(G76), .A2(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT7), .B1(new_n524), .B2(G651), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n511), .A2(G543), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT73), .B(G51), .Z(new_n527));
  AOI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G89), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n528), .B1(new_n529), .B2(new_n512), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n510), .A2(G63), .B1(KEYINPUT7), .B2(new_n524), .ZN(new_n531));
  INV_X1    g106(.A(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n530), .A2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n532), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  INV_X1    g113(.A(G52), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n512), .A2(new_n538), .B1(new_n539), .B2(new_n515), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n537), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n532), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  INV_X1    g120(.A(G43), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n512), .A2(new_n545), .B1(new_n546), .B2(new_n515), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(G188));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n515), .B2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n511), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n560), .B1(new_n559), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n507), .A2(new_n509), .ZN(new_n565));
  INV_X1    g140(.A(new_n505), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n565), .A2(G65), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT78), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(KEYINPUT78), .A3(new_n568), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n570), .A2(G651), .A3(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(KEYINPUT77), .B1(new_n512), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n510), .A2(new_n575), .A3(G91), .A4(new_n511), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n564), .A2(new_n572), .A3(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n567), .A2(KEYINPUT78), .A3(new_n568), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n569), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n577), .B1(new_n583), .B2(G651), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n584), .A2(KEYINPUT79), .A3(new_n564), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n581), .A2(new_n585), .ZN(G299));
  NAND2_X1  g161(.A1(new_n522), .A2(G651), .ZN(new_n587));
  INV_X1    g162(.A(new_n516), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(G303));
  NAND2_X1  g164(.A1(new_n526), .A2(G49), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT80), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n510), .A2(new_n511), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G87), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(G288));
  AOI21_X1  g170(.A(new_n508), .B1(KEYINPUT5), .B2(new_n504), .ZN(new_n596));
  NOR3_X1   g171(.A1(new_n506), .A2(KEYINPUT71), .A3(G543), .ZN(new_n597));
  OAI211_X1 g172(.A(G61), .B(new_n566), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n532), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND2_X1   g175(.A1(KEYINPUT6), .A2(G651), .ZN(new_n601));
  NOR2_X1   g176(.A1(KEYINPUT6), .A2(G651), .ZN(new_n602));
  OAI211_X1 g177(.A(G48), .B(G543), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g180(.A1(new_n511), .A2(KEYINPUT82), .A3(G48), .A4(G543), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g183(.A1(new_n565), .A2(G86), .A3(new_n566), .A4(new_n511), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g186(.A1(new_n510), .A2(KEYINPUT81), .A3(G86), .A4(new_n511), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n608), .A2(new_n613), .ZN(G305));
  AOI22_X1  g189(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n532), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT83), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n592), .A2(G85), .B1(G47), .B2(new_n526), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(G290));
  NAND2_X1  g194(.A1(G301), .A2(G868), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT10), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n592), .A2(new_n621), .A3(G92), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  OAI21_X1  g198(.A(KEYINPUT10), .B1(new_n512), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n526), .A2(G54), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n510), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n532), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n620), .B1(G868), .B2(new_n629), .ZN(G284));
  OAI21_X1  g205(.A(new_n620), .B1(G868), .B2(new_n629), .ZN(G321));
  NAND2_X1  g206(.A1(G286), .A2(G868), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n581), .A2(new_n585), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G297));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(G868), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n629), .B1(new_n636), .B2(G860), .ZN(G148));
  OAI21_X1  g212(.A(KEYINPUT84), .B1(new_n549), .B2(G868), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(new_n636), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  MUX2_X1   g215(.A(KEYINPUT84), .B(new_n638), .S(new_n640), .Z(G323));
  XOR2_X1   g216(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n642));
  XNOR2_X1  g217(.A(G323), .B(new_n642), .ZN(G282));
  INV_X1    g218(.A(G135), .ZN(new_n644));
  OR3_X1    g219(.A1(new_n484), .A2(KEYINPUT87), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n482), .A2(G123), .ZN(new_n646));
  OR2_X1    g221(.A1(G99), .A2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n647), .B(G2104), .C1(G111), .C2(new_n458), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT87), .B1(new_n484), .B2(new_n644), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n645), .A2(new_n646), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT88), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n458), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT13), .ZN(new_n659));
  INV_X1    g234(.A(G2100), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n655), .A2(new_n661), .ZN(G156));
  XNOR2_X1  g237(.A(KEYINPUT15), .B(G2435), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT90), .B(G2438), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2427), .B(G2430), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n667), .A2(KEYINPUT14), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT89), .B(KEYINPUT16), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2451), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n668), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2443), .B(G2446), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1341), .B(G1348), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(G14), .ZN(G401));
  XOR2_X1   g252(.A(G2067), .B(G2678), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT91), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT18), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n680), .B(KEYINPUT17), .ZN(new_n686));
  OAI211_X1 g261(.A(new_n685), .B(new_n682), .C1(new_n679), .C2(new_n686), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n679), .A2(new_n686), .A3(new_n681), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G2096), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(new_n660), .ZN(G227));
  XOR2_X1   g266(.A(G1956), .B(G2474), .Z(new_n692));
  XOR2_X1   g267(.A(G1961), .B(G1966), .Z(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT19), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n692), .A2(new_n693), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n698), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n702), .B(new_n703), .C1(new_n701), .C2(new_n700), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT92), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n708), .B(new_n710), .ZN(G229));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G26), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT28), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n482), .A2(G128), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n485), .A2(G140), .ZN(new_n716));
  OR2_X1    g291(.A1(G104), .A2(G2105), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n717), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G29), .ZN(new_n720));
  AND2_X1   g295(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n714), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(G2067), .ZN(new_n724));
  INV_X1    g299(.A(new_n654), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(G29), .B2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n712), .A2(G33), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n465), .A2(new_n469), .A3(G127), .ZN(new_n728));
  INV_X1    g303(.A(G115), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n728), .B1(new_n729), .B2(new_n459), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n485), .A2(G139), .B1(G2105), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT25), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n727), .B1(new_n734), .B2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(KEYINPUT96), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n738), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n712), .A2(G27), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G164), .B2(new_n712), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n743), .A2(G2078), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n735), .A2(new_n736), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n746), .A2(G34), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G34), .ZN(new_n748));
  AOI21_X1  g323(.A(G29), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n477), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT30), .B(G28), .Z(new_n752));
  OAI22_X1  g327(.A1(new_n750), .A2(new_n751), .B1(G29), .B2(new_n752), .ZN(new_n753));
  NOR4_X1   g328(.A1(new_n741), .A2(new_n744), .A3(new_n745), .A4(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G16), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n755), .A2(KEYINPUT23), .A3(G20), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT23), .ZN(new_n757));
  INV_X1    g332(.A(G20), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G16), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n759), .C1(new_n633), .C2(new_n755), .ZN(new_n760));
  INV_X1    g335(.A(G1956), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(G168), .A2(G16), .ZN(new_n763));
  OR2_X1    g338(.A1(G16), .A2(G21), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n763), .A2(G1966), .A3(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G1961), .ZN(new_n766));
  OR2_X1    g341(.A1(G5), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G301), .B2(new_n755), .ZN(new_n768));
  OR2_X1    g343(.A1(G29), .A2(G32), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n482), .A2(G129), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n485), .A2(G141), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n458), .A2(G105), .A3(G2104), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT26), .Z(new_n774));
  NAND4_X1  g349(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n769), .B1(new_n775), .B2(new_n712), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT27), .B(G1996), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n766), .A2(new_n768), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n750), .A2(new_n751), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n765), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(G1966), .B1(new_n763), .B2(new_n764), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n768), .A2(new_n766), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n743), .A2(G2078), .ZN(new_n784));
  NOR4_X1   g359(.A1(new_n781), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n726), .A2(new_n754), .A3(new_n762), .A4(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n755), .A2(G23), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G288), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT33), .B(G1976), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT94), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n789), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n755), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n755), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n755), .A2(G6), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G305), .B2(G16), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT32), .B(G1981), .Z(new_n800));
  XOR2_X1   g375(.A(new_n799), .B(new_n800), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n793), .A2(new_n797), .A3(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n793), .A2(new_n803), .A3(new_n797), .A4(new_n801), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(G290), .A2(G16), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n755), .A2(G24), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n810), .A2(G1986), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n810), .A2(G1986), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n482), .A2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n485), .A2(G131), .ZN(new_n814));
  OR2_X1    g389(.A1(G95), .A2(G2105), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n815), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  MUX2_X1   g392(.A(G25), .B(new_n817), .S(G29), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT35), .B(G1991), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n811), .A2(new_n812), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n787), .B1(new_n807), .B2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n807), .A2(new_n787), .A3(new_n821), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n786), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n712), .A2(G35), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G162), .B2(new_n712), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT29), .B(G2090), .Z(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n755), .A2(G4), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n629), .B2(new_n755), .ZN(new_n832));
  INV_X1    g407(.A(G1348), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G19), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n549), .B2(G16), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(G1341), .Z(new_n837));
  NAND4_X1  g412(.A1(new_n825), .A2(new_n830), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n838), .A2(KEYINPUT98), .ZN(new_n840));
  INV_X1    g415(.A(new_n786), .ZN(new_n841));
  INV_X1    g416(.A(new_n824), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n841), .B(new_n837), .C1(new_n842), .C2(new_n822), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n830), .A4(new_n834), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(new_n846), .ZN(G150));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  INV_X1    g423(.A(G55), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n512), .A2(new_n848), .B1(new_n849), .B2(new_n515), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT100), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(KEYINPUT100), .ZN(new_n852));
  AOI22_X1  g427(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n851), .A2(new_n852), .B1(new_n532), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n549), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n854), .A2(new_n548), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n629), .A2(G559), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n857), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n863), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n865), .B(new_n866), .C1(new_n862), .C2(new_n861), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT102), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n854), .A2(G860), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(KEYINPUT37), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(G145));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n654), .B(new_n477), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n490), .ZN(new_n874));
  INV_X1    g449(.A(new_n492), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n461), .B1(new_n462), .B2(G2104), .ZN(new_n876));
  NOR3_X1   g451(.A1(new_n459), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n877));
  OAI211_X1 g452(.A(G126), .B(new_n465), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(new_n493), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n875), .B1(new_n879), .B2(G2105), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n498), .A2(KEYINPUT103), .A3(new_n501), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT103), .B1(new_n498), .B2(new_n501), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n719), .ZN(new_n884));
  INV_X1    g459(.A(new_n775), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n734), .A2(KEYINPUT104), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n884), .B(new_n775), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n887), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n817), .B(new_n658), .ZN(new_n892));
  INV_X1    g467(.A(G142), .ZN(new_n893));
  NOR2_X1   g468(.A1(G106), .A2(G2105), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(new_n458), .B2(G118), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n484), .A2(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(G130), .B2(new_n482), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n892), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n889), .A2(new_n891), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n874), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n899), .B1(new_n889), .B2(new_n891), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n889), .A2(new_n891), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n898), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n889), .A2(new_n891), .A3(new_n904), .A4(new_n898), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI221_X1 g483(.A(new_n872), .B1(new_n901), .B2(new_n902), .C1(new_n874), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g485(.A1(new_n854), .A2(G868), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G288), .B(G303), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(G305), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(G305), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(G290), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n914), .A2(new_n618), .A3(new_n617), .A4(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n857), .B(new_n639), .ZN(new_n922));
  INV_X1    g497(.A(new_n629), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n633), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n629), .B1(new_n581), .B2(new_n585), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G299), .A2(new_n629), .ZN(new_n928));
  INV_X1    g503(.A(new_n925), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT41), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n924), .A2(new_n931), .A3(new_n925), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n922), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n927), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n927), .A2(KEYINPUT107), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n921), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(new_n936), .B2(new_n921), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n912), .B1(new_n939), .B2(G868), .ZN(G295));
  AOI21_X1  g515(.A(new_n912), .B1(new_n939), .B2(G868), .ZN(G331));
  XNOR2_X1  g516(.A(G286), .B(G301), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n857), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n855), .A3(new_n856), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n930), .B2(new_n932), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n944), .B(new_n945), .C1(new_n925), .C2(new_n924), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g524(.A1(new_n917), .A2(new_n918), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n919), .A2(new_n947), .A3(new_n948), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n872), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n951), .A2(new_n952), .A3(new_n956), .A4(new_n872), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n953), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n954), .A2(KEYINPUT44), .A3(new_n957), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(G397));
  NAND3_X1  g538(.A1(new_n468), .A2(new_n476), .A3(G40), .ZN(new_n964));
  INV_X1    g539(.A(G1384), .ZN(new_n965));
  AOI211_X1 g540(.A(KEYINPUT45), .B(new_n964), .C1(new_n883), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(G290), .A2(G1986), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n967), .B1(new_n968), .B2(KEYINPUT109), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(KEYINPUT109), .B2(new_n968), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT110), .ZN(new_n973));
  INV_X1    g548(.A(G1996), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n966), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n975), .B(KEYINPUT111), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n976), .A2(new_n775), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n719), .B(G2067), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n775), .A2(G1996), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n967), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n817), .B(new_n819), .Z(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n967), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n973), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n883), .A2(new_n965), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT45), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n964), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(G164), .A2(new_n987), .A3(G1384), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G2078), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n988), .A2(new_n990), .A3(KEYINPUT53), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n883), .A2(KEYINPUT45), .A3(new_n965), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n468), .A2(G40), .A3(new_n476), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n993), .A2(new_n994), .A3(new_n991), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT50), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n883), .A2(new_n1000), .A3(new_n965), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n999), .A2(new_n1001), .A3(new_n995), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n766), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n992), .A2(new_n998), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  XNOR2_X1  g580(.A(KEYINPUT114), .B(G8), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G286), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n883), .B2(new_n965), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1008), .A2(new_n989), .A3(new_n964), .ZN(new_n1009));
  OAI221_X1 g584(.A(new_n1007), .B1(G2084), .B2(new_n1002), .C1(new_n1009), .C2(G1966), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n988), .A2(new_n990), .ZN(new_n1011));
  INV_X1    g586(.A(G1966), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n999), .A2(new_n1001), .A3(new_n995), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1011), .A2(new_n1012), .B1(new_n1013), .B2(new_n751), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(G286), .B2(KEYINPUT114), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1010), .B(KEYINPUT51), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1006), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1018), .B(new_n1007), .C1(new_n1014), .C2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT62), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1005), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n1024));
  NAND3_X1  g599(.A1(G303), .A2(new_n1024), .A3(G8), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT55), .B1(G166), .B2(new_n1015), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n882), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n498), .A2(KEYINPUT103), .A3(new_n501), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n496), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(new_n1031), .B2(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(new_n502), .ZN(new_n1033));
  AOI21_X1  g608(.A(G1384), .B1(new_n880), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n964), .B1(new_n1034), .B2(new_n1000), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT117), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1000), .B1(new_n883), .B2(new_n965), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1000), .B(new_n965), .C1(new_n496), .C2(new_n502), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n995), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G2090), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n796), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1028), .B1(new_n1046), .B2(new_n1006), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1017), .A2(KEYINPUT62), .A3(new_n1020), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n1050));
  INV_X1    g625(.A(G1981), .ZN(new_n1051));
  AND3_X1   g626(.A1(new_n608), .A2(new_n1051), .A3(new_n613), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(new_n608), .B2(new_n609), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT49), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n995), .A2(new_n883), .A3(new_n965), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1056), .A2(new_n1006), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT49), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1050), .B(new_n1058), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(G1976), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1056), .B(new_n1006), .C1(new_n1061), .C2(G288), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT52), .ZN(new_n1063));
  INV_X1    g638(.A(G288), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1061), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1057), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1060), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  AOI22_X1  g643(.A1(new_n1013), .A2(new_n1042), .B1(new_n1044), .B2(new_n796), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(new_n1015), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1027), .A2(KEYINPUT113), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1025), .A2(new_n1072), .A3(new_n1026), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1071), .A2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1068), .B1(new_n1070), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1023), .A2(new_n1048), .A3(new_n1049), .A4(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1060), .A2(new_n1061), .A3(new_n1064), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1052), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1077), .A2(KEYINPUT116), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT116), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1014), .A2(G286), .A3(new_n1019), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1060), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1027), .B1(new_n1069), .B2(new_n1015), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1081), .A2(new_n1057), .B1(KEYINPUT63), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1045), .B1(G2090), .B2(new_n1002), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1074), .A2(new_n1087), .A3(G8), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1009), .A2(G1966), .B1(G2084), .B2(new_n1002), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT63), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(new_n1090), .A3(G168), .A4(new_n1006), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1088), .B1(new_n1047), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1083), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT118), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1085), .A2(KEYINPUT63), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1080), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1077), .A2(KEYINPUT116), .A3(new_n1078), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1096), .A2(new_n1057), .A3(new_n1097), .ZN(new_n1098));
  AND4_X1   g673(.A1(KEYINPUT118), .A2(new_n1093), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1076), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n988), .A2(KEYINPUT53), .A3(new_n991), .A4(new_n994), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1102), .A2(new_n998), .A3(new_n1003), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G171), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n996), .A2(new_n997), .B1(new_n1002), .B2(new_n766), .ZN(new_n1105));
  AOI21_X1  g680(.A(G301), .B1(new_n1105), .B2(new_n992), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1101), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1107), .A2(new_n1048), .A3(new_n1075), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(G171), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1105), .A2(G301), .A3(new_n992), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(KEYINPUT54), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1112));
  OAI21_X1  g687(.A(KEYINPUT125), .B1(new_n1108), .B2(new_n1112), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1111), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1019), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1088), .B(new_n1083), .C1(new_n1028), .C2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1105), .A2(G301), .A3(new_n1102), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT54), .B1(new_n1005), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1114), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n584), .B2(new_n564), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n559), .A2(new_n561), .ZN(new_n1125));
  AND4_X1   g700(.A1(new_n1123), .A2(new_n578), .A3(new_n572), .A4(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n579), .A2(KEYINPUT57), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n584), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n761), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT56), .B(G2072), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n1133), .ZN(new_n1134));
  AND4_X1   g709(.A1(new_n1127), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1056), .ZN(new_n1136));
  INV_X1    g711(.A(G2067), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1002), .A2(new_n833), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NOR3_X1   g713(.A1(new_n1138), .A2(KEYINPUT120), .A3(new_n923), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1127), .A2(new_n1131), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT120), .B1(new_n1138), .B2(new_n923), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1135), .B2(new_n1140), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1127), .A2(new_n1131), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT61), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1056), .A2(G2067), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1152), .B(new_n1153), .C1(new_n833), .C2(new_n1002), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT124), .B1(new_n1154), .B2(new_n923), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1154), .A2(new_n1156), .A3(new_n923), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1138), .A2(KEYINPUT60), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n1158), .B2(new_n629), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1158), .A2(new_n1160), .A3(new_n629), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1155), .A2(new_n1157), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1138), .A2(KEYINPUT60), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1151), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1044), .A2(KEYINPUT121), .A3(G1996), .ZN(new_n1165));
  XOR2_X1   g740(.A(KEYINPUT58), .B(G1341), .Z(new_n1166));
  NAND2_X1  g741(.A1(new_n1056), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT121), .B1(new_n1044), .B2(G1996), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(new_n549), .A3(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1170), .A2(KEYINPUT59), .ZN(new_n1173));
  XNOR2_X1  g748(.A(new_n1172), .B(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1143), .B1(new_n1164), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1122), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n985), .B1(new_n1100), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n817), .A2(new_n819), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n982), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n719), .A2(G2067), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1178), .B(new_n966), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n982), .B2(new_n1179), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT126), .B1(new_n1183), .B2(new_n967), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n967), .B1(new_n979), .B2(new_n885), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(KEYINPUT127), .B2(KEYINPUT46), .ZN(new_n1187));
  NOR2_X1   g762(.A1(KEYINPUT127), .A2(KEYINPUT46), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n976), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n976), .A2(new_n1188), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(new_n1191), .B(KEYINPUT47), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n970), .B(KEYINPUT48), .Z(new_n1193));
  OR2_X1    g768(.A1(new_n984), .A2(new_n1193), .ZN(new_n1194));
  AND3_X1   g769(.A1(new_n1185), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1177), .A2(new_n1195), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g771(.A(G319), .ZN(new_n1198));
  NOR2_X1   g772(.A1(G229), .A2(new_n1198), .ZN(new_n1199));
  AND2_X1   g773(.A1(new_n909), .A2(new_n1199), .ZN(new_n1200));
  NOR2_X1   g774(.A1(G401), .A2(G227), .ZN(new_n1201));
  AND4_X1   g775(.A1(new_n960), .A2(new_n1200), .A3(new_n958), .A4(new_n1201), .ZN(G308));
  NAND4_X1  g776(.A1(new_n1200), .A2(new_n958), .A3(new_n960), .A4(new_n1201), .ZN(G225));
endmodule


