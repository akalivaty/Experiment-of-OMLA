//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND4_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT84), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n187), .A2(new_n188), .A3(G214), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT82), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n187), .A2(new_n188), .A3(KEYINPUT82), .A4(G214), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT83), .ZN(new_n198));
  AOI21_X1  g012(.A(G143), .B1(new_n192), .B2(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n200), .A3(new_n196), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n191), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT18), .A2(G131), .ZN(new_n203));
  XNOR2_X1  g017(.A(G125), .B(G140), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(new_n204), .A2(new_n205), .ZN(new_n207));
  AOI22_X1  g021(.A1(new_n202), .A2(new_n203), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n189), .B(KEYINPUT84), .ZN(new_n209));
  AND4_X1   g023(.A1(new_n200), .A2(new_n194), .A3(new_n195), .A4(new_n196), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n200), .B1(new_n199), .B2(new_n196), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(KEYINPUT18), .A3(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g028(.A(G113), .B(G122), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT85), .B(G104), .ZN(new_n216));
  XOR2_X1   g030(.A(new_n215), .B(new_n216), .Z(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(G131), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n221), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n224));
  INV_X1    g038(.A(G125), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n225), .A2(G140), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n224), .B1(KEYINPUT16), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n205), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n224), .B(G146), .C1(KEYINPUT16), .C2(new_n226), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n231), .B1(new_n219), .B2(new_n220), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n214), .B(new_n218), .C1(new_n223), .C2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT87), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n219), .A2(new_n220), .A3(new_n222), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n202), .A2(new_n221), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT17), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n237), .A3(new_n231), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n238), .A2(new_n239), .A3(new_n214), .A4(new_n218), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n234), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n222), .ZN(new_n242));
  XOR2_X1   g056(.A(new_n204), .B(KEYINPUT19), .Z(new_n243));
  OAI21_X1  g057(.A(new_n229), .B1(new_n243), .B2(G146), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n242), .A2(new_n245), .B1(new_n208), .B2(new_n213), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT86), .B1(new_n246), .B2(new_n218), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT86), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n208), .A2(new_n213), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n219), .B2(new_n222), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n248), .B(new_n217), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n241), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT88), .ZN(new_n254));
  NOR2_X1   g068(.A1(G475), .A2(G902), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n254), .A3(KEYINPUT20), .A4(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT88), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(KEYINPUT88), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n234), .A2(new_n240), .B1(new_n247), .B2(new_n251), .ZN(new_n261));
  INV_X1    g075(.A(new_n255), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n258), .B(new_n260), .C1(new_n261), .C2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n218), .B1(new_n238), .B2(new_n214), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n264), .B1(new_n234), .B2(new_n240), .ZN(new_n265));
  OAI21_X1  g079(.A(G475), .B1(new_n265), .B2(G902), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n256), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT90), .B1(new_n195), .B2(G128), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT90), .ZN(new_n270));
  INV_X1    g084(.A(G128), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(G143), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n269), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n271), .B2(G143), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n195), .A2(KEYINPUT13), .A3(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G134), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n269), .A2(new_n272), .ZN(new_n279));
  INV_X1    g093(.A(G134), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n195), .A2(G128), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT92), .ZN(new_n283));
  AOI22_X1  g097(.A1(KEYINPUT91), .A2(new_n278), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n269), .A2(new_n272), .B1(G128), .B2(new_n195), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n285), .B2(new_n280), .ZN(new_n286));
  AND2_X1   g100(.A1(KEYINPUT89), .A2(G122), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT89), .A2(G122), .ZN(new_n288));
  OAI21_X1  g102(.A(G116), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G116), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G122), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n289), .A2(G107), .A3(new_n291), .ZN(new_n292));
  AOI21_X1  g106(.A(G107), .B1(new_n289), .B2(new_n291), .ZN(new_n293));
  NOR3_X1   g107(.A1(new_n286), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n278), .A2(KEYINPUT91), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT9), .B(G234), .ZN(new_n297));
  INV_X1    g111(.A(G217), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(G953), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT93), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n285), .A2(new_n280), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n301), .B2(new_n282), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n279), .A2(new_n281), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G134), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n285), .A2(new_n280), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(KEYINPUT93), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G107), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n289), .B2(KEYINPUT14), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n289), .A2(new_n291), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n302), .A2(new_n306), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n296), .A2(new_n299), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n299), .B1(new_n296), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n268), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT94), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G478), .ZN(new_n318));
  NOR2_X1   g132(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(KEYINPUT95), .A2(KEYINPUT15), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI211_X1 g136(.A(KEYINPUT94), .B(new_n268), .C1(new_n313), .C2(new_n314), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT96), .ZN(new_n325));
  INV_X1    g139(.A(new_n314), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n296), .A2(new_n312), .A3(new_n299), .ZN(new_n327));
  AOI21_X1  g141(.A(G902), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n322), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n317), .A2(new_n325), .A3(new_n322), .A4(new_n323), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT97), .A2(G952), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT97), .A2(G952), .ZN(new_n337));
  AOI21_X1  g151(.A(G953), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G234), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n339), .B2(new_n187), .ZN(new_n340));
  AOI211_X1 g154(.A(new_n268), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT21), .B(G898), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n267), .A2(new_n334), .A3(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(G214), .B1(G237), .B2(G902), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT64), .B1(new_n195), .B2(G146), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT64), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n205), .A3(G143), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n195), .A2(G146), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(KEYINPUT0), .A2(G128), .ZN(new_n354));
  NOR2_X1   g168(.A1(KEYINPUT0), .A2(G128), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G143), .B(G146), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n353), .A2(new_n356), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(new_n225), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n271), .A2(KEYINPUT1), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n205), .A2(G143), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n352), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(KEYINPUT65), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT65), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n365), .A3(new_n361), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n195), .A2(G146), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT1), .ZN(new_n368));
  OAI21_X1  g182(.A(G128), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n364), .A2(new_n366), .B1(new_n353), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n225), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n348), .B1(new_n360), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G224), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G953), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n359), .A2(KEYINPUT79), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n374), .B1(new_n372), .B2(new_n375), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G116), .ZN(new_n380));
  OAI21_X1  g194(.A(G113), .B1(new_n380), .B2(KEYINPUT5), .ZN(new_n381));
  XNOR2_X1  g195(.A(G116), .B(G119), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n381), .B1(KEYINPUT5), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(KEYINPUT2), .A2(G113), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT66), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT66), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT2), .A3(G113), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  OR2_X1    g202(.A1(KEYINPUT2), .A2(G113), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(new_n382), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  AOI21_X1  g207(.A(G101), .B1(new_n392), .B2(G107), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n395), .A2(new_n307), .A3(G104), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT74), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n393), .A2(new_n394), .A3(new_n396), .A4(KEYINPUT74), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(G107), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n307), .A2(G104), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(KEYINPUT76), .B1(new_n401), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n408));
  AOI211_X1 g222(.A(new_n408), .B(new_n405), .C1(new_n399), .C2(new_n400), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n391), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n393), .A2(new_n396), .A3(new_n403), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(G101), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT75), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT75), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n411), .A2(new_n415), .A3(new_n412), .A4(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n412), .B1(new_n411), .B2(G101), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n386), .B1(KEYINPUT2), .B2(G113), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n384), .A2(KEYINPUT66), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n389), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n382), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n388), .A2(new_n389), .A3(new_n382), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(KEYINPUT67), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT67), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n427), .B1(new_n390), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n417), .A2(new_n419), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n410), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT78), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n410), .A2(KEYINPUT78), .A3(new_n430), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G122), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n433), .A2(new_n434), .A3(new_n435), .A4(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n410), .A2(KEYINPUT78), .A3(new_n430), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT78), .B1(new_n410), .B2(new_n430), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(new_n436), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n410), .A2(new_n430), .A3(new_n436), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT6), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n378), .B(new_n438), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n436), .B(KEYINPUT8), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n401), .A2(new_n406), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n390), .B2(new_n383), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n445), .B1(new_n410), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n449), .B2(KEYINPUT7), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT7), .ZN(new_n451));
  OAI22_X1  g265(.A1(new_n372), .A2(new_n375), .B1(new_n451), .B2(new_n374), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(new_n442), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n444), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT81), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n444), .A2(new_n457), .A3(new_n454), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n455), .A2(KEYINPUT80), .ZN(new_n459));
  AOI22_X1  g273(.A1(KEYINPUT81), .A2(new_n456), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n459), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n444), .A2(new_n457), .A3(new_n454), .A4(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n347), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n379), .A2(G128), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n271), .A2(G119), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT71), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT24), .B(G110), .Z(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n271), .A2(KEYINPUT23), .A3(G119), .ZN(new_n470));
  INV_X1    g284(.A(new_n465), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n464), .B(new_n470), .C1(new_n471), .C2(KEYINPUT23), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(G110), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n229), .B(new_n206), .C1(new_n469), .C2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n467), .A2(new_n468), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(G110), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n230), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT22), .B(G137), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n479), .B(new_n480), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n474), .A2(new_n477), .A3(new_n481), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT25), .ZN(new_n485));
  AOI21_X1  g299(.A(G902), .B1(new_n485), .B2(KEYINPUT72), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n485), .A2(KEYINPUT72), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G217), .B1(new_n339), .B2(G902), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n487), .B2(new_n488), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n483), .A2(new_n484), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n339), .B2(G217), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n429), .A2(new_n426), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n353), .A2(new_n369), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n365), .B1(new_n357), .B2(new_n361), .ZN(new_n499));
  AND4_X1   g313(.A1(new_n365), .A2(new_n361), .A3(new_n362), .A4(new_n352), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT11), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n280), .B2(G137), .ZN(new_n503));
  INV_X1    g317(.A(G137), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(KEYINPUT11), .A3(G134), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n280), .A2(G137), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n503), .A2(new_n505), .A3(new_n221), .A4(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n280), .A2(G137), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n504), .A2(G134), .ZN(new_n509));
  OAI21_X1  g323(.A(G131), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n501), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n503), .A2(new_n505), .A3(new_n506), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G131), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n507), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n358), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n513), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n514), .B1(new_n513), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n497), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT68), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n518), .B1(new_n370), .B2(new_n511), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n522), .B1(new_n497), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n501), .A2(new_n512), .B1(new_n517), .B2(new_n358), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n429), .A2(new_n426), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT68), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n187), .A2(new_n188), .A3(G210), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT27), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT26), .B(G101), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n521), .A2(new_n524), .A3(new_n527), .A4(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT31), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT68), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT68), .B1(new_n525), .B2(new_n526), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(KEYINPUT31), .A3(new_n531), .A4(new_n521), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT28), .B1(new_n525), .B2(new_n526), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n525), .A2(new_n526), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n535), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT28), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n531), .B(KEYINPUT69), .Z(new_n545));
  AOI22_X1  g359(.A1(new_n534), .A2(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT32), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n534), .A2(new_n538), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n497), .A2(new_n523), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n543), .B1(new_n537), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n545), .B1(new_n552), .B2(new_n539), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n547), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n531), .A2(KEYINPUT29), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n524), .A2(new_n551), .A3(new_n527), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n539), .B(new_n558), .C1(new_n559), .C2(KEYINPUT28), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT70), .B1(new_n560), .B2(G902), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n562), .B(new_n268), .C1(new_n544), .C2(new_n558), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n537), .A2(new_n521), .ZN(new_n564));
  INV_X1    g378(.A(new_n531), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT29), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(new_n544), .B2(new_n545), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n561), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G472), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n496), .B1(new_n557), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  OR2_X1    g385(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(KEYINPUT77), .ZN(new_n573));
  INV_X1    g387(.A(new_n369), .ZN(new_n574));
  OAI22_X1  g388(.A1(new_n500), .A2(new_n499), .B1(new_n574), .B2(new_n357), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n405), .B1(new_n399), .B2(new_n400), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n407), .A2(new_n409), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n370), .ZN(new_n580));
  INV_X1    g394(.A(new_n517), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n572), .B(new_n573), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n446), .A2(new_n408), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n576), .A2(KEYINPUT76), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n370), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n577), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n586), .A2(KEYINPUT77), .A3(new_n571), .A4(new_n517), .ZN(new_n587));
  OAI211_X1 g401(.A(KEYINPUT10), .B(new_n501), .C1(new_n407), .C2(new_n409), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n577), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n417), .A2(new_n419), .A3(new_n358), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n581), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n582), .A2(new_n587), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(G110), .B(G140), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n188), .A2(G227), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(G469), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n517), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n596), .A3(new_n592), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n598), .A2(new_n599), .A3(new_n268), .A4(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n599), .A2(new_n268), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(new_n596), .B(KEYINPUT73), .Z(new_n606));
  NAND2_X1  g420(.A1(new_n593), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n601), .A2(new_n597), .A3(new_n592), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(G469), .A3(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(G221), .B1(new_n297), .B2(G902), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n345), .A2(new_n463), .A3(new_n570), .A4(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  INV_X1    g429(.A(new_n496), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n548), .B1(new_n550), .B2(new_n553), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n554), .A2(new_n268), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(G472), .ZN(new_n619));
  AND4_X1   g433(.A1(new_n616), .A2(new_n619), .A3(new_n611), .A4(new_n610), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n318), .A2(G902), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT33), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n326), .B2(new_n327), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT33), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n621), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n628));
  OAI211_X1 g442(.A(KEYINPUT98), .B(new_n621), .C1(new_n623), .C2(new_n624), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n267), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n344), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n444), .A2(new_n454), .A3(new_n455), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n455), .B1(new_n444), .B2(new_n454), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n633), .B(new_n346), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n620), .A2(new_n632), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND4_X1  g454(.A1(new_n256), .A2(new_n263), .A3(new_n331), .A4(new_n332), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n266), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(KEYINPUT99), .B(G475), .C1(new_n265), .C2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n620), .A2(new_n637), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NOR2_X1   g463(.A1(new_n482), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n478), .B(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n489), .A2(new_n491), .B1(new_n494), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT100), .B1(new_n619), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(G472), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n554), .B2(new_n268), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n656), .A2(new_n652), .A3(new_n617), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n458), .A2(new_n459), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n661), .A3(new_n462), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n346), .A2(new_n662), .A3(new_n611), .A4(new_n610), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n659), .A2(new_n663), .A3(new_n345), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  AOI22_X1  g480(.A1(new_n549), .A2(new_n556), .B1(new_n568), .B2(G472), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n346), .B1(new_n634), .B2(new_n635), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n667), .A2(new_n668), .A3(new_n652), .ZN(new_n669));
  INV_X1    g483(.A(new_n340), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n670), .B1(new_n671), .B2(new_n341), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n641), .A2(new_n645), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n673), .A3(new_n613), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XOR2_X1   g489(.A(new_n672), .B(KEYINPUT39), .Z(new_n676));
  NAND3_X1  g490(.A1(new_n610), .A2(new_n611), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT40), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n267), .A2(new_n334), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n559), .A2(new_n545), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n532), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n655), .B1(new_n682), .B2(new_n268), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n549), .B2(new_n556), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n680), .A2(new_n684), .A3(new_n347), .A4(new_n653), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n662), .B(KEYINPUT38), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G143), .ZN(G45));
  INV_X1    g502(.A(new_n672), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n267), .A2(new_n630), .A3(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n652), .B1(new_n557), .B2(new_n569), .ZN(new_n692));
  INV_X1    g506(.A(new_n668), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n691), .A2(new_n692), .A3(new_n693), .A4(new_n613), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND3_X1  g509(.A1(new_n598), .A2(new_n268), .A3(new_n602), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n697), .A3(G469), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(G469), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n598), .A2(new_n268), .A3(new_n602), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n611), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n632), .A2(new_n702), .A3(new_n570), .A4(new_n637), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT41), .B(G113), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NAND4_X1  g519(.A1(new_n646), .A2(new_n570), .A3(new_n637), .A4(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G116), .ZN(G18));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n668), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n345), .A2(new_n708), .A3(new_n692), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  INV_X1    g524(.A(new_n656), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n539), .B1(new_n559), .B2(KEYINPUT28), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(KEYINPUT102), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n545), .B1(new_n712), .B2(KEYINPUT102), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n550), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n547), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n711), .A2(new_n716), .A3(new_n616), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n701), .A3(new_n344), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n668), .B1(new_n680), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n267), .A2(KEYINPUT103), .A3(new_n334), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n718), .A2(new_n720), .A3(new_n724), .A4(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND3_X1  g541(.A1(new_n711), .A2(new_n716), .A3(new_n653), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n690), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n708), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT105), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n608), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n601), .A2(KEYINPUT105), .A3(new_n597), .A4(new_n592), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n607), .A2(G469), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n603), .A2(new_n737), .A3(new_n605), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(KEYINPUT106), .A3(new_n611), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT106), .B1(new_n738), .B2(new_n611), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n662), .B2(new_n347), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n460), .A2(KEYINPUT107), .A3(new_n346), .A4(new_n462), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n741), .A2(new_n570), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n733), .B1(new_n745), .B2(new_n690), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n738), .A2(new_n611), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT106), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n738), .A2(KEYINPUT106), .A3(new_n611), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n743), .A2(new_n744), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT108), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(KEYINPUT42), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n751), .A2(new_n570), .A3(new_n691), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n746), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  INV_X1    g571(.A(new_n673), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n745), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n280), .ZN(G36));
  INV_X1    g574(.A(new_n611), .ZN(new_n761));
  INV_X1    g575(.A(new_n603), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n607), .A2(new_n608), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n607), .A2(KEYINPUT45), .A3(new_n735), .A4(new_n736), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(G469), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT109), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT109), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n769), .A3(G469), .A4(new_n766), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n605), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n762), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n773), .B(new_n604), .C1(new_n768), .C2(new_n770), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n761), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n256), .A2(new_n263), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT43), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n266), .A4(new_n630), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n630), .A2(new_n256), .A3(new_n263), .A4(new_n266), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT43), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n619), .A2(new_n652), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n780), .A2(new_n782), .A3(KEYINPUT44), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT110), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n743), .A2(new_n744), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n780), .A2(new_n782), .A3(new_n783), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT44), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n777), .A2(new_n785), .A3(new_n676), .A4(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  AOI21_X1  g605(.A(new_n604), .B1(new_n768), .B2(new_n770), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n603), .B1(new_n792), .B2(KEYINPUT46), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n611), .B1(new_n793), .B2(new_n775), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g610(.A(KEYINPUT47), .B(new_n611), .C1(new_n793), .C2(new_n775), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n743), .A2(new_n744), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(new_n667), .A3(new_n496), .A4(new_n691), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT111), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n798), .A2(KEYINPUT111), .A3(new_n801), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n652), .A2(new_n689), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n747), .A2(new_n684), .A3(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n720), .A2(new_n811), .A3(new_n721), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n674), .A3(new_n694), .A4(new_n730), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n667), .A2(new_n612), .A3(new_n668), .A4(new_n652), .ZN(new_n816));
  AOI22_X1  g630(.A1(new_n816), .A2(new_n673), .B1(new_n729), .B2(new_n708), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n817), .A2(KEYINPUT52), .A3(new_n694), .A4(new_n812), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n749), .A2(new_n750), .ZN(new_n820));
  INV_X1    g634(.A(new_n570), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n786), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n822), .A2(new_n673), .B1(new_n729), .B2(new_n751), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n333), .A2(KEYINPUT112), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n331), .A2(new_n825), .A3(new_n332), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n631), .B1(new_n827), .B2(new_n267), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n620), .A3(new_n633), .A4(new_n463), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n664), .A2(new_n829), .A3(new_n614), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n331), .A2(new_n825), .A3(new_n332), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n331), .B2(new_n332), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n689), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n778), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n645), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n613), .A3(new_n836), .A4(new_n692), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT113), .B1(new_n837), .B2(new_n786), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n672), .B1(new_n824), .B2(new_n826), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n778), .A2(new_n692), .A3(new_n839), .A4(new_n836), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n799), .A3(new_n841), .A4(new_n613), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n830), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n819), .A2(new_n823), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n703), .A2(new_n709), .A3(new_n706), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n845), .B1(new_n723), .B2(new_n725), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n756), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n809), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n838), .A2(new_n842), .ZN(new_n849));
  INV_X1    g663(.A(new_n830), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n849), .A2(new_n823), .A3(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n756), .A2(new_n846), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n809), .B1(new_n817), .B2(new_n814), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n819), .A4(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n808), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n817), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n809), .B1(new_n856), .B2(KEYINPUT52), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n819), .A2(new_n843), .A3(new_n823), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n756), .A2(new_n846), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n860), .B1(new_n756), .B2(new_n846), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n851), .A2(new_n852), .A3(new_n819), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n859), .A2(new_n863), .B1(new_n864), .B2(new_n809), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n855), .B1(new_n808), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n780), .A2(new_n782), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n670), .A2(new_n799), .A3(new_n702), .A4(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n570), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n869), .A2(new_n870), .A3(KEYINPUT48), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n867), .A2(new_n670), .ZN(new_n872));
  INV_X1    g686(.A(new_n717), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n708), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT116), .ZN(new_n875));
  XNOR2_X1  g689(.A(KEYINPUT117), .B(KEYINPUT48), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n338), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n684), .A2(new_n616), .A3(new_n670), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n786), .A2(new_n701), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n878), .B1(new_n880), .B2(new_n632), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n871), .A2(new_n875), .A3(new_n877), .A4(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n686), .A2(new_n346), .A3(new_n701), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n872), .A2(new_n883), .A3(KEYINPUT50), .A4(new_n873), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n662), .B(KEYINPUT38), .Z(new_n886));
  NAND3_X1  g700(.A1(new_n886), .A2(new_n347), .A3(new_n702), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n867), .A2(new_n670), .A3(new_n873), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(new_n728), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n267), .A2(new_n630), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n868), .A2(new_n891), .B1(new_n880), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n698), .A2(new_n700), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n796), .B(new_n797), .C1(new_n611), .C2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n888), .A2(new_n786), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n882), .B1(KEYINPUT51), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(KEYINPUT51), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(KEYINPUT115), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n866), .B(new_n899), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(G952), .A2(G953), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n895), .A2(KEYINPUT49), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n496), .A2(new_n347), .A3(new_n761), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n684), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n895), .A2(KEYINPUT49), .ZN(new_n909));
  OR4_X1    g723(.A1(new_n686), .A2(new_n908), .A3(new_n781), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n910), .ZN(G75));
  NAND2_X1  g725(.A1(new_n863), .A2(new_n859), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n848), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n913), .A2(G210), .A3(G902), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n441), .A2(new_n443), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n434), .B2(new_n441), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n378), .ZN(new_n918));
  XOR2_X1   g732(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n914), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n920), .B1(new_n914), .B2(new_n915), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n188), .A2(G952), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G51));
  AND3_X1   g738(.A1(new_n819), .A2(new_n823), .A3(new_n843), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n925), .B2(new_n852), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT54), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n862), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n756), .A2(new_n846), .A3(new_n860), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n848), .B(new_n808), .C1(new_n931), .C2(new_n858), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n604), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n598), .A3(new_n602), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n913), .A2(G902), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(new_n771), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n923), .B1(new_n937), .B2(new_n939), .ZN(G54));
  NAND2_X1  g754(.A1(KEYINPUT58), .A2(G475), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n261), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n923), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n938), .A2(new_n261), .A3(new_n941), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n944), .A2(new_n945), .ZN(G60));
  INV_X1    g760(.A(KEYINPUT120), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n623), .A2(new_n624), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(G478), .A2(G902), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT59), .Z(new_n951));
  OAI211_X1 g765(.A(new_n947), .B(new_n949), .C1(new_n866), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n848), .A2(new_n854), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(new_n932), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT120), .B1(new_n955), .B2(new_n948), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n949), .A2(new_n951), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n923), .B1(new_n933), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n952), .A2(new_n956), .A3(new_n958), .ZN(G63));
  XNOR2_X1  g773(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n298), .A2(new_n268), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n926), .B2(new_n927), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n493), .B(KEYINPUT123), .Z(new_n964));
  AOI21_X1  g778(.A(new_n923), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n913), .A2(new_n651), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n963), .A2(new_n964), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT122), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n969), .A3(new_n943), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n967), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n965), .B(new_n966), .C1(new_n969), .C2(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(G66));
  NAND2_X1  g788(.A1(new_n846), .A2(new_n850), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n188), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n342), .B2(new_n373), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(KEYINPUT124), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(KEYINPUT124), .B2(new_n976), .ZN(new_n979));
  INV_X1    g793(.A(G898), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n917), .B1(new_n980), .B2(G953), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n979), .B(new_n981), .ZN(G69));
  NAND3_X1  g796(.A1(new_n720), .A2(new_n570), .A3(new_n721), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n777), .A2(new_n676), .A3(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n674), .A2(new_n694), .A3(new_n730), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n759), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n790), .A2(new_n756), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n988), .B1(new_n804), .B2(new_n805), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n188), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n519), .A2(new_n520), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(new_n243), .Z(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n990), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n817), .A2(new_n687), .A3(new_n694), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(KEYINPUT62), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n995), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n784), .A2(KEYINPUT110), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n784), .A2(KEYINPUT110), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n789), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n611), .B(new_n676), .C1(new_n793), .C2(new_n775), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n817), .A2(new_n687), .A3(new_n1006), .A4(new_n694), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n821), .A2(new_n677), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n799), .A2(new_n1008), .A3(new_n828), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1005), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(KEYINPUT111), .B1(new_n798), .B2(new_n801), .ZN(new_n1012));
  AOI211_X1 g826(.A(new_n803), .B(new_n800), .C1(new_n796), .C2(new_n797), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1000), .B(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1014));
  AND2_X1   g828(.A1(new_n1014), .A2(new_n188), .ZN(new_n1015));
  INV_X1    g829(.A(new_n992), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n994), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n1017), .B(new_n1018), .ZN(G72));
  INV_X1    g833(.A(new_n564), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n565), .ZN(new_n1021));
  OAI211_X1 g835(.A(new_n756), .B(new_n987), .C1(new_n1004), .C2(new_n983), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(new_n1005), .ZN(new_n1023));
  INV_X1    g837(.A(new_n975), .ZN(new_n1024));
  OAI211_X1 g838(.A(new_n1023), .B(new_n1024), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  AOI21_X1  g841(.A(new_n1021), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(KEYINPUT127), .B1(new_n1028), .B2(new_n923), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT127), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1027), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1031), .B1(new_n989), .B2(new_n1024), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1030), .B(new_n943), .C1(new_n1032), .C2(new_n1021), .ZN(new_n1033));
  AND2_X1   g847(.A1(new_n1029), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1020), .A2(new_n565), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1035), .A2(new_n1031), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n953), .A2(new_n1021), .A3(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1027), .B1(new_n1014), .B2(new_n975), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT126), .ZN(new_n1039));
  AND3_X1   g853(.A1(new_n1038), .A2(new_n1039), .A3(new_n1035), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1039), .B1(new_n1038), .B2(new_n1035), .ZN(new_n1041));
  OAI21_X1  g855(.A(new_n1037), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1034), .A2(new_n1042), .ZN(G57));
endmodule


