//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n558, new_n559, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n455));
  XOR2_X1   g030(.A(KEYINPUT69), .B(KEYINPUT2), .Z(new_n456));
  XNOR2_X1  g031(.A(new_n455), .B(new_n456), .ZN(new_n457));
  NOR4_X1   g032(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n457), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n457), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT70), .B(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n465), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(G137), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n466), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n469), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2104), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT3), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n464), .ZN(new_n485));
  OR3_X1    g060(.A1(new_n485), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT71), .B1(new_n485), .B2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G136), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n485), .A2(new_n468), .ZN(new_n491));
  OR2_X1    g066(.A1(new_n468), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n491), .A2(G124), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G162));
  NAND4_X1  g072(.A1(new_n484), .A2(G126), .A3(G2105), .A4(new_n464), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n484), .A2(new_n464), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT72), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n484), .A2(new_n506), .A3(new_n464), .A4(new_n503), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n505), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n508));
  NOR4_X1   g083(.A1(new_n473), .A2(KEYINPUT4), .A3(new_n502), .A4(G2105), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n501), .B1(new_n508), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n512), .B2(G651), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n512), .A2(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n517), .A2(new_n518), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G88), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n524), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(new_n515), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n526), .A2(G89), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n520), .A2(G51), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AND2_X1   g111(.A1(G63), .A2(G651), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n535), .A2(new_n536), .B1(new_n524), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n532), .A2(new_n533), .A3(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n526), .A2(G90), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n520), .A2(G52), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n524), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n515), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(G301));
  INV_X1    g120(.A(G301), .ZN(G171));
  AOI22_X1  g121(.A1(new_n524), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n515), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n549), .A2(new_n519), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  AND2_X1   g126(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(KEYINPUT74), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n548), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n520), .A2(G53), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n561), .A2(KEYINPUT75), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n524), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n526), .A2(G91), .B1(new_n567), .B2(G651), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n561), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n520), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(KEYINPUT9), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n569), .A2(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n520), .A2(G49), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n526), .A2(G87), .ZN(new_n576));
  OAI21_X1  g151(.A(G651), .B1(new_n524), .B2(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  NAND2_X1  g153(.A1(new_n526), .A2(G86), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n520), .A2(G48), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n565), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G651), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n526), .A2(G85), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n520), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n586), .B(new_n587), .C1(new_n515), .C2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G54), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n519), .B1(new_n592), .B2(new_n515), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n517), .A2(G92), .A3(new_n518), .A4(new_n524), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(KEYINPUT76), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n596), .ZN(new_n600));
  AND2_X1   g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n590), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  AND2_X1   g179(.A1(new_n569), .A2(new_n573), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G297));
  OAI21_X1  g181(.A(new_n604), .B1(new_n605), .B2(G868), .ZN(G280));
  XNOR2_X1  g182(.A(KEYINPUT77), .B(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n601), .B1(G860), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT78), .ZN(G148));
  NOR2_X1   g185(.A1(new_n555), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n601), .A2(new_n608), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(G868), .B2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT79), .Z(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g190(.A(new_n473), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n477), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT12), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n468), .A2(G111), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n621), .A2(KEYINPUT80), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n621), .B2(KEYINPUT80), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n491), .A2(G123), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(G135), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n488), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n620), .A2(new_n628), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n641), .B2(new_n644), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(G401));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT83), .Z(new_n650));
  NOR2_X1   g225(.A1(G2072), .A2(G2078), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n444), .A2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n648), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n652), .B(KEYINPUT17), .Z(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n655), .B2(new_n650), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n652), .A2(new_n649), .A3(new_n648), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n650), .A3(new_n648), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT84), .B(G2096), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n668));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n670), .A2(new_n664), .A3(new_n665), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n664), .B(new_n665), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n673), .B(new_n674), .C1(new_n670), .C2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1991), .B(G1996), .Z(new_n677));
  XOR2_X1   g252(.A(new_n676), .B(new_n677), .Z(new_n678));
  XOR2_X1   g253(.A(G1981), .B(G1986), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT87), .ZN(new_n680));
  XOR2_X1   g255(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n678), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(G229));
  NAND2_X1  g259(.A1(new_n489), .A2(G131), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n491), .A2(G119), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT88), .ZN(new_n687));
  OAI21_X1  g262(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR3_X1   g264(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n690));
  OAI221_X1 g265(.A(G2104), .B1(G107), .B2(new_n468), .C1(new_n689), .C2(new_n690), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n685), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G29), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G25), .B2(G29), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT35), .B(G1991), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  MUX2_X1   g273(.A(G24), .B(G290), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1986), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n697), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT32), .B(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1971), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(G23), .ZN(new_n709));
  INV_X1    g284(.A(G288), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n705), .ZN(new_n711));
  XOR2_X1   g286(.A(KEYINPUT33), .B(G1976), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR3_X1   g288(.A1(new_n704), .A2(new_n708), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT34), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  NAND3_X1  g292(.A1(new_n701), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT36), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n705), .A2(G4), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n601), .B2(new_n705), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1348), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT93), .ZN(new_n724));
  INV_X1    g299(.A(G29), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G26), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n724), .B(new_n726), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n491), .A2(G128), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n468), .A2(G116), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n730));
  INV_X1    g305(.A(G140), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n728), .B1(new_n729), .B2(new_n730), .C1(new_n488), .C2(new_n731), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n732), .A2(KEYINPUT91), .A3(G29), .ZN(new_n733));
  AOI21_X1  g308(.A(KEYINPUT91), .B1(new_n732), .B2(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT94), .B(G2067), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1341), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G19), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(new_n555), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT90), .Z(new_n741));
  AOI211_X1 g316(.A(new_n722), .B(new_n737), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G33), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT95), .Z(new_n744));
  NAND3_X1  g319(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT25), .Z(new_n746));
  AOI22_X1  g321(.A1(new_n616), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n747));
  INV_X1    g322(.A(G139), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n746), .B1(new_n468), .B2(new_n747), .C1(new_n488), .C2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n744), .B1(new_n749), .B2(new_n725), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(new_n442), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT97), .Z(new_n753));
  OR2_X1    g328(.A1(new_n751), .A2(new_n442), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n705), .A2(G20), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT23), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(new_n605), .B2(new_n705), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT100), .B(G1956), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G29), .A2(G35), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(G162), .B2(G29), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT29), .B(G2090), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n725), .A2(G32), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n489), .A2(G141), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n477), .A2(G105), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n767), .B(new_n768), .C1(G129), .C2(new_n491), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(new_n725), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  NAND4_X1  g349(.A1(new_n754), .A2(new_n759), .A3(new_n763), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n627), .A2(new_n725), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(KEYINPUT98), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n705), .A2(G21), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G168), .B2(new_n705), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n777), .B1(G1966), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n705), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n705), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1961), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n779), .A2(G1966), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n776), .B2(KEYINPUT98), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT30), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G28), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n725), .B1(new_n786), .B2(G28), .ZN(new_n788));
  AND2_X1   g363(.A1(KEYINPUT31), .A2(G11), .ZN(new_n789));
  NOR2_X1   g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  OAI22_X1  g365(.A1(new_n787), .A2(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G34), .ZN(new_n792));
  AOI21_X1  g367(.A(G29), .B1(new_n792), .B2(KEYINPUT24), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(KEYINPUT24), .B2(new_n792), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n479), .B2(new_n725), .ZN(new_n795));
  INV_X1    g370(.A(G2084), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n791), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  NOR4_X1   g373(.A1(new_n780), .A2(new_n783), .A3(new_n785), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n725), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n725), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT99), .B(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n803), .C1(new_n741), .C2(new_n738), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n753), .A2(new_n775), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n719), .A2(new_n742), .A3(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n526), .A2(G93), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n520), .A2(G55), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n808), .B(new_n809), .C1(new_n515), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G860), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT37), .Z(new_n813));
  NAND2_X1  g388(.A1(new_n601), .A2(G559), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OR2_X1    g391(.A1(new_n554), .A2(new_n811), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n554), .A2(new_n811), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n816), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT39), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT102), .Z(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n820), .B2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n813), .B1(new_n822), .B2(new_n824), .ZN(G145));
  AOI21_X1  g400(.A(new_n506), .B1(new_n467), .B2(new_n503), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n510), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n501), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n732), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n749), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(new_n771), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n771), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n692), .B(new_n618), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n491), .A2(G130), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n468), .A2(G118), .ZN(new_n839));
  OAI21_X1  g414(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n840));
  INV_X1    g415(.A(G142), .ZN(new_n841));
  OAI221_X1 g416(.A(new_n838), .B1(new_n839), .B2(new_n840), .C1(new_n488), .C2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n837), .B(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n835), .A2(new_n836), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n843), .ZN(new_n845));
  OAI22_X1  g420(.A1(new_n833), .A2(new_n834), .B1(new_n845), .B2(KEYINPUT103), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n627), .B(new_n479), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n496), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n844), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n835), .A2(new_n845), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n843), .B1(new_n833), .B2(new_n834), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n851), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(G37), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g431(.A(new_n819), .B(new_n612), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n599), .A2(new_n600), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n858), .B1(new_n605), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n601), .A2(G299), .A3(KEYINPUT104), .ZN(new_n861));
  AOI22_X1  g436(.A1(new_n860), .A2(new_n861), .B1(new_n605), .B2(new_n859), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n605), .A2(new_n859), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT105), .ZN(new_n867));
  OR3_X1    g442(.A1(new_n601), .A2(G299), .A3(KEYINPUT105), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(new_n860), .B2(new_n861), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n869), .A2(new_n870), .B1(new_n871), .B2(new_n866), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n864), .B1(new_n872), .B2(new_n857), .ZN(new_n873));
  XOR2_X1   g448(.A(G290), .B(G305), .Z(new_n874));
  XOR2_X1   g449(.A(G303), .B(G288), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(KEYINPUT42), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n873), .B(new_n877), .ZN(new_n878));
  MUX2_X1   g453(.A(new_n811), .B(new_n878), .S(G868), .Z(G295));
  MUX2_X1   g454(.A(new_n811), .B(new_n878), .S(G868), .Z(G331));
  XOR2_X1   g455(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n881));
  OR2_X1    g456(.A1(G301), .A2(KEYINPUT107), .ZN(new_n882));
  NAND2_X1  g457(.A1(G301), .A2(KEYINPUT107), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(G168), .ZN(new_n884));
  AOI21_X1  g459(.A(G168), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n819), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n882), .A2(G168), .A3(new_n883), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n818), .B(new_n817), .C1(new_n888), .C2(new_n885), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n887), .A2(KEYINPUT108), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n819), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n886), .A2(new_n884), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n891), .A2(KEYINPUT109), .A3(new_n893), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT109), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n889), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n898), .A3(new_n887), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n872), .A2(new_n895), .B1(new_n899), .B2(new_n862), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n876), .ZN(new_n903));
  OAI221_X1 g478(.A(KEYINPUT110), .B1(new_n899), .B2(new_n862), .C1(new_n872), .C2(new_n895), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n869), .A2(new_n870), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n871), .A2(new_n866), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n890), .A2(new_n894), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n896), .A2(new_n898), .A3(new_n887), .ZN(new_n910));
  AOI22_X1  g485(.A1(new_n908), .A2(new_n909), .B1(new_n910), .B2(new_n863), .ZN(new_n911));
  AOI21_X1  g486(.A(G37), .B1(new_n911), .B2(new_n876), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n881), .B1(new_n905), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n854), .B1(new_n900), .B2(new_n903), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n871), .A2(new_n867), .A3(new_n868), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(KEYINPUT41), .B2(new_n862), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(new_n899), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n895), .A2(new_n863), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n876), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n881), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n913), .A2(KEYINPUT44), .A3(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n905), .A2(new_n912), .A3(new_n881), .ZN(new_n924));
  OAI21_X1  g499(.A(KEYINPUT43), .B1(new_n914), .B2(new_n919), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n922), .A2(new_n926), .ZN(G397));
  INV_X1    g502(.A(G1996), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n770), .B(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G2067), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n732), .B(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g507(.A(new_n692), .B(new_n696), .Z(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(G290), .A2(G1986), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G290), .A2(G1986), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(KEYINPUT111), .B(G1384), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n828), .B2(new_n829), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(KEYINPUT45), .ZN(new_n941));
  INV_X1    g516(.A(G40), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n479), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(G303), .A2(G8), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT55), .ZN(new_n948));
  OR3_X1    g523(.A1(new_n947), .A2(KEYINPUT113), .A3(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT113), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n948), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n939), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n509), .B1(new_n954), .B2(new_n505), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT45), .B(new_n953), .C1(new_n955), .C2(new_n501), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT112), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT112), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n940), .A2(new_n958), .A3(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n943), .ZN(new_n961));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n955), .B2(new_n501), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(G1971), .B1(new_n960), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n968), .B(new_n962), .C1(new_n955), .C2(new_n501), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n967), .A2(new_n969), .A3(new_n943), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n970), .A2(G2090), .ZN(new_n971));
  OAI211_X1 g546(.A(G8), .B(new_n952), .C1(new_n966), .C2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT114), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n961), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n974));
  INV_X1    g549(.A(G2090), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n969), .ZN(new_n976));
  AOI21_X1  g551(.A(G1384), .B1(new_n828), .B2(new_n829), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n943), .B1(new_n977), .B2(KEYINPUT45), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n957), .B2(new_n959), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n976), .B1(new_n979), .B2(G1971), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT114), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n980), .A2(new_n981), .A3(G8), .A4(new_n952), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n973), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n952), .B1(new_n980), .B2(G8), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(KEYINPUT45), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n964), .B1(G164), .B2(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n987), .A3(new_n943), .ZN(new_n988));
  INV_X1    g563(.A(G1966), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n974), .A2(new_n796), .A3(new_n969), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(G8), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n993), .A2(G286), .ZN(new_n994));
  INV_X1    g569(.A(G8), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n977), .B2(new_n943), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n710), .A2(G1976), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G1976), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT52), .B1(G288), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g577(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1981), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1005), .B1(new_n584), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1002), .A2(new_n1007), .A3(new_n1003), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n996), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1001), .B(new_n1011), .C1(new_n1012), .C2(new_n998), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n994), .A2(new_n1014), .A3(KEYINPUT63), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n984), .A2(new_n985), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1013), .B1(new_n985), .B2(KEYINPUT116), .ZN(new_n1017));
  INV_X1    g592(.A(new_n952), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n960), .A2(new_n965), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n971), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1018), .B1(new_n1021), .B2(new_n995), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AND4_X1   g599(.A1(new_n983), .A2(new_n1017), .A3(new_n1024), .A4(new_n994), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT63), .B1(new_n1025), .B2(KEYINPUT117), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT117), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n983), .A2(new_n1017), .A3(new_n1024), .ZN(new_n1028));
  INV_X1    g603(.A(new_n994), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1016), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AND3_X1   g606(.A1(new_n983), .A2(new_n1017), .A3(new_n1024), .ZN(new_n1032));
  INV_X1    g607(.A(new_n970), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1033), .A2(new_n796), .B1(new_n988), .B2(new_n989), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G286), .A2(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n1035), .B2(KEYINPUT123), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1035), .B(new_n1039), .C1(new_n1034), .C2(new_n995), .ZN(new_n1040));
  OAI211_X1 g615(.A(G8), .B(new_n1038), .C1(new_n992), .C2(G286), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT62), .ZN(new_n1043));
  OR2_X1    g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n958), .B1(new_n940), .B2(KEYINPUT45), .ZN(new_n1045));
  NOR4_X1   g620(.A1(G164), .A2(KEYINPUT112), .A3(new_n964), .A4(new_n939), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n965), .B(new_n443), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(G2078), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n965), .A2(new_n986), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1961), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n970), .A2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G171), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1055), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1032), .A2(new_n1044), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1011), .A2(new_n999), .A3(new_n710), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(G1981), .B2(G305), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n984), .A2(new_n1014), .B1(new_n996), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G299), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n569), .A2(new_n573), .A3(new_n1061), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(new_n1065), .B(KEYINPUT119), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT56), .B(G2072), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n965), .B(new_n1067), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1068));
  INV_X1    g643(.A(G1956), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n970), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(new_n1065), .A3(new_n1070), .ZN(new_n1072));
  INV_X1    g647(.A(G1348), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n970), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n977), .A2(new_n930), .A3(new_n943), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n859), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1066), .A2(new_n1071), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n965), .B(new_n928), .C1(new_n1045), .C2(new_n1046), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n977), .A2(new_n943), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT120), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1080), .A2(new_n1084), .A3(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n555), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n599), .A2(new_n1090), .A3(new_n600), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1090), .B1(new_n599), .B2(new_n600), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1093), .A2(new_n1074), .A3(KEYINPUT60), .A4(new_n1075), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT60), .ZN(new_n1095));
  AOI21_X1  g670(.A(G1348), .B1(new_n974), .B2(new_n969), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1075), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1074), .A2(KEYINPUT60), .A3(new_n1075), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1092), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1094), .B(new_n1098), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1088), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n555), .B(new_n1102), .C1(new_n1079), .C2(new_n1086), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1089), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1065), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1072), .B1(new_n1105), .B2(KEYINPUT61), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT61), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1068), .A2(new_n1065), .A3(new_n1107), .A4(new_n1070), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1077), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n964), .B1(G164), .B2(new_n939), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n960), .A2(new_n943), .A3(new_n1050), .A4(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1049), .A2(new_n1112), .A3(G301), .A4(new_n1053), .ZN(new_n1113));
  AOI21_X1  g688(.A(KEYINPUT54), .B1(new_n1055), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1114), .A2(new_n1042), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1032), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1049), .A2(new_n1053), .A3(new_n1112), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(G171), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1049), .A2(G301), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT54), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1119), .B1(new_n1118), .B2(G171), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1117), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1121), .A2(KEYINPUT54), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT125), .A4(new_n1120), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1057), .B(new_n1060), .C1(new_n1116), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n946), .B1(new_n1031), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n944), .B1(new_n931), .B2(new_n771), .ZN(new_n1131));
  XNOR2_X1  g706(.A(new_n1131), .B(KEYINPUT126), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n944), .A2(G1996), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT46), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n1135), .B(KEYINPUT47), .Z(new_n1136));
  NOR2_X1   g711(.A1(new_n934), .A2(new_n944), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n944), .A2(new_n936), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(KEYINPUT48), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(KEYINPUT48), .B2(new_n1138), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n693), .A2(new_n696), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n932), .A2(new_n1141), .B1(G2067), .B2(new_n732), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n945), .ZN(new_n1143));
  AND3_X1   g718(.A1(new_n1136), .A2(new_n1140), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1130), .A2(new_n1144), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g720(.A(G319), .B1(new_n645), .B2(new_n646), .ZN(new_n1147));
  OR2_X1    g721(.A1(G227), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1149));
  AND2_X1   g723(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1151));
  NOR3_X1   g725(.A1(new_n1150), .A2(new_n1151), .A3(G229), .ZN(new_n1152));
  OAI211_X1 g726(.A(new_n855), .B(new_n1152), .C1(new_n913), .C2(new_n921), .ZN(G225));
  INV_X1    g727(.A(G225), .ZN(G308));
endmodule


