

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U551 ( .A(n762), .B(n761), .ZN(n767) );
  XNOR2_X1 U552 ( .A(n544), .B(KEYINPUT65), .ZN(G160) );
  NOR2_X1 U553 ( .A1(n781), .A2(n921), .ZN(n749) );
  NOR2_X1 U554 ( .A1(n757), .A2(G299), .ZN(n752) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n776) );
  INV_X1 U556 ( .A(KEYINPUT29), .ZN(n761) );
  XNOR2_X1 U557 ( .A(n776), .B(KEYINPUT31), .ZN(n777) );
  XNOR2_X1 U558 ( .A(n778), .B(n777), .ZN(n779) );
  NOR2_X1 U559 ( .A1(G1966), .A2(n811), .ZN(n792) );
  NAND2_X1 U560 ( .A1(n730), .A2(n729), .ZN(n781) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n638) );
  NOR2_X2 U562 ( .A1(n531), .A2(n529), .ZN(n877) );
  NOR2_X1 U563 ( .A1(G651), .A2(n656), .ZN(n650) );
  XOR2_X1 U564 ( .A(KEYINPUT1), .B(n520), .Z(n655) );
  NOR2_X1 U565 ( .A1(n536), .A2(n535), .ZN(G164) );
  NAND2_X1 U566 ( .A1(G91), .A2(n638), .ZN(n518) );
  XOR2_X1 U567 ( .A(KEYINPUT0), .B(G543), .Z(n656) );
  INV_X1 U568 ( .A(G651), .ZN(n519) );
  NOR2_X1 U569 ( .A1(n656), .A2(n519), .ZN(n641) );
  NAND2_X1 U570 ( .A1(G78), .A2(n641), .ZN(n517) );
  NAND2_X1 U571 ( .A1(n518), .A2(n517), .ZN(n524) );
  NOR2_X1 U572 ( .A1(G543), .A2(n519), .ZN(n520) );
  NAND2_X1 U573 ( .A1(G65), .A2(n655), .ZN(n522) );
  NAND2_X1 U574 ( .A1(G53), .A2(n650), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n523) );
  OR2_X1 U576 ( .A1(n524), .A2(n523), .ZN(G299) );
  NOR2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n525), .Z(n873) );
  NAND2_X1 U579 ( .A1(G138), .A2(n873), .ZN(n527) );
  INV_X1 U580 ( .A(G2104), .ZN(n529) );
  NOR2_X2 U581 ( .A1(G2105), .A2(n529), .ZN(n874) );
  NAND2_X1 U582 ( .A1(G102), .A2(n874), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U584 ( .A(KEYINPUT86), .B(n528), .ZN(n536) );
  INV_X1 U585 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n877), .A2(G114), .ZN(n530) );
  XNOR2_X1 U587 ( .A(n530), .B(KEYINPUT84), .ZN(n533) );
  NOR2_X1 U588 ( .A1(G2104), .A2(n531), .ZN(n878) );
  NAND2_X1 U589 ( .A1(G126), .A2(n878), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT85), .B(n534), .Z(n535) );
  NAND2_X1 U592 ( .A1(G137), .A2(n873), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G113), .A2(n877), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G125), .A2(n878), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n541) );
  NAND2_X1 U596 ( .A1(G101), .A2(n874), .ZN(n539) );
  XNOR2_X1 U597 ( .A(KEYINPUT23), .B(n539), .ZN(n540) );
  NOR2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n638), .A2(G89), .ZN(n545) );
  XNOR2_X1 U601 ( .A(KEYINPUT4), .B(n545), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n641), .A2(G76), .ZN(n546) );
  XOR2_X1 U603 ( .A(KEYINPUT71), .B(n546), .Z(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U605 ( .A(n549), .B(KEYINPUT5), .ZN(n554) );
  NAND2_X1 U606 ( .A1(G63), .A2(n655), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G51), .A2(n650), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U609 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(n555), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U613 ( .A(G2443), .B(G2446), .Z(n557) );
  XNOR2_X1 U614 ( .A(G2427), .B(G2451), .ZN(n556) );
  XNOR2_X1 U615 ( .A(n557), .B(n556), .ZN(n563) );
  XOR2_X1 U616 ( .A(G2430), .B(G2454), .Z(n559) );
  XNOR2_X1 U617 ( .A(G1341), .B(G1348), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U619 ( .A(G2435), .B(G2438), .Z(n560) );
  XNOR2_X1 U620 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U621 ( .A(n563), .B(n562), .Z(n564) );
  AND2_X1 U622 ( .A1(G14), .A2(n564), .ZN(G401) );
  AND2_X1 U623 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U624 ( .A(G132), .ZN(G219) );
  INV_X1 U625 ( .A(G82), .ZN(G220) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G120), .ZN(G236) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n565) );
  XNOR2_X1 U629 ( .A(n565), .B(KEYINPUT10), .ZN(n566) );
  XNOR2_X1 U630 ( .A(KEYINPUT68), .B(n566), .ZN(G223) );
  INV_X1 U631 ( .A(G223), .ZN(n831) );
  NAND2_X1 U632 ( .A1(n831), .A2(G567), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT11), .B(n567), .Z(G234) );
  XNOR2_X1 U634 ( .A(KEYINPUT69), .B(KEYINPUT70), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n638), .A2(G81), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n568), .B(KEYINPUT12), .ZN(n570) );
  NAND2_X1 U637 ( .A1(G68), .A2(n641), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n571), .B(KEYINPUT13), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n655), .A2(G56), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n574), .B(KEYINPUT14), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G43), .A2(n650), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n959) );
  NAND2_X1 U646 ( .A1(n959), .A2(G860), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G90), .A2(n638), .ZN(n580) );
  NAND2_X1 U648 ( .A1(G77), .A2(n641), .ZN(n579) );
  NAND2_X1 U649 ( .A1(n580), .A2(n579), .ZN(n582) );
  XOR2_X1 U650 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n581) );
  XNOR2_X1 U651 ( .A(n582), .B(n581), .ZN(n586) );
  NAND2_X1 U652 ( .A1(G64), .A2(n655), .ZN(n584) );
  NAND2_X1 U653 ( .A1(G52), .A2(n650), .ZN(n583) );
  AND2_X1 U654 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U655 ( .A1(n586), .A2(n585), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G66), .A2(n655), .ZN(n588) );
  NAND2_X1 U658 ( .A1(G54), .A2(n650), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U660 ( .A1(G92), .A2(n638), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G79), .A2(n641), .ZN(n589) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U664 ( .A(n593), .B(KEYINPUT15), .ZN(n972) );
  INV_X1 U665 ( .A(G868), .ZN(n668) );
  NAND2_X1 U666 ( .A1(n972), .A2(n668), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G284) );
  NOR2_X1 U668 ( .A1(G286), .A2(n668), .ZN(n597) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n596) );
  NOR2_X1 U670 ( .A1(n597), .A2(n596), .ZN(G297) );
  INV_X1 U671 ( .A(G860), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n598), .A2(G559), .ZN(n599) );
  INV_X1 U673 ( .A(n972), .ZN(n621) );
  NAND2_X1 U674 ( .A1(n599), .A2(n621), .ZN(n600) );
  XNOR2_X1 U675 ( .A(n600), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U676 ( .A1(n621), .A2(G868), .ZN(n601) );
  NOR2_X1 U677 ( .A1(G559), .A2(n601), .ZN(n603) );
  AND2_X1 U678 ( .A1(n668), .A2(n959), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G282) );
  XOR2_X1 U680 ( .A(G2100), .B(KEYINPUT74), .Z(n614) );
  NAND2_X1 U681 ( .A1(G123), .A2(n878), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n877), .A2(G111), .ZN(n605) );
  XNOR2_X1 U684 ( .A(n605), .B(KEYINPUT72), .ZN(n607) );
  NAND2_X1 U685 ( .A1(G135), .A2(n873), .ZN(n606) );
  NAND2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U687 ( .A1(G99), .A2(n874), .ZN(n608) );
  XNOR2_X1 U688 ( .A(KEYINPUT73), .B(n608), .ZN(n609) );
  NOR2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n918) );
  XOR2_X1 U691 ( .A(G2096), .B(n918), .Z(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U693 ( .A1(G93), .A2(n638), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G80), .A2(n641), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U696 ( .A1(G67), .A2(n655), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G55), .A2(n650), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  OR2_X1 U699 ( .A1(n620), .A2(n619), .ZN(n669) );
  NAND2_X1 U700 ( .A1(G559), .A2(n621), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n622), .B(n959), .ZN(n666) );
  XNOR2_X1 U702 ( .A(KEYINPUT75), .B(n666), .ZN(n623) );
  NOR2_X1 U703 ( .A1(G860), .A2(n623), .ZN(n624) );
  XOR2_X1 U704 ( .A(n669), .B(n624), .Z(G145) );
  NAND2_X1 U705 ( .A1(G88), .A2(n638), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G75), .A2(n641), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U708 ( .A1(G62), .A2(n655), .ZN(n628) );
  NAND2_X1 U709 ( .A1(G50), .A2(n650), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U711 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U712 ( .A1(G85), .A2(n638), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G72), .A2(n641), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n650), .A2(G47), .ZN(n633) );
  XOR2_X1 U716 ( .A(KEYINPUT66), .B(n633), .Z(n634) );
  NOR2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n655), .A2(G60), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(G290) );
  NAND2_X1 U720 ( .A1(n655), .A2(G61), .ZN(n640) );
  NAND2_X1 U721 ( .A1(n638), .A2(G86), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(n646) );
  XOR2_X1 U723 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n643) );
  NAND2_X1 U724 ( .A1(G73), .A2(n641), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n643), .B(n642), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT77), .B(n644), .Z(n645) );
  NOR2_X1 U727 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n647), .Z(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(G48), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(G305) );
  NAND2_X1 U731 ( .A1(G49), .A2(n650), .ZN(n652) );
  NAND2_X1 U732 ( .A1(G74), .A2(G651), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(KEYINPUT76), .B(n653), .ZN(n654) );
  NOR2_X1 U735 ( .A1(n655), .A2(n654), .ZN(n658) );
  NAND2_X1 U736 ( .A1(n656), .A2(G87), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(G288) );
  XOR2_X1 U738 ( .A(n669), .B(G299), .Z(n659) );
  XNOR2_X1 U739 ( .A(G166), .B(n659), .ZN(n663) );
  XNOR2_X1 U740 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n661) );
  XNOR2_X1 U741 ( .A(G290), .B(KEYINPUT81), .ZN(n660) );
  XNOR2_X1 U742 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U743 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U744 ( .A(n664), .B(G305), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(G288), .ZN(n897) );
  XOR2_X1 U746 ( .A(n897), .B(n666), .Z(n667) );
  NOR2_X1 U747 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U748 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U749 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n673), .ZN(n675) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(KEYINPUT82), .ZN(n674) );
  XNOR2_X1 U754 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U755 ( .A1(G2072), .A2(n676), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G236), .A2(G237), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G69), .A2(n677), .ZN(n678) );
  XNOR2_X1 U759 ( .A(KEYINPUT83), .B(n678), .ZN(n679) );
  NAND2_X1 U760 ( .A1(n679), .A2(G108), .ZN(n835) );
  NAND2_X1 U761 ( .A1(n835), .A2(G567), .ZN(n684) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U764 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U765 ( .A1(G96), .A2(n682), .ZN(n836) );
  NAND2_X1 U766 ( .A1(n836), .A2(G2106), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n684), .A2(n683), .ZN(n854) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U769 ( .A1(n854), .A2(n685), .ZN(n834) );
  NAND2_X1 U770 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U771 ( .A(G166), .ZN(G303) );
  INV_X1 U772 ( .A(G301), .ZN(G171) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n730) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n728) );
  NOR2_X1 U775 ( .A1(n730), .A2(n728), .ZN(n686) );
  XOR2_X1 U776 ( .A(KEYINPUT88), .B(n686), .Z(n823) );
  XOR2_X1 U777 ( .A(G2067), .B(KEYINPUT37), .Z(n697) );
  NAND2_X1 U778 ( .A1(G116), .A2(n877), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G128), .A2(n878), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U781 ( .A(n689), .B(KEYINPUT35), .ZN(n695) );
  XNOR2_X1 U782 ( .A(KEYINPUT89), .B(KEYINPUT34), .ZN(n693) );
  NAND2_X1 U783 ( .A1(G140), .A2(n873), .ZN(n691) );
  NAND2_X1 U784 ( .A1(G104), .A2(n874), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U786 ( .A(n693), .B(n692), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U788 ( .A(KEYINPUT36), .B(n696), .ZN(n893) );
  NOR2_X1 U789 ( .A1(n697), .A2(n893), .ZN(n932) );
  NAND2_X1 U790 ( .A1(n697), .A2(n893), .ZN(n929) );
  NOR2_X1 U791 ( .A1(n929), .A2(n823), .ZN(n698) );
  XNOR2_X1 U792 ( .A(n698), .B(KEYINPUT90), .ZN(n819) );
  NAND2_X1 U793 ( .A1(G117), .A2(n877), .ZN(n700) );
  NAND2_X1 U794 ( .A1(G129), .A2(n878), .ZN(n699) );
  NAND2_X1 U795 ( .A1(n700), .A2(n699), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G105), .A2(n874), .ZN(n701) );
  XNOR2_X1 U797 ( .A(n701), .B(KEYINPUT38), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n702), .B(KEYINPUT93), .ZN(n703) );
  NOR2_X1 U799 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U800 ( .A1(n873), .A2(G141), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n888) );
  NOR2_X1 U802 ( .A1(G1996), .A2(n888), .ZN(n912) );
  NAND2_X1 U803 ( .A1(G107), .A2(n877), .ZN(n708) );
  NAND2_X1 U804 ( .A1(G119), .A2(n878), .ZN(n707) );
  NAND2_X1 U805 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U806 ( .A(KEYINPUT91), .B(n709), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G131), .A2(n873), .ZN(n711) );
  NAND2_X1 U808 ( .A1(G95), .A2(n874), .ZN(n710) );
  AND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U810 ( .A1(n713), .A2(n712), .ZN(n885) );
  NAND2_X1 U811 ( .A1(G1991), .A2(n885), .ZN(n714) );
  XNOR2_X1 U812 ( .A(n714), .B(KEYINPUT92), .ZN(n716) );
  NAND2_X1 U813 ( .A1(G1996), .A2(n888), .ZN(n715) );
  NAND2_X1 U814 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U815 ( .A(KEYINPUT94), .B(n717), .Z(n925) );
  NOR2_X1 U816 ( .A1(n823), .A2(n925), .ZN(n820) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n718) );
  XOR2_X1 U818 ( .A(n718), .B(KEYINPUT105), .Z(n719) );
  NOR2_X1 U819 ( .A1(G1991), .A2(n885), .ZN(n917) );
  NOR2_X1 U820 ( .A1(n719), .A2(n917), .ZN(n720) );
  NOR2_X1 U821 ( .A1(n820), .A2(n720), .ZN(n721) );
  NOR2_X1 U822 ( .A1(n912), .A2(n721), .ZN(n722) );
  XOR2_X1 U823 ( .A(KEYINPUT39), .B(n722), .Z(n723) );
  NOR2_X1 U824 ( .A1(n819), .A2(n723), .ZN(n724) );
  XNOR2_X1 U825 ( .A(n724), .B(KEYINPUT106), .ZN(n725) );
  NOR2_X1 U826 ( .A1(n932), .A2(n725), .ZN(n726) );
  NOR2_X1 U827 ( .A1(n823), .A2(n726), .ZN(n727) );
  XNOR2_X1 U828 ( .A(n727), .B(KEYINPUT107), .ZN(n829) );
  INV_X1 U829 ( .A(n728), .ZN(n729) );
  NAND2_X1 U830 ( .A1(G8), .A2(n781), .ZN(n811) );
  NOR2_X1 U831 ( .A1(G1981), .A2(G305), .ZN(n731) );
  XOR2_X1 U832 ( .A(n731), .B(KEYINPUT24), .Z(n732) );
  NOR2_X1 U833 ( .A1(n811), .A2(n732), .ZN(n802) );
  NAND2_X1 U834 ( .A1(G1348), .A2(n972), .ZN(n976) );
  XOR2_X1 U835 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n735) );
  NOR2_X1 U836 ( .A1(G1341), .A2(n735), .ZN(n733) );
  NAND2_X1 U837 ( .A1(n976), .A2(n733), .ZN(n734) );
  NAND2_X1 U838 ( .A1(n734), .A2(n781), .ZN(n740) );
  NAND2_X1 U839 ( .A1(n972), .A2(G2067), .ZN(n737) );
  INV_X1 U840 ( .A(n735), .ZN(n741) );
  NAND2_X1 U841 ( .A1(G1996), .A2(n741), .ZN(n736) );
  NAND2_X1 U842 ( .A1(n737), .A2(n736), .ZN(n738) );
  INV_X1 U843 ( .A(n781), .ZN(n763) );
  NAND2_X1 U844 ( .A1(n738), .A2(n763), .ZN(n739) );
  NAND2_X1 U845 ( .A1(n740), .A2(n739), .ZN(n743) );
  NOR2_X1 U846 ( .A1(G1996), .A2(n741), .ZN(n742) );
  NOR2_X1 U847 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U848 ( .A1(n959), .A2(n744), .ZN(n756) );
  NAND2_X1 U849 ( .A1(G1348), .A2(n781), .ZN(n746) );
  NAND2_X1 U850 ( .A1(n763), .A2(G2067), .ZN(n745) );
  NAND2_X1 U851 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U852 ( .A1(n972), .A2(n747), .ZN(n754) );
  INV_X1 U853 ( .A(G2072), .ZN(n921) );
  XOR2_X1 U854 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n748) );
  XNOR2_X1 U855 ( .A(n749), .B(n748), .ZN(n751) );
  NAND2_X1 U856 ( .A1(n781), .A2(G1956), .ZN(n750) );
  NAND2_X1 U857 ( .A1(n751), .A2(n750), .ZN(n757) );
  XNOR2_X1 U858 ( .A(n752), .B(KEYINPUT98), .ZN(n753) );
  NOR2_X1 U859 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U860 ( .A1(n756), .A2(n755), .ZN(n760) );
  NAND2_X1 U861 ( .A1(G299), .A2(n757), .ZN(n758) );
  XNOR2_X1 U862 ( .A(KEYINPUT28), .B(n758), .ZN(n759) );
  NAND2_X1 U863 ( .A1(n760), .A2(n759), .ZN(n762) );
  XNOR2_X1 U864 ( .A(G2078), .B(KEYINPUT25), .ZN(n940) );
  NOR2_X1 U865 ( .A1(n781), .A2(n940), .ZN(n765) );
  INV_X1 U866 ( .A(G1961), .ZN(n987) );
  NOR2_X1 U867 ( .A1(n763), .A2(n987), .ZN(n764) );
  NOR2_X1 U868 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U869 ( .A1(n768), .A2(G171), .ZN(n766) );
  NAND2_X1 U870 ( .A1(n767), .A2(n766), .ZN(n780) );
  OR2_X1 U871 ( .A1(G171), .A2(n768), .ZN(n769) );
  XNOR2_X1 U872 ( .A(n769), .B(KEYINPUT99), .ZN(n775) );
  NOR2_X1 U873 ( .A1(n781), .A2(G2084), .ZN(n770) );
  XNOR2_X1 U874 ( .A(n770), .B(KEYINPUT96), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n792), .A2(n789), .ZN(n771) );
  NAND2_X1 U876 ( .A1(G8), .A2(n771), .ZN(n772) );
  XNOR2_X1 U877 ( .A(KEYINPUT30), .B(n772), .ZN(n773) );
  NOR2_X1 U878 ( .A1(n773), .A2(G168), .ZN(n774) );
  NOR2_X1 U879 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U880 ( .A1(n780), .A2(n779), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n790), .A2(G286), .ZN(n786) );
  NOR2_X1 U882 ( .A1(G1971), .A2(n811), .ZN(n783) );
  NOR2_X1 U883 ( .A1(G2090), .A2(n781), .ZN(n782) );
  NOR2_X1 U884 ( .A1(n783), .A2(n782), .ZN(n784) );
  NAND2_X1 U885 ( .A1(G303), .A2(n784), .ZN(n785) );
  NAND2_X1 U886 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U887 ( .A1(n787), .A2(G8), .ZN(n788) );
  XNOR2_X1 U888 ( .A(KEYINPUT32), .B(n788), .ZN(n796) );
  NAND2_X1 U889 ( .A1(n789), .A2(G8), .ZN(n794) );
  INV_X1 U890 ( .A(n790), .ZN(n791) );
  NOR2_X1 U891 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n804) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n797) );
  NAND2_X1 U895 ( .A1(G8), .A2(n797), .ZN(n798) );
  NAND2_X1 U896 ( .A1(n804), .A2(n798), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n811), .A2(n799), .ZN(n800) );
  XOR2_X1 U898 ( .A(KEYINPUT104), .B(n800), .Z(n801) );
  NOR2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n818) );
  NAND2_X1 U900 ( .A1(G1976), .A2(G288), .ZN(n970) );
  NOR2_X1 U901 ( .A1(G1976), .A2(G288), .ZN(n810) );
  NOR2_X1 U902 ( .A1(G1971), .A2(G303), .ZN(n803) );
  NOR2_X1 U903 ( .A1(n810), .A2(n803), .ZN(n960) );
  NAND2_X1 U904 ( .A1(n804), .A2(n960), .ZN(n805) );
  NAND2_X1 U905 ( .A1(n970), .A2(n805), .ZN(n806) );
  NOR2_X1 U906 ( .A1(n811), .A2(n806), .ZN(n807) );
  NOR2_X1 U907 ( .A1(KEYINPUT33), .A2(n807), .ZN(n808) );
  XNOR2_X1 U908 ( .A(n808), .B(KEYINPUT101), .ZN(n816) );
  XOR2_X1 U909 ( .A(KEYINPUT103), .B(G1981), .Z(n809) );
  XNOR2_X1 U910 ( .A(G305), .B(n809), .ZN(n963) );
  NAND2_X1 U911 ( .A1(n810), .A2(KEYINPUT33), .ZN(n812) );
  NOR2_X1 U912 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U913 ( .A(KEYINPUT102), .B(n813), .ZN(n814) );
  NOR2_X1 U914 ( .A1(n963), .A2(n814), .ZN(n815) );
  NAND2_X1 U915 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n827) );
  NOR2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n821), .B(KEYINPUT95), .ZN(n825) );
  XNOR2_X1 U919 ( .A(KEYINPUT87), .B(G1986), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n822), .B(G290), .ZN(n967) );
  NOR2_X1 U921 ( .A1(n967), .A2(n823), .ZN(n824) );
  NOR2_X1 U922 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U928 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(G188) );
  XOR2_X1 U931 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  NOR2_X1 U934 ( .A1(n836), .A2(n835), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(G2096), .B(G2100), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT43), .B(G2090), .Z(n840) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2084), .B(G2078), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U945 ( .A(G1986), .B(G1966), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1976), .B(G1971), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(KEYINPUT41), .B(G1956), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1981), .B(G1961), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(G229) );
  INV_X1 U955 ( .A(n854), .ZN(G319) );
  NAND2_X1 U956 ( .A1(G124), .A2(n878), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U958 ( .A1(n877), .A2(G112), .ZN(n856) );
  NAND2_X1 U959 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G136), .A2(n873), .ZN(n859) );
  NAND2_X1 U961 ( .A1(G100), .A2(n874), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U963 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U964 ( .A1(G118), .A2(n877), .ZN(n863) );
  NAND2_X1 U965 ( .A1(G130), .A2(n878), .ZN(n862) );
  NAND2_X1 U966 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G142), .A2(n873), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G106), .A2(n874), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT108), .B(n866), .Z(n867) );
  XNOR2_X1 U971 ( .A(KEYINPUT45), .B(n867), .ZN(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(G160), .B(n870), .ZN(n892) );
  XNOR2_X1 U974 ( .A(KEYINPUT48), .B(KEYINPUT109), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n918), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U976 ( .A(n872), .B(n871), .ZN(n887) );
  NAND2_X1 U977 ( .A1(G139), .A2(n873), .ZN(n876) );
  NAND2_X1 U978 ( .A1(G103), .A2(n874), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G115), .A2(n877), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G127), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n920) );
  XOR2_X1 U985 ( .A(G164), .B(n920), .Z(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n888), .B(G162), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U992 ( .A1(G37), .A2(n895), .ZN(n896) );
  XNOR2_X1 U993 ( .A(KEYINPUT110), .B(n896), .ZN(G395) );
  XNOR2_X1 U994 ( .A(n897), .B(KEYINPUT111), .ZN(n899) );
  XNOR2_X1 U995 ( .A(n972), .B(G286), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U997 ( .A(n959), .B(G171), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U999 ( .A1(G37), .A2(n902), .ZN(G397) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n903) );
  XOR2_X1 U1001 ( .A(KEYINPUT112), .B(n903), .Z(n904) );
  XNOR2_X1 U1002 ( .A(KEYINPUT49), .B(n904), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n905) );
  XOR2_X1 U1004 ( .A(KEYINPUT113), .B(n905), .Z(n906) );
  NAND2_X1 U1005 ( .A1(G319), .A2(n906), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(G401), .A2(n907), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(n909), .A2(n908), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  INV_X1 U1010 ( .A(KEYINPUT55), .ZN(n936) );
  XOR2_X1 U1011 ( .A(KEYINPUT115), .B(KEYINPUT52), .Z(n910) );
  XNOR2_X1 U1012 ( .A(KEYINPUT116), .B(n910), .ZN(n934) );
  XNOR2_X1 U1013 ( .A(G160), .B(G2084), .ZN(n915) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n911) );
  NOR2_X1 U1015 ( .A1(n912), .A2(n911), .ZN(n913) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n913), .Z(n914) );
  NAND2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n928) );
  XOR2_X1 U1020 ( .A(G164), .B(G2078), .Z(n923) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n924), .B(KEYINPUT50), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1028 ( .A(n934), .B(n933), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n937), .A2(G29), .ZN(n1020) );
  XNOR2_X1 U1031 ( .A(G1996), .B(G32), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G2067), .B(G26), .ZN(n938) );
  NOR2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n944) );
  XOR2_X1 U1034 ( .A(n940), .B(G27), .Z(n942) );
  XNOR2_X1 U1035 ( .A(G2072), .B(G33), .ZN(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n949) );
  XNOR2_X1 U1038 ( .A(G1991), .B(KEYINPUT117), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n945), .B(G25), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(G28), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT118), .B(n947), .ZN(n948) );
  NOR2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1043 ( .A(KEYINPUT53), .B(n950), .Z(n954) );
  XNOR2_X1 U1044 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(n951), .B(G34), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G2084), .B(n952), .ZN(n953) );
  NAND2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G35), .B(G2090), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1050 ( .A(KEYINPUT55), .B(n957), .Z(n958) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n958), .ZN(n1016) );
  XOR2_X1 U1052 ( .A(G16), .B(KEYINPUT56), .Z(n986) );
  XNOR2_X1 U1053 ( .A(n959), .B(G1341), .ZN(n961) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n983) );
  XOR2_X1 U1055 ( .A(G1966), .B(G168), .Z(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT120), .B(n964), .Z(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT57), .B(n965), .ZN(n981) );
  NAND2_X1 U1059 ( .A1(G1971), .A2(G303), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(G1956), .B(G299), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(G301), .B(G1961), .ZN(n974) );
  NOR2_X1 U1065 ( .A1(n972), .A2(G1348), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1068 ( .A(KEYINPUT121), .B(n977), .Z(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1071 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(n984), .B(KEYINPUT122), .ZN(n985) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n1013) );
  XOR2_X1 U1074 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n1010) );
  XOR2_X1 U1075 ( .A(G1966), .B(G21), .Z(n989) );
  XNOR2_X1 U1076 ( .A(n987), .B(G5), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n996) );
  XNOR2_X1 U1078 ( .A(G1976), .B(G23), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(G1971), .B(G22), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n993) );
  XOR2_X1 U1081 ( .A(G1986), .B(G24), .Z(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(KEYINPUT58), .B(n994), .ZN(n995) );
  NOR2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1008) );
  XNOR2_X1 U1085 ( .A(G1981), .B(G6), .ZN(n998) );
  XNOR2_X1 U1086 ( .A(G20), .B(G1956), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1005) );
  XOR2_X1 U1088 ( .A(G4), .B(KEYINPUT124), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(n1000), .B(n999), .ZN(n1003) );
  XOR2_X1 U1091 ( .A(KEYINPUT123), .B(G1341), .Z(n1001) );
  XNOR2_X1 U1092 ( .A(G19), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1006), .Z(n1007) );
  NAND2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(G16), .A2(n1011), .ZN(n1012) );
  NOR2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1100 ( .A(KEYINPUT126), .B(n1014), .Z(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1102 ( .A1(G11), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1021), .Z(G311) );
  INV_X1 U1106 ( .A(G311), .ZN(G150) );
endmodule

