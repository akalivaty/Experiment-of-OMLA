

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786;

  AND2_X1 U387 ( .A1(n401), .A2(n402), .ZN(n400) );
  NAND2_X1 U388 ( .A1(n601), .A2(n591), .ZN(n593) );
  AND2_X1 U389 ( .A1(n403), .A2(n595), .ZN(n401) );
  INV_X1 U390 ( .A(G953), .ZN(n755) );
  XOR2_X1 U391 ( .A(n569), .B(KEYINPUT19), .Z(n365) );
  INV_X1 U392 ( .A(n537), .ZN(n406) );
  XNOR2_X2 U393 ( .A(n419), .B(KEYINPUT32), .ZN(n786) );
  NOR2_X1 U394 ( .A1(n664), .A2(n663), .ZN(n601) );
  XNOR2_X2 U395 ( .A(n393), .B(n554), .ZN(n781) );
  XNOR2_X2 U396 ( .A(n486), .B(n761), .ZN(n394) );
  INV_X1 U397 ( .A(n596), .ZN(n416) );
  NOR2_X1 U398 ( .A1(n561), .A2(n560), .ZN(n727) );
  XNOR2_X1 U399 ( .A(n457), .B(n398), .ZN(n596) );
  INV_X1 U400 ( .A(KEYINPUT35), .ZN(n412) );
  INV_X1 U401 ( .A(KEYINPUT74), .ZN(n367) );
  INV_X1 U402 ( .A(KEYINPUT66), .ZN(n417) );
  NOR2_X1 U403 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U404 ( .A1(n781), .A2(n783), .ZN(n556) );
  NAND2_X1 U405 ( .A1(n404), .A2(n537), .ZN(n399) );
  NAND2_X1 U406 ( .A1(n381), .A2(n416), .ZN(n600) );
  XNOR2_X1 U407 ( .A(n382), .B(n417), .ZN(n381) );
  NOR2_X1 U408 ( .A1(n493), .A2(n492), .ZN(n494) );
  AND2_X1 U409 ( .A1(n596), .A2(n466), .ZN(n605) );
  OR2_X1 U410 ( .A1(n713), .A2(G902), .ZN(n410) );
  NAND2_X1 U411 ( .A1(n400), .A2(n399), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n569), .B(KEYINPUT19), .ZN(n531) );
  BUF_X1 U413 ( .A(n418), .Z(n366) );
  XNOR2_X1 U414 ( .A(n494), .B(n367), .ZN(n550) );
  NOR2_X1 U415 ( .A1(n623), .A2(n436), .ZN(n369) );
  NAND2_X2 U416 ( .A1(n540), .A2(n653), .ZN(n569) );
  BUF_X1 U417 ( .A(n623), .Z(n368) );
  XNOR2_X2 U418 ( .A(n369), .B(n370), .ZN(n540) );
  XOR2_X1 U419 ( .A(n438), .B(KEYINPUT93), .Z(n370) );
  BUF_X1 U420 ( .A(n640), .Z(n756) );
  XNOR2_X1 U421 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n471) );
  XNOR2_X1 U422 ( .A(n414), .B(G134), .ZN(n481) );
  INV_X1 U423 ( .A(G131), .ZN(n414) );
  XNOR2_X1 U424 ( .A(n384), .B(KEYINPUT72), .ZN(n383) );
  AND2_X1 U425 ( .A1(n600), .A2(n396), .ZN(n395) );
  XNOR2_X1 U426 ( .A(G137), .B(G146), .ZN(n482) );
  XNOR2_X1 U427 ( .A(G116), .B(G113), .ZN(n432) );
  XNOR2_X1 U428 ( .A(KEYINPUT3), .B(G119), .ZN(n431) );
  XOR2_X1 U429 ( .A(G137), .B(G140), .Z(n461) );
  INV_X1 U430 ( .A(KEYINPUT11), .ZN(n509) );
  XOR2_X1 U431 ( .A(G140), .B(G122), .Z(n514) );
  XNOR2_X1 U432 ( .A(n481), .B(n413), .ZN(n769) );
  INV_X1 U433 ( .A(KEYINPUT95), .ZN(n413) );
  XNOR2_X1 U434 ( .A(G146), .B(G125), .ZN(n445) );
  NAND2_X1 U435 ( .A1(n576), .A2(n371), .ZN(n577) );
  XNOR2_X1 U436 ( .A(n389), .B(n541), .ZN(n657) );
  INV_X1 U437 ( .A(KEYINPUT109), .ZN(n541) );
  OR2_X1 U438 ( .A1(n549), .A2(n390), .ZN(n389) );
  XNOR2_X1 U439 ( .A(n520), .B(n519), .ZN(n553) );
  XNOR2_X1 U440 ( .A(KEYINPUT13), .B(G475), .ZN(n519) );
  XNOR2_X1 U441 ( .A(G128), .B(G119), .ZN(n446) );
  XNOR2_X1 U442 ( .A(n552), .B(n551), .ZN(n580) );
  INV_X1 U443 ( .A(KEYINPUT39), .ZN(n551) );
  XNOR2_X1 U444 ( .A(n458), .B(n375), .ZN(n398) );
  INV_X1 U445 ( .A(KEYINPUT22), .ZN(n409) );
  INV_X1 U446 ( .A(KEYINPUT46), .ZN(n555) );
  NAND2_X1 U447 ( .A1(n596), .A2(n590), .ZN(n663) );
  XNOR2_X1 U448 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n424) );
  XNOR2_X1 U449 ( .A(n485), .B(n484), .ZN(n487) );
  XNOR2_X1 U450 ( .A(G122), .B(G107), .ZN(n499) );
  XNOR2_X1 U451 ( .A(G116), .B(G134), .ZN(n495) );
  XNOR2_X1 U452 ( .A(n512), .B(n511), .ZN(n518) );
  XNOR2_X1 U453 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U454 ( .A(G146), .B(G107), .Z(n464) );
  XNOR2_X1 U455 ( .A(n542), .B(n422), .ZN(n687) );
  NOR2_X1 U456 ( .A1(n657), .A2(n656), .ZN(n542) );
  NOR2_X1 U457 ( .A1(n686), .A2(KEYINPUT34), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n447), .B(n373), .ZN(n455) );
  XNOR2_X1 U459 ( .A(n628), .B(KEYINPUT91), .ZN(n752) );
  XNOR2_X1 U460 ( .A(n392), .B(n391), .ZN(n783) );
  XNOR2_X1 U461 ( .A(n548), .B(KEYINPUT42), .ZN(n391) );
  NOR2_X1 U462 ( .A1(n687), .A2(n557), .ZN(n392) );
  INV_X1 U463 ( .A(KEYINPUT111), .ZN(n548) );
  NAND2_X1 U464 ( .A1(n580), .A2(n730), .ZN(n393) );
  NAND2_X1 U465 ( .A1(n408), .A2(n377), .ZN(n419) );
  INV_X1 U466 ( .A(n675), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n489), .B(G472), .ZN(n671) );
  XOR2_X1 U468 ( .A(n575), .B(KEYINPUT80), .Z(n371) );
  XOR2_X1 U469 ( .A(KEYINPUT23), .B(G110), .Z(n372) );
  XNOR2_X1 U470 ( .A(KEYINPUT24), .B(KEYINPUT76), .ZN(n373) );
  AND2_X1 U471 ( .A1(n564), .A2(n563), .ZN(n374) );
  XOR2_X1 U472 ( .A(KEYINPUT75), .B(KEYINPUT25), .Z(n375) );
  AND2_X1 U473 ( .A1(n664), .A2(n566), .ZN(n376) );
  AND2_X1 U474 ( .A1(n599), .A2(n598), .ZN(n377) );
  AND2_X1 U475 ( .A1(n610), .A2(n664), .ZN(n378) );
  AND2_X1 U476 ( .A1(n605), .A2(n566), .ZN(n379) );
  XOR2_X1 U477 ( .A(KEYINPUT88), .B(KEYINPUT0), .Z(n380) );
  NAND2_X1 U478 ( .A1(n408), .A2(n376), .ZN(n382) );
  XNOR2_X2 U479 ( .A(n538), .B(n409), .ZN(n408) );
  NAND2_X1 U480 ( .A1(n385), .A2(n383), .ZN(n617) );
  NAND2_X1 U481 ( .A1(n395), .A2(n366), .ZN(n384) );
  XNOR2_X1 U482 ( .A(n386), .B(n613), .ZN(n385) );
  NAND2_X1 U483 ( .A1(n387), .A2(n612), .ZN(n386) );
  NAND2_X1 U484 ( .A1(n397), .A2(KEYINPUT44), .ZN(n387) );
  XNOR2_X2 U485 ( .A(n388), .B(n423), .ZN(n486) );
  XNOR2_X1 U486 ( .A(n388), .B(n769), .ZN(n771) );
  XNOR2_X2 U487 ( .A(n498), .B(KEYINPUT4), .ZN(n388) );
  INV_X1 U488 ( .A(n549), .ZN(n654) );
  INV_X1 U489 ( .A(n653), .ZN(n390) );
  XNOR2_X1 U490 ( .A(n394), .B(n435), .ZN(n623) );
  XNOR2_X1 U491 ( .A(n394), .B(n411), .ZN(n713) );
  NAND2_X1 U492 ( .A1(n418), .A2(n600), .ZN(n397) );
  INV_X1 U493 ( .A(KEYINPUT44), .ZN(n396) );
  XNOR2_X1 U494 ( .A(n617), .B(n616), .ZN(n640) );
  NAND2_X1 U495 ( .A1(n686), .A2(KEYINPUT34), .ZN(n402) );
  NAND2_X1 U496 ( .A1(n406), .A2(KEYINPUT34), .ZN(n403) );
  XNOR2_X2 U497 ( .A(n405), .B(n412), .ZN(n420) );
  NAND2_X1 U498 ( .A1(n407), .A2(n537), .ZN(n604) );
  NAND2_X1 U499 ( .A1(n537), .A2(n379), .ZN(n724) );
  XNOR2_X2 U500 ( .A(n532), .B(n380), .ZN(n537) );
  NAND2_X1 U501 ( .A1(n408), .A2(n378), .ZN(n718) );
  XNOR2_X2 U502 ( .A(n410), .B(G469), .ZN(n546) );
  XNOR2_X1 U503 ( .A(n465), .B(n464), .ZN(n411) );
  INV_X1 U504 ( .A(n420), .ZN(n782) );
  XNOR2_X2 U505 ( .A(n415), .B(G143), .ZN(n498) );
  XNOR2_X2 U506 ( .A(G128), .B(KEYINPUT65), .ZN(n415) );
  AND2_X2 U507 ( .A1(n420), .A2(n786), .ZN(n418) );
  XNOR2_X1 U508 ( .A(n540), .B(KEYINPUT38), .ZN(n549) );
  AND2_X1 U509 ( .A1(n530), .A2(n529), .ZN(n421) );
  XNOR2_X1 U510 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n422) );
  NOR2_X1 U511 ( .A1(n730), .A2(n581), .ZN(n658) );
  INV_X1 U512 ( .A(KEYINPUT86), .ZN(n613) );
  XNOR2_X1 U513 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U514 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U515 ( .A(KEYINPUT70), .B(G101), .ZN(n423) );
  XNOR2_X1 U516 ( .A(G110), .B(G104), .ZN(n761) );
  XOR2_X1 U517 ( .A(KEYINPUT78), .B(KEYINPUT92), .Z(n427) );
  NAND2_X1 U518 ( .A1(G224), .A2(n755), .ZN(n425) );
  XNOR2_X1 U519 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U520 ( .A(n427), .B(n426), .ZN(n430) );
  XNOR2_X1 U521 ( .A(KEYINPUT77), .B(KEYINPUT89), .ZN(n428) );
  XNOR2_X1 U522 ( .A(n445), .B(n428), .ZN(n429) );
  XNOR2_X1 U523 ( .A(n430), .B(n429), .ZN(n434) );
  XNOR2_X1 U524 ( .A(n432), .B(n431), .ZN(n477) );
  XNOR2_X1 U525 ( .A(n499), .B(KEYINPUT16), .ZN(n433) );
  XNOR2_X1 U526 ( .A(n477), .B(n433), .ZN(n763) );
  XNOR2_X1 U527 ( .A(n434), .B(n763), .ZN(n435) );
  XNOR2_X1 U528 ( .A(KEYINPUT15), .B(G902), .ZN(n620) );
  INV_X1 U529 ( .A(n620), .ZN(n436) );
  INV_X1 U530 ( .A(G902), .ZN(n488) );
  INV_X1 U531 ( .A(G237), .ZN(n437) );
  NAND2_X1 U532 ( .A1(n488), .A2(n437), .ZN(n490) );
  NAND2_X1 U533 ( .A1(n490), .A2(G210), .ZN(n438) );
  NAND2_X1 U534 ( .A1(G952), .A2(n755), .ZN(n526) );
  INV_X1 U535 ( .A(n526), .ZN(n440) );
  NAND2_X1 U536 ( .A1(G953), .A2(G902), .ZN(n523) );
  NOR2_X1 U537 ( .A1(G900), .A2(n523), .ZN(n439) );
  NOR2_X1 U538 ( .A1(n440), .A2(n439), .ZN(n442) );
  NAND2_X1 U539 ( .A1(G234), .A2(G237), .ZN(n441) );
  XOR2_X1 U540 ( .A(n441), .B(KEYINPUT14), .Z(n522) );
  NOR2_X1 U541 ( .A1(n442), .A2(n522), .ZN(n544) );
  NAND2_X1 U542 ( .A1(n620), .A2(G234), .ZN(n444) );
  XNOR2_X1 U543 ( .A(KEYINPUT20), .B(KEYINPUT96), .ZN(n443) );
  XNOR2_X1 U544 ( .A(n444), .B(n443), .ZN(n459) );
  NAND2_X1 U545 ( .A1(G217), .A2(n459), .ZN(n458) );
  XNOR2_X1 U546 ( .A(n445), .B(KEYINPUT10), .ZN(n515) );
  XNOR2_X1 U547 ( .A(n461), .B(n515), .ZN(n770) );
  XNOR2_X1 U548 ( .A(n372), .B(n446), .ZN(n447) );
  INV_X1 U549 ( .A(KEYINPUT8), .ZN(n448) );
  NAND2_X1 U550 ( .A1(KEYINPUT82), .A2(n448), .ZN(n451) );
  INV_X1 U551 ( .A(KEYINPUT82), .ZN(n449) );
  NAND2_X1 U552 ( .A1(n449), .A2(KEYINPUT8), .ZN(n450) );
  NAND2_X1 U553 ( .A1(n451), .A2(n450), .ZN(n453) );
  NAND2_X1 U554 ( .A1(G234), .A2(n755), .ZN(n452) );
  XNOR2_X1 U555 ( .A(n453), .B(n452), .ZN(n502) );
  NAND2_X1 U556 ( .A1(G221), .A2(n502), .ZN(n454) );
  XNOR2_X1 U557 ( .A(n770), .B(n456), .ZN(n749) );
  NOR2_X1 U558 ( .A1(n749), .A2(G902), .ZN(n457) );
  NAND2_X1 U559 ( .A1(n459), .A2(G221), .ZN(n460) );
  XNOR2_X1 U560 ( .A(KEYINPUT21), .B(n460), .ZN(n666) );
  XNOR2_X1 U561 ( .A(n666), .B(KEYINPUT97), .ZN(n590) );
  NAND2_X1 U562 ( .A1(n755), .A2(G227), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U564 ( .A(n463), .B(n769), .Z(n465) );
  AND2_X1 U565 ( .A1(n590), .A2(n546), .ZN(n466) );
  NAND2_X1 U566 ( .A1(n544), .A2(n605), .ZN(n493) );
  INV_X1 U567 ( .A(KEYINPUT5), .ZN(n467) );
  NAND2_X1 U568 ( .A1(KEYINPUT100), .A2(n467), .ZN(n470) );
  INV_X1 U569 ( .A(KEYINPUT100), .ZN(n468) );
  NAND2_X1 U570 ( .A1(n468), .A2(KEYINPUT5), .ZN(n469) );
  NAND2_X1 U571 ( .A1(n470), .A2(n469), .ZN(n472) );
  XNOR2_X1 U572 ( .A(n472), .B(n471), .ZN(n474) );
  NOR2_X1 U573 ( .A1(G953), .A2(G237), .ZN(n506) );
  NAND2_X1 U574 ( .A1(n506), .A2(G210), .ZN(n473) );
  XNOR2_X1 U575 ( .A(n474), .B(n473), .ZN(n478) );
  INV_X1 U576 ( .A(n478), .ZN(n476) );
  INV_X1 U577 ( .A(n477), .ZN(n475) );
  NAND2_X1 U578 ( .A1(n476), .A2(n475), .ZN(n480) );
  NAND2_X1 U579 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U580 ( .A1(n480), .A2(n479), .ZN(n485) );
  INV_X1 U581 ( .A(n481), .ZN(n483) );
  XNOR2_X1 U582 ( .A(n487), .B(n486), .ZN(n633) );
  NAND2_X1 U583 ( .A1(n633), .A2(n488), .ZN(n489) );
  INV_X1 U584 ( .A(G472), .ZN(n632) );
  NAND2_X1 U585 ( .A1(n490), .A2(G214), .ZN(n653) );
  NAND2_X1 U586 ( .A1(n671), .A2(n653), .ZN(n491) );
  XNOR2_X1 U587 ( .A(n491), .B(KEYINPUT30), .ZN(n492) );
  XOR2_X1 U588 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n496) );
  XNOR2_X1 U589 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U590 ( .A(n497), .B(KEYINPUT103), .Z(n501) );
  XOR2_X1 U591 ( .A(n498), .B(n499), .Z(n500) );
  XNOR2_X1 U592 ( .A(n501), .B(n500), .ZN(n504) );
  NAND2_X1 U593 ( .A1(G217), .A2(n502), .ZN(n503) );
  XOR2_X1 U594 ( .A(n504), .B(n503), .Z(n744) );
  NOR2_X1 U595 ( .A1(n744), .A2(G902), .ZN(n505) );
  XOR2_X1 U596 ( .A(n505), .B(G478), .Z(n533) );
  XOR2_X1 U597 ( .A(KEYINPUT12), .B(KEYINPUT101), .Z(n508) );
  NAND2_X1 U598 ( .A1(G214), .A2(n506), .ZN(n507) );
  XNOR2_X1 U599 ( .A(n508), .B(n507), .ZN(n512) );
  XNOR2_X1 U600 ( .A(G143), .B(G113), .ZN(n510) );
  XNOR2_X1 U601 ( .A(G131), .B(G104), .ZN(n513) );
  XNOR2_X1 U602 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U603 ( .A(n516), .B(n515), .Z(n517) );
  XNOR2_X1 U604 ( .A(n518), .B(n517), .ZN(n705) );
  NOR2_X1 U605 ( .A1(G902), .A2(n705), .ZN(n520) );
  NAND2_X1 U606 ( .A1(n533), .A2(n553), .ZN(n594) );
  NOR2_X1 U607 ( .A1(n550), .A2(n594), .ZN(n521) );
  NAND2_X1 U608 ( .A1(n540), .A2(n521), .ZN(n573) );
  XNOR2_X1 U609 ( .A(n573), .B(G143), .ZN(G45) );
  INV_X1 U610 ( .A(n522), .ZN(n683) );
  OR2_X1 U611 ( .A1(n523), .A2(G898), .ZN(n525) );
  NOR2_X1 U612 ( .A1(KEYINPUT94), .A2(n525), .ZN(n524) );
  NAND2_X1 U613 ( .A1(n683), .A2(n524), .ZN(n530) );
  NAND2_X1 U614 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U615 ( .A1(n527), .A2(n683), .ZN(n528) );
  NAND2_X1 U616 ( .A1(n528), .A2(KEYINPUT94), .ZN(n529) );
  NAND2_X1 U617 ( .A1(n531), .A2(n421), .ZN(n532) );
  INV_X1 U618 ( .A(n553), .ZN(n534) );
  INV_X1 U619 ( .A(n533), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n534), .A2(n561), .ZN(n656) );
  INV_X1 U621 ( .A(n590), .ZN(n535) );
  NOR2_X1 U622 ( .A1(n656), .A2(n535), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U624 ( .A(KEYINPUT67), .B(KEYINPUT1), .ZN(n539) );
  XNOR2_X2 U625 ( .A(n546), .B(n539), .ZN(n664) );
  XNOR2_X1 U626 ( .A(n600), .B(G110), .ZN(G12) );
  NOR2_X1 U627 ( .A1(n666), .A2(n596), .ZN(n543) );
  NAND2_X1 U628 ( .A1(n544), .A2(n543), .ZN(n567) );
  NOR2_X1 U629 ( .A1(n566), .A2(n567), .ZN(n545) );
  XNOR2_X1 U630 ( .A(KEYINPUT28), .B(n545), .ZN(n547) );
  NAND2_X1 U631 ( .A1(n547), .A2(n546), .ZN(n557) );
  XOR2_X1 U632 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n554) );
  NOR2_X1 U633 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U634 ( .A(n553), .B(KEYINPUT102), .ZN(n560) );
  NAND2_X1 U635 ( .A1(n561), .A2(n560), .ZN(n734) );
  INV_X1 U636 ( .A(n734), .ZN(n730) );
  XNOR2_X1 U637 ( .A(n556), .B(n555), .ZN(n578) );
  NOR2_X1 U638 ( .A1(n557), .A2(n365), .ZN(n731) );
  INV_X1 U639 ( .A(KEYINPUT71), .ZN(n558) );
  NAND2_X1 U640 ( .A1(n731), .A2(n558), .ZN(n559) );
  XNOR2_X1 U641 ( .A(n559), .B(KEYINPUT47), .ZN(n564) );
  INV_X1 U642 ( .A(n727), .ZN(n738) );
  XOR2_X1 U643 ( .A(KEYINPUT104), .B(n738), .Z(n581) );
  XNOR2_X1 U644 ( .A(n658), .B(KEYINPUT81), .ZN(n607) );
  INV_X1 U645 ( .A(n607), .ZN(n562) );
  NAND2_X1 U646 ( .A1(n562), .A2(n731), .ZN(n563) );
  INV_X1 U647 ( .A(n671), .ZN(n566) );
  INV_X1 U648 ( .A(KEYINPUT6), .ZN(n565) );
  XNOR2_X1 U649 ( .A(n566), .B(n565), .ZN(n609) );
  INV_X1 U650 ( .A(n609), .ZN(n591) );
  NOR2_X1 U651 ( .A1(n734), .A2(n567), .ZN(n568) );
  NAND2_X1 U652 ( .A1(n591), .A2(n568), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n582), .A2(n569), .ZN(n571) );
  XNOR2_X1 U654 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n570) );
  XNOR2_X1 U655 ( .A(n571), .B(n570), .ZN(n572) );
  NOR2_X1 U656 ( .A1(n664), .A2(n572), .ZN(n740) );
  NOR2_X1 U657 ( .A1(n374), .A2(n740), .ZN(n576) );
  NAND2_X1 U658 ( .A1(n658), .A2(KEYINPUT47), .ZN(n574) );
  NAND2_X1 U659 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U660 ( .A(KEYINPUT48), .B(n579), .ZN(n589) );
  AND2_X1 U661 ( .A1(n581), .A2(n580), .ZN(n742) );
  INV_X1 U662 ( .A(n742), .ZN(n587) );
  INV_X1 U663 ( .A(n664), .ZN(n598) );
  NOR2_X1 U664 ( .A1(n598), .A2(n582), .ZN(n583) );
  NAND2_X1 U665 ( .A1(n583), .A2(n653), .ZN(n584) );
  XOR2_X1 U666 ( .A(KEYINPUT43), .B(n584), .Z(n585) );
  NOR2_X1 U667 ( .A1(n585), .A2(n540), .ZN(n586) );
  XNOR2_X1 U668 ( .A(n586), .B(KEYINPUT107), .ZN(n784) );
  AND2_X1 U669 ( .A1(n587), .A2(n784), .ZN(n588) );
  AND2_X2 U670 ( .A1(n589), .A2(n588), .ZN(n772) );
  XOR2_X1 U671 ( .A(KEYINPUT106), .B(KEYINPUT33), .Z(n592) );
  XNOR2_X2 U672 ( .A(n593), .B(n592), .ZN(n686) );
  INV_X1 U673 ( .A(n594), .ZN(n595) );
  XNOR2_X1 U674 ( .A(KEYINPUT79), .B(n609), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT105), .ZN(n667) );
  INV_X1 U676 ( .A(n667), .ZN(n608) );
  NOR2_X1 U677 ( .A1(n597), .A2(n608), .ZN(n599) );
  INV_X1 U678 ( .A(n601), .ZN(n602) );
  OR2_X1 U679 ( .A1(n566), .A2(n602), .ZN(n675) );
  INV_X1 U680 ( .A(KEYINPUT31), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n604), .B(n603), .ZN(n737) );
  NAND2_X1 U682 ( .A1(n737), .A2(n724), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n607), .A2(n606), .ZN(n611) );
  AND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  AND2_X1 U685 ( .A1(n611), .A2(n718), .ZN(n612) );
  XNOR2_X1 U686 ( .A(KEYINPUT85), .B(KEYINPUT45), .ZN(n615) );
  INV_X1 U687 ( .A(KEYINPUT64), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n615), .B(n614), .ZN(n616) );
  NAND2_X1 U689 ( .A1(n772), .A2(n640), .ZN(n647) );
  INV_X1 U690 ( .A(KEYINPUT2), .ZN(n641) );
  NOR2_X1 U691 ( .A1(n641), .A2(KEYINPUT73), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n647), .B(n618), .ZN(n622) );
  INV_X1 U693 ( .A(KEYINPUT73), .ZN(n644) );
  NOR2_X1 U694 ( .A1(n644), .A2(KEYINPUT2), .ZN(n619) );
  NOR2_X1 U695 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n703) );
  INV_X1 U697 ( .A(n703), .ZN(n712) );
  NAND2_X1 U698 ( .A1(n712), .A2(G210), .ZN(n626) );
  XNOR2_X1 U699 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n624) );
  XNOR2_X1 U700 ( .A(n368), .B(n624), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n626), .B(n625), .ZN(n629) );
  INV_X1 U702 ( .A(G952), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n627), .A2(G953), .ZN(n628) );
  INV_X1 U704 ( .A(n752), .ZN(n708) );
  NAND2_X1 U705 ( .A1(n629), .A2(n708), .ZN(n631) );
  INV_X1 U706 ( .A(KEYINPUT56), .ZN(n630) );
  XNOR2_X1 U707 ( .A(n631), .B(n630), .ZN(G51) );
  NOR2_X1 U708 ( .A1(n703), .A2(n632), .ZN(n635) );
  XOR2_X1 U709 ( .A(KEYINPUT62), .B(n633), .Z(n634) );
  XNOR2_X1 U710 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n636), .A2(n708), .ZN(n639) );
  XNOR2_X1 U712 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(KEYINPUT90), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n639), .B(n638), .ZN(G57) );
  NAND2_X1 U715 ( .A1(n647), .A2(KEYINPUT2), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n756), .A2(n641), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U719 ( .A1(KEYINPUT2), .A2(KEYINPUT73), .ZN(n646) );
  OR2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n648) );
  AND2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U722 ( .A1(n650), .A2(KEYINPUT83), .ZN(n694) );
  NOR2_X1 U723 ( .A1(KEYINPUT73), .A2(KEYINPUT2), .ZN(n651) );
  NAND2_X1 U724 ( .A1(n651), .A2(KEYINPUT83), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n756), .A2(n652), .ZN(n692) );
  NOR2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n660) );
  NOR2_X1 U728 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U730 ( .A(KEYINPUT121), .B(n661), .Z(n662) );
  NOR2_X1 U731 ( .A1(n686), .A2(n662), .ZN(n680) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U733 ( .A(n665), .B(KEYINPUT50), .ZN(n674) );
  XOR2_X1 U734 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n669) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U736 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(KEYINPUT120), .B(n672), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n677), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n687), .A2(n678), .ZN(n679) );
  NOR2_X1 U743 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U744 ( .A(n681), .B(KEYINPUT52), .ZN(n682) );
  XNOR2_X1 U745 ( .A(n682), .B(KEYINPUT122), .ZN(n685) );
  NAND2_X1 U746 ( .A1(G952), .A2(n683), .ZN(n684) );
  NOR2_X1 U747 ( .A1(n685), .A2(n684), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n688), .B(KEYINPUT123), .ZN(n689) );
  NAND2_X1 U750 ( .A1(n689), .A2(n755), .ZN(n690) );
  OR2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n697) );
  OR2_X1 U752 ( .A1(n692), .A2(n697), .ZN(n693) );
  OR2_X1 U753 ( .A1(n694), .A2(n693), .ZN(n699) );
  NOR2_X1 U754 ( .A1(n772), .A2(KEYINPUT2), .ZN(n695) );
  XOR2_X1 U755 ( .A(KEYINPUT84), .B(n695), .Z(n696) );
  OR2_X1 U756 ( .A1(n697), .A2(n696), .ZN(n698) );
  AND2_X1 U757 ( .A1(n699), .A2(n698), .ZN(n701) );
  INV_X1 U758 ( .A(KEYINPUT53), .ZN(n700) );
  XNOR2_X1 U759 ( .A(n701), .B(n700), .ZN(G75) );
  INV_X1 U760 ( .A(G475), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n707) );
  XOR2_X1 U762 ( .A(KEYINPUT68), .B(KEYINPUT59), .Z(n704) );
  XNOR2_X1 U763 ( .A(n705), .B(n704), .ZN(n706) );
  XNOR2_X1 U764 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U765 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U766 ( .A(KEYINPUT69), .B(KEYINPUT60), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n711), .B(n710), .ZN(G60) );
  BUF_X2 U768 ( .A(n712), .Z(n748) );
  NAND2_X1 U769 ( .A1(n748), .A2(G469), .ZN(n716) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n714) );
  XNOR2_X1 U771 ( .A(n713), .B(n714), .ZN(n715) );
  XNOR2_X1 U772 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n717), .A2(n752), .ZN(G54) );
  INV_X1 U774 ( .A(n718), .ZN(n719) );
  XNOR2_X1 U775 ( .A(G101), .B(n719), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n720), .B(KEYINPUT113), .ZN(G3) );
  NOR2_X1 U777 ( .A1(n734), .A2(n724), .ZN(n721) );
  XOR2_X1 U778 ( .A(G104), .B(n721), .Z(G6) );
  XOR2_X1 U779 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n723) );
  XNOR2_X1 U780 ( .A(G107), .B(KEYINPUT26), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n723), .B(n722), .ZN(n726) );
  NOR2_X1 U782 ( .A1(n738), .A2(n724), .ZN(n725) );
  XOR2_X1 U783 ( .A(n726), .B(n725), .Z(G9) );
  XOR2_X1 U784 ( .A(G128), .B(KEYINPUT29), .Z(n729) );
  NAND2_X1 U785 ( .A1(n731), .A2(n727), .ZN(n728) );
  XNOR2_X1 U786 ( .A(n729), .B(n728), .ZN(G30) );
  XOR2_X1 U787 ( .A(G146), .B(KEYINPUT115), .Z(n733) );
  NAND2_X1 U788 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U789 ( .A(n733), .B(n732), .ZN(G48) );
  NOR2_X1 U790 ( .A1(n734), .A2(n737), .ZN(n735) );
  XOR2_X1 U791 ( .A(KEYINPUT116), .B(n735), .Z(n736) );
  XNOR2_X1 U792 ( .A(G113), .B(n736), .ZN(G15) );
  NOR2_X1 U793 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U794 ( .A(G116), .B(n739), .Z(G18) );
  XNOR2_X1 U795 ( .A(G125), .B(n740), .ZN(n741) );
  XNOR2_X1 U796 ( .A(n741), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U797 ( .A(G134), .B(n742), .ZN(n743) );
  XNOR2_X1 U798 ( .A(n743), .B(KEYINPUT117), .ZN(G36) );
  NAND2_X1 U799 ( .A1(n748), .A2(G478), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n744), .B(KEYINPUT124), .ZN(n745) );
  XNOR2_X1 U801 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U802 ( .A1(n752), .A2(n747), .ZN(G63) );
  NAND2_X1 U803 ( .A1(n748), .A2(G217), .ZN(n750) );
  XNOR2_X1 U804 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(G66) );
  INV_X1 U806 ( .A(G898), .ZN(n760) );
  NAND2_X1 U807 ( .A1(G953), .A2(G224), .ZN(n753) );
  XOR2_X1 U808 ( .A(KEYINPUT61), .B(n753), .Z(n754) );
  NOR2_X1 U809 ( .A1(n760), .A2(n754), .ZN(n759) );
  NAND2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(KEYINPUT125), .ZN(n758) );
  NOR2_X1 U812 ( .A1(n759), .A2(n758), .ZN(n768) );
  NAND2_X1 U813 ( .A1(n760), .A2(G953), .ZN(n765) );
  XOR2_X1 U814 ( .A(G101), .B(n761), .Z(n762) );
  XNOR2_X1 U815 ( .A(n763), .B(n762), .ZN(n764) );
  NAND2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U817 ( .A(n766), .B(KEYINPUT126), .ZN(n767) );
  XNOR2_X1 U818 ( .A(n768), .B(n767), .ZN(G69) );
  XNOR2_X1 U819 ( .A(n771), .B(n770), .ZN(n776) );
  INV_X1 U820 ( .A(n772), .ZN(n773) );
  XOR2_X1 U821 ( .A(n776), .B(n773), .Z(n774) );
  NOR2_X1 U822 ( .A1(G953), .A2(n774), .ZN(n775) );
  XNOR2_X1 U823 ( .A(n775), .B(KEYINPUT127), .ZN(n780) );
  XNOR2_X1 U824 ( .A(G227), .B(n776), .ZN(n777) );
  NAND2_X1 U825 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U826 ( .A1(n778), .A2(G953), .ZN(n779) );
  NAND2_X1 U827 ( .A1(n780), .A2(n779), .ZN(G72) );
  XOR2_X1 U828 ( .A(G131), .B(n781), .Z(G33) );
  XOR2_X1 U829 ( .A(n782), .B(G122), .Z(G24) );
  XOR2_X1 U830 ( .A(n783), .B(G137), .Z(G39) );
  XNOR2_X1 U831 ( .A(G140), .B(KEYINPUT118), .ZN(n785) );
  XNOR2_X1 U832 ( .A(n785), .B(n784), .ZN(G42) );
  XNOR2_X1 U833 ( .A(G119), .B(n786), .ZN(G21) );
endmodule

