

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U547 ( .A1(n520), .A2(G2105), .ZN(n885) );
  BUF_X2 U548 ( .A(n877), .Z(n515) );
  XOR2_X1 U549 ( .A(KEYINPUT17), .B(n519), .Z(n877) );
  AND2_X1 U550 ( .A1(n740), .A2(n739), .ZN(n742) );
  NOR2_X1 U551 ( .A1(n784), .A2(n797), .ZN(n785) );
  NOR2_X1 U552 ( .A1(G164), .A2(G1384), .ZN(n718) );
  XOR2_X1 U553 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  XNOR2_X1 U554 ( .A(n726), .B(KEYINPUT99), .ZN(n733) );
  INV_X1 U555 ( .A(KEYINPUT100), .ZN(n741) );
  XNOR2_X1 U556 ( .A(n742), .B(n741), .ZN(n746) );
  INV_X1 U557 ( .A(KEYINPUT31), .ZN(n760) );
  XNOR2_X1 U558 ( .A(n760), .B(KEYINPUT102), .ZN(n761) );
  XNOR2_X1 U559 ( .A(n762), .B(n761), .ZN(n763) );
  NOR2_X1 U560 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U561 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U562 ( .A(G651), .ZN(n535) );
  INV_X1 U563 ( .A(KEYINPUT77), .ZN(n604) );
  NOR2_X1 U564 ( .A1(n803), .A2(n802), .ZN(n805) );
  XNOR2_X1 U565 ( .A(KEYINPUT1), .B(n537), .ZN(n652) );
  XNOR2_X1 U566 ( .A(n604), .B(KEYINPUT6), .ZN(n605) );
  XNOR2_X1 U567 ( .A(n606), .B(n605), .ZN(n607) );
  NOR2_X1 U568 ( .A1(n532), .A2(n531), .ZN(G160) );
  INV_X1 U569 ( .A(G2104), .ZN(n520) );
  NAND2_X1 U570 ( .A1(G126), .A2(n885), .ZN(n517) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U572 ( .A1(G114), .A2(n882), .ZN(n516) );
  NAND2_X1 U573 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U574 ( .A(n518), .B(KEYINPUT90), .ZN(n524) );
  NOR2_X1 U575 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  NAND2_X1 U576 ( .A1(G138), .A2(n515), .ZN(n522) );
  NOR2_X4 U577 ( .A1(G2105), .A2(n520), .ZN(n878) );
  NAND2_X1 U578 ( .A1(G102), .A2(n878), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U581 ( .A1(G101), .A2(n878), .ZN(n525) );
  XOR2_X1 U582 ( .A(KEYINPUT23), .B(n525), .Z(n528) );
  NAND2_X1 U583 ( .A1(G113), .A2(n882), .ZN(n526) );
  XOR2_X1 U584 ( .A(KEYINPUT65), .B(n526), .Z(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n532) );
  NAND2_X1 U586 ( .A1(G125), .A2(n885), .ZN(n530) );
  NAND2_X1 U587 ( .A1(G137), .A2(n515), .ZN(n529) );
  NAND2_X1 U588 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U589 ( .A1(G543), .A2(G651), .ZN(n648) );
  NAND2_X1 U590 ( .A1(G85), .A2(n648), .ZN(n534) );
  NOR2_X1 U591 ( .A1(n634), .A2(n535), .ZN(n649) );
  NAND2_X1 U592 ( .A1(G72), .A2(n649), .ZN(n533) );
  NAND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n542) );
  NOR2_X1 U594 ( .A1(G543), .A2(n535), .ZN(n536) );
  XOR2_X1 U595 ( .A(KEYINPUT66), .B(n536), .Z(n537) );
  NAND2_X1 U596 ( .A1(G60), .A2(n652), .ZN(n540) );
  NOR2_X1 U597 ( .A1(n634), .A2(G651), .ZN(n538) );
  XNOR2_X2 U598 ( .A(KEYINPUT64), .B(n538), .ZN(n653) );
  NAND2_X1 U599 ( .A1(G47), .A2(n653), .ZN(n539) );
  NAND2_X1 U600 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U601 ( .A1(n542), .A2(n541), .ZN(G290) );
  XOR2_X1 U602 ( .A(G2430), .B(G2443), .Z(n544) );
  XNOR2_X1 U603 ( .A(KEYINPUT107), .B(G2451), .ZN(n543) );
  XNOR2_X1 U604 ( .A(n544), .B(n543), .ZN(n551) );
  XOR2_X1 U605 ( .A(G2435), .B(G2427), .Z(n546) );
  XNOR2_X1 U606 ( .A(G2446), .B(G2454), .ZN(n545) );
  XNOR2_X1 U607 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U608 ( .A(n547), .B(G2438), .Z(n549) );
  XNOR2_X1 U609 ( .A(G1341), .B(G1348), .ZN(n548) );
  XNOR2_X1 U610 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n551), .B(n550), .ZN(n552) );
  AND2_X1 U612 ( .A1(n552), .A2(G14), .ZN(G401) );
  NAND2_X1 U613 ( .A1(n885), .A2(G123), .ZN(n553) );
  XNOR2_X1 U614 ( .A(n553), .B(KEYINPUT18), .ZN(n555) );
  NAND2_X1 U615 ( .A1(G135), .A2(n515), .ZN(n554) );
  NAND2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U617 ( .A(KEYINPUT79), .B(n556), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G111), .A2(n882), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G99), .A2(n878), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT80), .B(n559), .Z(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n973) );
  XNOR2_X1 U623 ( .A(G2096), .B(n973), .ZN(n562) );
  OR2_X1 U624 ( .A1(G2100), .A2(n562), .ZN(G156) );
  INV_X1 U625 ( .A(G57), .ZN(G237) );
  NAND2_X1 U626 ( .A1(G94), .A2(G452), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U630 ( .A(G223), .ZN(n823) );
  NAND2_X1 U631 ( .A1(n823), .A2(G567), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U633 ( .A1(n648), .A2(G81), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U635 ( .A1(G68), .A2(n649), .ZN(n567) );
  NAND2_X1 U636 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U637 ( .A(KEYINPUT13), .B(n569), .ZN(n575) );
  NAND2_X1 U638 ( .A1(n652), .A2(G56), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT14), .B(n570), .Z(n573) );
  NAND2_X1 U640 ( .A1(G43), .A2(n653), .ZN(n571) );
  XNOR2_X1 U641 ( .A(KEYINPUT71), .B(n571), .ZN(n572) );
  NOR2_X1 U642 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n988) );
  XOR2_X1 U644 ( .A(G860), .B(KEYINPUT72), .Z(n619) );
  NOR2_X1 U645 ( .A1(n988), .A2(n619), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT73), .ZN(G153) );
  NAND2_X1 U647 ( .A1(G64), .A2(n652), .ZN(n577) );
  XNOR2_X1 U648 ( .A(KEYINPUT67), .B(n577), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G90), .A2(n648), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G77), .A2(n649), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT9), .B(n580), .Z(n581) );
  XNOR2_X1 U653 ( .A(KEYINPUT68), .B(n581), .ZN(n582) );
  NOR2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G52), .A2(n653), .ZN(n584) );
  NAND2_X1 U656 ( .A1(n585), .A2(n584), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U658 ( .A1(n652), .A2(G66), .ZN(n592) );
  NAND2_X1 U659 ( .A1(G92), .A2(n648), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G79), .A2(n649), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n653), .A2(G54), .ZN(n588) );
  XOR2_X1 U663 ( .A(KEYINPUT74), .B(n588), .Z(n589) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X2 U665 ( .A(n593), .B(KEYINPUT15), .ZN(n1001) );
  OR2_X1 U666 ( .A1(n1001), .A2(G868), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n595), .A2(n594), .ZN(G284) );
  XNOR2_X1 U668 ( .A(KEYINPUT5), .B(KEYINPUT75), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n648), .A2(G89), .ZN(n596) );
  XNOR2_X1 U670 ( .A(n596), .B(KEYINPUT4), .ZN(n598) );
  NAND2_X1 U671 ( .A1(G76), .A2(n649), .ZN(n597) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n600), .B(n599), .ZN(n608) );
  NAND2_X1 U674 ( .A1(G63), .A2(n652), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT76), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G51), .A2(n653), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n606) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U679 ( .A(KEYINPUT7), .B(n609), .Z(G168) );
  XOR2_X1 U680 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U681 ( .A1(G91), .A2(n648), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G65), .A2(n652), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n649), .A2(G78), .ZN(n612) );
  XOR2_X1 U685 ( .A(KEYINPUT70), .B(n612), .Z(n613) );
  NOR2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G53), .A2(n653), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(G299) );
  INV_X1 U689 ( .A(G868), .ZN(n667) );
  NOR2_X1 U690 ( .A1(G286), .A2(n667), .ZN(n618) );
  NOR2_X1 U691 ( .A1(G868), .A2(G299), .ZN(n617) );
  NOR2_X1 U692 ( .A1(n618), .A2(n617), .ZN(G297) );
  NAND2_X1 U693 ( .A1(n619), .A2(G559), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n620), .A2(n1001), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT16), .ZN(n622) );
  XNOR2_X1 U696 ( .A(KEYINPUT78), .B(n622), .ZN(G148) );
  NOR2_X1 U697 ( .A1(G868), .A2(n988), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G868), .A2(n1001), .ZN(n623) );
  NOR2_X1 U699 ( .A1(G559), .A2(n623), .ZN(n624) );
  NOR2_X1 U700 ( .A1(n625), .A2(n624), .ZN(G282) );
  NAND2_X1 U701 ( .A1(G62), .A2(n652), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G50), .A2(n653), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U704 ( .A(KEYINPUT84), .B(n628), .Z(n632) );
  NAND2_X1 U705 ( .A1(G88), .A2(n648), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G75), .A2(n649), .ZN(n629) );
  AND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(G303) );
  INV_X1 U709 ( .A(G303), .ZN(G166) );
  NAND2_X1 U710 ( .A1(n653), .A2(G49), .ZN(n633) );
  XNOR2_X1 U711 ( .A(n633), .B(KEYINPUT82), .ZN(n639) );
  NAND2_X1 U712 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U713 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U715 ( .A1(n652), .A2(n637), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U717 ( .A(KEYINPUT83), .B(n640), .Z(G288) );
  NAND2_X1 U718 ( .A1(G86), .A2(n648), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G61), .A2(n652), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n649), .A2(G73), .ZN(n643) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U723 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U724 ( .A1(G48), .A2(n653), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(G305) );
  XNOR2_X1 U726 ( .A(G166), .B(G288), .ZN(n664) );
  NAND2_X1 U727 ( .A1(G93), .A2(n648), .ZN(n651) );
  NAND2_X1 U728 ( .A1(G80), .A2(n649), .ZN(n650) );
  NAND2_X1 U729 ( .A1(n651), .A2(n650), .ZN(n657) );
  NAND2_X1 U730 ( .A1(G67), .A2(n652), .ZN(n655) );
  NAND2_X1 U731 ( .A1(G55), .A2(n653), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U733 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U734 ( .A(KEYINPUT81), .B(n658), .Z(n830) );
  XNOR2_X1 U735 ( .A(KEYINPUT19), .B(n830), .ZN(n660) );
  XNOR2_X1 U736 ( .A(G290), .B(KEYINPUT85), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(n661) );
  XOR2_X1 U738 ( .A(n661), .B(G299), .Z(n662) );
  XNOR2_X1 U739 ( .A(G305), .B(n662), .ZN(n663) );
  XNOR2_X1 U740 ( .A(n664), .B(n663), .ZN(n896) );
  NAND2_X1 U741 ( .A1(G559), .A2(n1001), .ZN(n665) );
  XNOR2_X1 U742 ( .A(n988), .B(n665), .ZN(n829) );
  XNOR2_X1 U743 ( .A(n896), .B(n829), .ZN(n666) );
  NOR2_X1 U744 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U745 ( .A1(n830), .A2(G868), .ZN(n668) );
  NOR2_X1 U746 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U747 ( .A(KEYINPUT86), .B(n670), .Z(G295) );
  NAND2_X1 U748 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n671), .Z(n672) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n672), .ZN(n673) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n673), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n674), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n675) );
  NOR2_X1 U755 ( .A1(G237), .A2(n675), .ZN(n676) );
  NAND2_X1 U756 ( .A1(G108), .A2(n676), .ZN(n828) );
  NAND2_X1 U757 ( .A1(n828), .A2(G567), .ZN(n683) );
  XOR2_X1 U758 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n678) );
  NAND2_X1 U759 ( .A1(G132), .A2(G82), .ZN(n677) );
  XNOR2_X1 U760 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U761 ( .A1(n679), .A2(G218), .ZN(n680) );
  NAND2_X1 U762 ( .A1(G96), .A2(n680), .ZN(n827) );
  NAND2_X1 U763 ( .A1(G2106), .A2(n827), .ZN(n681) );
  XNOR2_X1 U764 ( .A(KEYINPUT88), .B(n681), .ZN(n682) );
  NAND2_X1 U765 ( .A1(n683), .A2(n682), .ZN(n832) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U767 ( .A1(n832), .A2(n684), .ZN(n826) );
  NAND2_X1 U768 ( .A1(n826), .A2(G36), .ZN(n685) );
  XOR2_X1 U769 ( .A(KEYINPUT89), .B(n685), .Z(G176) );
  NAND2_X1 U770 ( .A1(G160), .A2(G40), .ZN(n716) );
  NOR2_X1 U771 ( .A1(n718), .A2(n716), .ZN(n817) );
  NAND2_X1 U772 ( .A1(G140), .A2(n515), .ZN(n687) );
  NAND2_X1 U773 ( .A1(G104), .A2(n878), .ZN(n686) );
  NAND2_X1 U774 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U775 ( .A(KEYINPUT34), .B(n688), .ZN(n693) );
  NAND2_X1 U776 ( .A1(G128), .A2(n885), .ZN(n690) );
  NAND2_X1 U777 ( .A1(G116), .A2(n882), .ZN(n689) );
  NAND2_X1 U778 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U779 ( .A(n691), .B(KEYINPUT35), .Z(n692) );
  NOR2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U781 ( .A(KEYINPUT36), .B(n694), .Z(n695) );
  XNOR2_X1 U782 ( .A(KEYINPUT91), .B(n695), .ZN(n893) );
  XNOR2_X1 U783 ( .A(G2067), .B(KEYINPUT37), .ZN(n806) );
  NOR2_X1 U784 ( .A1(n893), .A2(n806), .ZN(n963) );
  NAND2_X1 U785 ( .A1(n817), .A2(n963), .ZN(n813) );
  NAND2_X1 U786 ( .A1(G119), .A2(n885), .ZN(n697) );
  NAND2_X1 U787 ( .A1(G131), .A2(n515), .ZN(n696) );
  NAND2_X1 U788 ( .A1(n697), .A2(n696), .ZN(n700) );
  NAND2_X1 U789 ( .A1(n878), .A2(G95), .ZN(n698) );
  XOR2_X1 U790 ( .A(KEYINPUT92), .B(n698), .Z(n699) );
  NOR2_X1 U791 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n882), .A2(G107), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n702), .A2(n701), .ZN(n870) );
  AND2_X1 U794 ( .A1(n870), .A2(G1991), .ZN(n713) );
  XOR2_X1 U795 ( .A(KEYINPUT93), .B(KEYINPUT38), .Z(n704) );
  NAND2_X1 U796 ( .A1(G105), .A2(n878), .ZN(n703) );
  XNOR2_X1 U797 ( .A(n704), .B(n703), .ZN(n711) );
  NAND2_X1 U798 ( .A1(G129), .A2(n885), .ZN(n706) );
  NAND2_X1 U799 ( .A1(G117), .A2(n882), .ZN(n705) );
  NAND2_X1 U800 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n515), .A2(G141), .ZN(n707) );
  XOR2_X1 U802 ( .A(KEYINPUT94), .B(n707), .Z(n708) );
  NOR2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n874) );
  AND2_X1 U805 ( .A1(n874), .A2(G1996), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n962) );
  INV_X1 U807 ( .A(n817), .ZN(n714) );
  NOR2_X1 U808 ( .A1(n962), .A2(n714), .ZN(n809) );
  XNOR2_X1 U809 ( .A(KEYINPUT95), .B(n809), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n813), .A2(n715), .ZN(n803) );
  INV_X1 U811 ( .A(G1341), .ZN(n989) );
  XOR2_X1 U812 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n729) );
  NAND2_X1 U813 ( .A1(n989), .A2(n729), .ZN(n719) );
  INV_X1 U814 ( .A(n716), .ZN(n717) );
  NAND2_X2 U815 ( .A1(n718), .A2(n717), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n719), .A2(n765), .ZN(n722) );
  INV_X1 U817 ( .A(n765), .ZN(n748) );
  AND2_X1 U818 ( .A1(G1996), .A2(n748), .ZN(n720) );
  NAND2_X1 U819 ( .A1(n720), .A2(n729), .ZN(n721) );
  NAND2_X1 U820 ( .A1(n722), .A2(n721), .ZN(n728) );
  NAND2_X1 U821 ( .A1(G1348), .A2(n765), .ZN(n723) );
  XNOR2_X1 U822 ( .A(n723), .B(KEYINPUT98), .ZN(n725) );
  NAND2_X1 U823 ( .A1(n748), .A2(G2067), .ZN(n724) );
  NAND2_X1 U824 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U825 ( .A1(n1001), .A2(n733), .ZN(n727) );
  NOR2_X1 U826 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n729), .ZN(n730) );
  NOR2_X1 U828 ( .A1(n730), .A2(n988), .ZN(n731) );
  NAND2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n740) );
  AND2_X1 U830 ( .A1(n733), .A2(n1001), .ZN(n738) );
  NAND2_X1 U831 ( .A1(n748), .A2(G2072), .ZN(n734) );
  XOR2_X1 U832 ( .A(KEYINPUT27), .B(n734), .Z(n736) );
  NAND2_X1 U833 ( .A1(G1956), .A2(n765), .ZN(n735) );
  NAND2_X1 U834 ( .A1(n736), .A2(n735), .ZN(n743) );
  NOR2_X1 U835 ( .A1(G299), .A2(n743), .ZN(n737) );
  NOR2_X1 U836 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U837 ( .A1(G299), .A2(n743), .ZN(n744) );
  XNOR2_X1 U838 ( .A(KEYINPUT28), .B(n744), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U840 ( .A(n747), .B(KEYINPUT29), .ZN(n752) );
  XOR2_X1 U841 ( .A(KEYINPUT25), .B(G2078), .Z(n934) );
  NOR2_X1 U842 ( .A1(n934), .A2(n765), .ZN(n750) );
  XNOR2_X1 U843 ( .A(G1961), .B(KEYINPUT96), .ZN(n907) );
  NOR2_X1 U844 ( .A1(n748), .A2(n907), .ZN(n749) );
  NOR2_X1 U845 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U846 ( .A1(G301), .A2(n754), .ZN(n751) );
  NOR2_X1 U847 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U848 ( .A(n753), .B(KEYINPUT101), .ZN(n764) );
  AND2_X1 U849 ( .A1(G301), .A2(n754), .ZN(n759) );
  NAND2_X1 U850 ( .A1(G8), .A2(n765), .ZN(n797) );
  NOR2_X1 U851 ( .A1(G1966), .A2(n797), .ZN(n777) );
  NOR2_X1 U852 ( .A1(G2084), .A2(n765), .ZN(n774) );
  NOR2_X1 U853 ( .A1(n777), .A2(n774), .ZN(n755) );
  NAND2_X1 U854 ( .A1(G8), .A2(n755), .ZN(n756) );
  XNOR2_X1 U855 ( .A(KEYINPUT30), .B(n756), .ZN(n757) );
  NOR2_X1 U856 ( .A1(G168), .A2(n757), .ZN(n758) );
  NOR2_X1 U857 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U858 ( .A1(n764), .A2(n763), .ZN(n775) );
  NAND2_X1 U859 ( .A1(n775), .A2(G286), .ZN(n771) );
  NOR2_X1 U860 ( .A1(G1971), .A2(n797), .ZN(n767) );
  NOR2_X1 U861 ( .A1(G2090), .A2(n765), .ZN(n766) );
  NOR2_X1 U862 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U863 ( .A1(n768), .A2(G303), .ZN(n769) );
  XOR2_X1 U864 ( .A(KEYINPUT103), .B(n769), .Z(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U866 ( .A1(n772), .A2(G8), .ZN(n773) );
  XNOR2_X1 U867 ( .A(n773), .B(KEYINPUT32), .ZN(n781) );
  NAND2_X1 U868 ( .A1(G8), .A2(n774), .ZN(n779) );
  INV_X1 U869 ( .A(n775), .ZN(n776) );
  NOR2_X1 U870 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n791) );
  NOR2_X1 U873 ( .A1(G1976), .A2(G288), .ZN(n786) );
  NOR2_X1 U874 ( .A1(G1971), .A2(G303), .ZN(n782) );
  NOR2_X1 U875 ( .A1(n786), .A2(n782), .ZN(n1005) );
  NAND2_X1 U876 ( .A1(n791), .A2(n1005), .ZN(n783) );
  NAND2_X1 U877 ( .A1(G1976), .A2(G288), .ZN(n996) );
  NAND2_X1 U878 ( .A1(n783), .A2(n996), .ZN(n784) );
  NOR2_X1 U879 ( .A1(KEYINPUT33), .A2(n785), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n786), .A2(KEYINPUT33), .ZN(n787) );
  NOR2_X1 U881 ( .A1(n797), .A2(n787), .ZN(n788) );
  XOR2_X1 U882 ( .A(G1981), .B(G305), .Z(n990) );
  AND2_X1 U883 ( .A1(n790), .A2(n990), .ZN(n801) );
  NOR2_X1 U884 ( .A1(G2090), .A2(G303), .ZN(n792) );
  NAND2_X1 U885 ( .A1(G8), .A2(n792), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n791), .A2(n793), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n794), .A2(n797), .ZN(n799) );
  NOR2_X1 U888 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U889 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  OR2_X1 U890 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U891 ( .A1(n799), .A2(n798), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n998) );
  NAND2_X1 U894 ( .A1(n998), .A2(n817), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n805), .A2(n804), .ZN(n820) );
  NAND2_X1 U896 ( .A1(n893), .A2(n806), .ZN(n965) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n874), .ZN(n959) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n870), .ZN(n976) );
  NOR2_X1 U900 ( .A1(n807), .A2(n976), .ZN(n808) );
  NOR2_X1 U901 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U902 ( .A1(n959), .A2(n810), .ZN(n811) );
  XNOR2_X1 U903 ( .A(KEYINPUT104), .B(n811), .ZN(n812) );
  XNOR2_X1 U904 ( .A(n812), .B(KEYINPUT39), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n965), .A2(n815), .ZN(n816) );
  XOR2_X1 U907 ( .A(KEYINPUT105), .B(n816), .Z(n818) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n820), .A2(n819), .ZN(n822) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n821) );
  XNOR2_X1 U911 ( .A(n822), .B(n821), .ZN(G329) );
  NAND2_X1 U912 ( .A1(G2106), .A2(n823), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n824) );
  NAND2_X1 U914 ( .A1(G661), .A2(n824), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U916 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U918 ( .A(G132), .ZN(G219) );
  INV_X1 U919 ( .A(G120), .ZN(G236) );
  INV_X1 U920 ( .A(G96), .ZN(G221) );
  INV_X1 U921 ( .A(G82), .ZN(G220) );
  INV_X1 U922 ( .A(G69), .ZN(G235) );
  NOR2_X1 U923 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  NOR2_X1 U925 ( .A1(n829), .A2(G860), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(n830), .ZN(G145) );
  INV_X1 U927 ( .A(n832), .ZN(G319) );
  XOR2_X1 U928 ( .A(G2096), .B(KEYINPUT108), .Z(n834) );
  XNOR2_X1 U929 ( .A(G2090), .B(KEYINPUT43), .ZN(n833) );
  XNOR2_X1 U930 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U931 ( .A(n835), .B(KEYINPUT42), .Z(n837) );
  XNOR2_X1 U932 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U933 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U934 ( .A(G2678), .B(G2100), .Z(n839) );
  XNOR2_X1 U935 ( .A(G2084), .B(G2078), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U937 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U938 ( .A(KEYINPUT110), .B(G1981), .Z(n843) );
  XNOR2_X1 U939 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n844), .B(KEYINPUT41), .Z(n846) );
  XNOR2_X1 U942 ( .A(G1971), .B(G1976), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(G1956), .B(G1961), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1986), .B(G1966), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U947 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U948 ( .A(KEYINPUT109), .B(G2474), .ZN(n851) );
  XNOR2_X1 U949 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n885), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U952 ( .A1(G112), .A2(n882), .ZN(n854) );
  XOR2_X1 U953 ( .A(KEYINPUT111), .B(n854), .Z(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U955 ( .A1(G136), .A2(n515), .ZN(n858) );
  NAND2_X1 U956 ( .A1(G100), .A2(n878), .ZN(n857) );
  NAND2_X1 U957 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U958 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n872) );
  NAND2_X1 U960 ( .A1(G139), .A2(n515), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G103), .A2(n878), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G127), .A2(n885), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G115), .A2(n882), .ZN(n863) );
  NAND2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(KEYINPUT47), .B(n865), .ZN(n866) );
  XNOR2_X1 U967 ( .A(KEYINPUT113), .B(n866), .ZN(n867) );
  NOR2_X1 U968 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U969 ( .A(KEYINPUT114), .B(n869), .Z(n966) );
  XOR2_X1 U970 ( .A(n870), .B(n966), .Z(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n973), .B(n873), .ZN(n876) );
  XOR2_X1 U973 ( .A(G164), .B(n874), .Z(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n890) );
  NAND2_X1 U975 ( .A1(G142), .A2(n515), .ZN(n880) );
  NAND2_X1 U976 ( .A1(G106), .A2(n878), .ZN(n879) );
  NAND2_X1 U977 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n881), .B(KEYINPUT45), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G118), .A2(n882), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n884), .A2(n883), .ZN(n888) );
  NAND2_X1 U981 ( .A1(n885), .A2(G130), .ZN(n886) );
  XOR2_X1 U982 ( .A(KEYINPUT112), .B(n886), .Z(n887) );
  NOR2_X1 U983 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U984 ( .A(n890), .B(n889), .Z(n892) );
  XNOR2_X1 U985 ( .A(G160), .B(G162), .ZN(n891) );
  XNOR2_X1 U986 ( .A(n892), .B(n891), .ZN(n894) );
  XNOR2_X1 U987 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U988 ( .A1(G37), .A2(n895), .ZN(G395) );
  INV_X1 U989 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U990 ( .A(n988), .B(n896), .ZN(n898) );
  XNOR2_X1 U991 ( .A(G171), .B(n1001), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n899), .B(G286), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G37), .A2(n900), .ZN(G397) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT49), .B(n901), .Z(n902) );
  NAND2_X1 U997 ( .A1(G319), .A2(n902), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G401), .A2(n903), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G395), .A2(G397), .ZN(n904) );
  XOR2_X1 U1000 ( .A(KEYINPUT115), .B(n904), .Z(n905) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(G225) );
  INV_X1 U1002 ( .A(G225), .ZN(G308) );
  INV_X1 U1003 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1004 ( .A(n907), .B(G5), .Z(n921) );
  XNOR2_X1 U1005 ( .A(G1348), .B(KEYINPUT59), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n908), .B(G4), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(G1956), .B(G20), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(G19), .B(G1341), .ZN(n909) );
  NOR2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(n915) );
  XOR2_X1 U1011 ( .A(KEYINPUT125), .B(G1981), .Z(n913) );
  XNOR2_X1 U1012 ( .A(G6), .B(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1014 ( .A(KEYINPUT60), .B(n916), .Z(n918) );
  XNOR2_X1 U1015 ( .A(G1966), .B(G21), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1017 ( .A(KEYINPUT126), .B(n919), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1971), .B(G22), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(G23), .B(G1976), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n925) );
  XOR2_X1 U1022 ( .A(G1986), .B(G24), .Z(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(KEYINPUT58), .B(n926), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n930) );
  XOR2_X1 U1026 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n929) );
  XNOR2_X1 U1027 ( .A(n930), .B(n929), .ZN(n932) );
  INV_X1 U1028 ( .A(G16), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(G11), .ZN(n957) );
  XOR2_X1 U1031 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n953) );
  XNOR2_X1 U1032 ( .A(G2090), .B(G35), .ZN(n948) );
  XNOR2_X1 U1033 ( .A(G1996), .B(G32), .ZN(n936) );
  XNOR2_X1 U1034 ( .A(n934), .B(G27), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(KEYINPUT120), .B(n937), .ZN(n943) );
  XOR2_X1 U1037 ( .A(G2072), .B(G33), .Z(n938) );
  NAND2_X1 U1038 ( .A1(n938), .A2(G28), .ZN(n941) );
  XOR2_X1 U1039 ( .A(G25), .B(G1991), .Z(n939) );
  XNOR2_X1 U1040 ( .A(KEYINPUT119), .B(n939), .ZN(n940) );
  NOR2_X1 U1041 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n945) );
  XNOR2_X1 U1043 ( .A(G26), .B(G2067), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1045 ( .A(KEYINPUT53), .B(n946), .ZN(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1047 ( .A(G2084), .B(G34), .Z(n949) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(n949), .ZN(n950) );
  NAND2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1050 ( .A(n953), .B(n952), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n954), .A2(G29), .ZN(n955) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n955), .ZN(n956) );
  NOR2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n987) );
  XOR2_X1 U1054 ( .A(G2090), .B(G162), .Z(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1056 ( .A(KEYINPUT51), .B(n960), .Z(n961) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n981) );
  INV_X1 U1058 ( .A(n963), .ZN(n964) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n972) );
  XOR2_X1 U1060 ( .A(G2072), .B(n966), .Z(n968) );
  XNOR2_X1 U1061 ( .A(G164), .B(G2078), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(KEYINPUT50), .B(n969), .Z(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT117), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n979) );
  XNOR2_X1 U1066 ( .A(G160), .B(G2084), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(KEYINPUT116), .ZN(n978) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1072 ( .A(KEYINPUT52), .B(n982), .Z(n983) );
  NOR2_X1 U1073 ( .A1(KEYINPUT55), .A2(n983), .ZN(n984) );
  XOR2_X1 U1074 ( .A(KEYINPUT118), .B(n984), .Z(n985) );
  NAND2_X1 U1075 ( .A1(G29), .A2(n985), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n1015) );
  XOR2_X1 U1077 ( .A(G16), .B(KEYINPUT56), .Z(n1013) );
  XNOR2_X1 U1078 ( .A(n989), .B(n988), .ZN(n994) );
  XNOR2_X1 U1079 ( .A(G1966), .B(G168), .ZN(n991) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(n992), .B(KEYINPUT57), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1010) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n995) );
  NAND2_X1 U1084 ( .A1(n996), .A2(n995), .ZN(n1007) );
  XNOR2_X1 U1085 ( .A(G171), .B(G1961), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(G1956), .B(G299), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XOR2_X1 U1089 ( .A(n1001), .B(G1348), .Z(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(n1008), .B(KEYINPUT123), .ZN(n1009) );
  NOR2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT124), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1096 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1097 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1098 ( .A(n1016), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

