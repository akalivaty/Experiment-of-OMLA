

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595;

  XNOR2_X1 U320 ( .A(n457), .B(n456), .ZN(n489) );
  OR2_X1 U321 ( .A1(n476), .A2(n475), .ZN(n500) );
  XNOR2_X1 U322 ( .A(n390), .B(KEYINPUT48), .ZN(n559) );
  XOR2_X1 U323 ( .A(n311), .B(n310), .Z(n538) );
  XOR2_X1 U324 ( .A(n396), .B(n418), .Z(n288) );
  XNOR2_X1 U325 ( .A(n346), .B(KEYINPUT111), .ZN(n347) );
  XNOR2_X1 U326 ( .A(n348), .B(n347), .ZN(n382) );
  XNOR2_X1 U327 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U328 ( .A(n338), .B(n337), .ZN(n343) );
  XNOR2_X1 U329 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n456) );
  XNOR2_X1 U330 ( .A(n445), .B(KEYINPUT55), .ZN(n446) );
  XNOR2_X1 U331 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U332 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U333 ( .A(n380), .B(n379), .ZN(n592) );
  XNOR2_X1 U334 ( .A(KEYINPUT122), .B(G183GAT), .ZN(n449) );
  XNOR2_X1 U335 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U336 ( .A(n450), .B(n449), .ZN(G1350GAT) );
  XNOR2_X1 U337 ( .A(n486), .B(n485), .ZN(G1330GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n290) );
  XNOR2_X1 U339 ( .A(G15GAT), .B(G71GAT), .ZN(n289) );
  XNOR2_X1 U340 ( .A(n290), .B(n289), .ZN(n311) );
  INV_X1 U341 ( .A(KEYINPUT17), .ZN(n291) );
  NAND2_X1 U342 ( .A1(KEYINPUT19), .A2(n291), .ZN(n294) );
  INV_X1 U343 ( .A(KEYINPUT19), .ZN(n292) );
  NAND2_X1 U344 ( .A1(n292), .A2(KEYINPUT17), .ZN(n293) );
  NAND2_X1 U345 ( .A1(n294), .A2(n293), .ZN(n296) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n396) );
  XOR2_X1 U348 ( .A(G113GAT), .B(KEYINPUT0), .Z(n418) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U350 ( .A(n288), .B(n297), .ZN(n309) );
  XOR2_X1 U351 ( .A(G99GAT), .B(G134GAT), .Z(n299) );
  XNOR2_X1 U352 ( .A(G43GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U354 ( .A(G183GAT), .B(G176GAT), .Z(n301) );
  XNOR2_X1 U355 ( .A(G127GAT), .B(G120GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U357 ( .A(n303), .B(n302), .Z(n307) );
  XOR2_X1 U358 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n305) );
  XNOR2_X1 U359 ( .A(KEYINPUT20), .B(KEYINPUT65), .ZN(n304) );
  XNOR2_X1 U360 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U361 ( .A(G113GAT), .B(G50GAT), .Z(n313) );
  XNOR2_X1 U362 ( .A(G36GAT), .B(G29GAT), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U364 ( .A(G8GAT), .B(G141GAT), .Z(n315) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G1GAT), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(n317), .B(n316), .Z(n322) );
  XOR2_X1 U368 ( .A(KEYINPUT68), .B(KEYINPUT70), .Z(n319) );
  NAND2_X1 U369 ( .A1(G229GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U370 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U371 ( .A(KEYINPUT69), .B(n320), .ZN(n321) );
  XNOR2_X1 U372 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U373 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n324) );
  XNOR2_X1 U374 ( .A(G197GAT), .B(KEYINPUT29), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U376 ( .A(n326), .B(n325), .Z(n330) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n327), .B(KEYINPUT8), .ZN(n361) );
  XNOR2_X1 U379 ( .A(G15GAT), .B(KEYINPUT71), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n328), .B(G22GAT), .ZN(n378) );
  XNOR2_X1 U381 ( .A(n361), .B(n378), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n584) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(G57GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n331), .B(G148GAT), .ZN(n410) );
  XNOR2_X1 U385 ( .A(G176GAT), .B(G64GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n332), .B(KEYINPUT74), .ZN(n392) );
  XNOR2_X1 U387 ( .A(n410), .B(n392), .ZN(n345) );
  XOR2_X1 U388 ( .A(G71GAT), .B(KEYINPUT13), .Z(n366) );
  XOR2_X1 U389 ( .A(G204GAT), .B(G78GAT), .Z(n436) );
  XOR2_X1 U390 ( .A(n366), .B(n436), .Z(n338) );
  XOR2_X1 U391 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n334) );
  XNOR2_X1 U392 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n336) );
  NAND2_X1 U394 ( .A1(G230GAT), .A2(G233GAT), .ZN(n335) );
  XOR2_X1 U395 ( .A(G99GAT), .B(G106GAT), .Z(n353) );
  XOR2_X1 U396 ( .A(KEYINPUT73), .B(KEYINPUT75), .Z(n340) );
  XNOR2_X1 U397 ( .A(G85GAT), .B(G92GAT), .ZN(n339) );
  XNOR2_X1 U398 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U399 ( .A(n353), .B(n341), .Z(n342) );
  XNOR2_X1 U400 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n481) );
  XOR2_X1 U402 ( .A(KEYINPUT41), .B(n481), .Z(n567) );
  INV_X1 U403 ( .A(n567), .ZN(n451) );
  NAND2_X1 U404 ( .A1(n584), .A2(n451), .ZN(n348) );
  INV_X1 U405 ( .A(KEYINPUT46), .ZN(n346) );
  XNOR2_X1 U406 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n350) );
  AND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U408 ( .A(n350), .B(n349), .ZN(n352) );
  INV_X1 U409 ( .A(KEYINPUT10), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n355) );
  XOR2_X1 U411 ( .A(G50GAT), .B(G162GAT), .Z(n440) );
  XNOR2_X1 U412 ( .A(n353), .B(n440), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U414 ( .A(G218GAT), .B(G92GAT), .Z(n357) );
  XNOR2_X1 U415 ( .A(G190GAT), .B(KEYINPUT76), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U417 ( .A(G36GAT), .B(n358), .Z(n405) );
  XOR2_X1 U418 ( .A(n359), .B(n405), .Z(n363) );
  XNOR2_X1 U419 ( .A(G29GAT), .B(G134GAT), .ZN(n360) );
  XNOR2_X1 U420 ( .A(n360), .B(G85GAT), .ZN(n411) );
  XNOR2_X1 U421 ( .A(n361), .B(n411), .ZN(n362) );
  XNOR2_X1 U422 ( .A(n363), .B(n362), .ZN(n575) );
  XOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT79), .Z(n365) );
  XNOR2_X1 U424 ( .A(KEYINPUT14), .B(KEYINPUT80), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n365), .B(n364), .ZN(n370) );
  XOR2_X1 U426 ( .A(G1GAT), .B(G127GAT), .Z(n419) );
  XOR2_X1 U427 ( .A(n366), .B(n419), .Z(n368) );
  XNOR2_X1 U428 ( .A(G155GAT), .B(G57GAT), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U430 ( .A(n370), .B(n369), .Z(n372) );
  NAND2_X1 U431 ( .A1(G231GAT), .A2(G233GAT), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n376) );
  XOR2_X1 U433 ( .A(KEYINPUT12), .B(G78GAT), .Z(n374) );
  XNOR2_X1 U434 ( .A(G211GAT), .B(G64GAT), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U436 ( .A(n376), .B(n375), .Z(n380) );
  XNOR2_X1 U437 ( .A(G8GAT), .B(G183GAT), .ZN(n377) );
  XNOR2_X1 U438 ( .A(n377), .B(KEYINPUT78), .ZN(n391) );
  XNOR2_X1 U439 ( .A(n378), .B(n391), .ZN(n379) );
  INV_X1 U440 ( .A(n592), .ZN(n572) );
  AND2_X1 U441 ( .A1(n575), .A2(n572), .ZN(n381) );
  AND2_X1 U442 ( .A1(n382), .A2(n381), .ZN(n383) );
  XOR2_X1 U443 ( .A(KEYINPUT47), .B(n383), .Z(n389) );
  XNOR2_X1 U444 ( .A(n575), .B(KEYINPUT77), .ZN(n578) );
  XOR2_X1 U445 ( .A(KEYINPUT36), .B(n578), .Z(n493) );
  NOR2_X1 U446 ( .A1(n572), .A2(n493), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n384), .B(KEYINPUT45), .ZN(n385) );
  NAND2_X1 U448 ( .A1(n385), .A2(n481), .ZN(n386) );
  NOR2_X1 U449 ( .A1(n584), .A2(n386), .ZN(n387) );
  XNOR2_X1 U450 ( .A(KEYINPUT112), .B(n387), .ZN(n388) );
  NOR2_X1 U451 ( .A1(n389), .A2(n388), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n403) );
  XOR2_X1 U453 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n394) );
  XNOR2_X1 U454 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U456 ( .A(G197GAT), .B(n395), .Z(n428) );
  XOR2_X1 U457 ( .A(KEYINPUT95), .B(G204GAT), .Z(n398) );
  XNOR2_X1 U458 ( .A(n396), .B(KEYINPUT94), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U460 ( .A(n428), .B(n399), .Z(n401) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U463 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n536) );
  NOR2_X1 U465 ( .A1(n559), .A2(n536), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n406), .B(KEYINPUT54), .ZN(n426) );
  XOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n408) );
  NAND2_X1 U468 ( .A1(G225GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U470 ( .A(n409), .B(KEYINPUT6), .Z(n413) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n415) );
  XNOR2_X1 U474 ( .A(G162GAT), .B(KEYINPUT92), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U479 ( .A(KEYINPUT2), .B(KEYINPUT90), .Z(n423) );
  XNOR2_X1 U480 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(G141GAT), .B(n424), .Z(n429) );
  XOR2_X1 U483 ( .A(n425), .B(n429), .Z(n473) );
  XNOR2_X1 U484 ( .A(KEYINPUT93), .B(n473), .ZN(n560) );
  NAND2_X1 U485 ( .A1(n426), .A2(n560), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n427), .B(KEYINPUT64), .ZN(n490) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n444) );
  XOR2_X1 U488 ( .A(G106GAT), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U489 ( .A(G22GAT), .B(G148GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U491 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n433) );
  XNOR2_X1 U492 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U494 ( .A(n435), .B(n434), .Z(n442) );
  XOR2_X1 U495 ( .A(n436), .B(KEYINPUT24), .Z(n438) );
  NAND2_X1 U496 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n464) );
  NOR2_X1 U501 ( .A1(n490), .A2(n464), .ZN(n447) );
  INV_X1 U502 ( .A(KEYINPUT119), .ZN(n445) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U504 ( .A1(n538), .A2(n448), .ZN(n577) );
  NAND2_X1 U505 ( .A1(n577), .A2(n592), .ZN(n450) );
  NAND2_X1 U506 ( .A1(n577), .A2(n451), .ZN(n455) );
  XOR2_X1 U507 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n453) );
  XOR2_X1 U508 ( .A(G176GAT), .B(KEYINPUT56), .Z(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U510 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XNOR2_X1 U511 ( .A(KEYINPUT27), .B(n536), .ZN(n466) );
  NAND2_X1 U512 ( .A1(n464), .A2(n538), .ZN(n457) );
  NOR2_X1 U513 ( .A1(n466), .A2(n489), .ZN(n562) );
  INV_X1 U514 ( .A(KEYINPUT97), .ZN(n458) );
  NAND2_X1 U515 ( .A1(n562), .A2(n458), .ZN(n461) );
  INV_X1 U516 ( .A(n562), .ZN(n459) );
  NAND2_X1 U517 ( .A1(n459), .A2(KEYINPUT97), .ZN(n460) );
  NAND2_X1 U518 ( .A1(n461), .A2(n460), .ZN(n471) );
  NOR2_X1 U519 ( .A1(n538), .A2(n536), .ZN(n462) );
  NOR2_X1 U520 ( .A1(n464), .A2(n462), .ZN(n463) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n463), .Z(n469) );
  XNOR2_X1 U522 ( .A(n464), .B(KEYINPUT66), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(KEYINPUT28), .ZN(n508) );
  NOR2_X1 U524 ( .A1(n508), .A2(n560), .ZN(n468) );
  INV_X1 U525 ( .A(n466), .ZN(n467) );
  NAND2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n545) );
  INV_X1 U527 ( .A(n538), .ZN(n547) );
  NOR2_X1 U528 ( .A1(n545), .A2(n547), .ZN(n472) );
  OR2_X1 U529 ( .A1(n469), .A2(n472), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n471), .A2(n470), .ZN(n476) );
  INV_X1 U531 ( .A(n472), .ZN(n474) );
  AND2_X1 U532 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n592), .A2(n500), .ZN(n478) );
  INV_X1 U534 ( .A(KEYINPUT102), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n493), .A2(n479), .ZN(n480) );
  XOR2_X1 U537 ( .A(KEYINPUT37), .B(n480), .Z(n534) );
  INV_X1 U538 ( .A(n584), .ZN(n563) );
  INV_X1 U539 ( .A(n481), .ZN(n589) );
  NOR2_X1 U540 ( .A1(n563), .A2(n589), .ZN(n501) );
  AND2_X1 U541 ( .A1(n534), .A2(n501), .ZN(n482) );
  XOR2_X2 U542 ( .A(KEYINPUT38), .B(n482), .Z(n520) );
  NOR2_X1 U543 ( .A1(n538), .A2(n520), .ZN(n486) );
  XNOR2_X1 U544 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n484) );
  INV_X1 U545 ( .A(G43GAT), .ZN(n483) );
  NAND2_X1 U546 ( .A1(n577), .A2(n584), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT120), .B(G169GAT), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1348GAT) );
  INV_X1 U549 ( .A(KEYINPUT125), .ZN(n492) );
  OR2_X1 U550 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n492), .B(n491), .ZN(n583) );
  NOR2_X1 U552 ( .A1(n493), .A2(n583), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT62), .B(n494), .ZN(n496) );
  INV_X1 U554 ( .A(G218GAT), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n496), .B(n495), .ZN(G1355GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT16), .B(KEYINPUT81), .Z(n498) );
  OR2_X1 U557 ( .A1(n578), .A2(n572), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(n499) );
  NOR2_X1 U559 ( .A1(n500), .A2(n499), .ZN(n523) );
  NAND2_X1 U560 ( .A1(n501), .A2(n523), .ZN(n509) );
  NOR2_X1 U561 ( .A1(n560), .A2(n509), .ZN(n503) );
  XNOR2_X1 U562 ( .A(KEYINPUT34), .B(KEYINPUT98), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U564 ( .A(G1GAT), .B(n504), .Z(G1324GAT) );
  NOR2_X1 U565 ( .A1(n536), .A2(n509), .ZN(n505) );
  XOR2_X1 U566 ( .A(G8GAT), .B(n505), .Z(G1325GAT) );
  NOR2_X1 U567 ( .A1(n538), .A2(n509), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n506) );
  XNOR2_X1 U569 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  INV_X1 U570 ( .A(n508), .ZN(n542) );
  NOR2_X1 U571 ( .A1(n542), .A2(n509), .ZN(n511) );
  XNOR2_X1 U572 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(n512), .ZN(G1327GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n514) );
  XNOR2_X1 U576 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(n516) );
  NOR2_X1 U578 ( .A1(n520), .A2(n560), .ZN(n515) );
  XOR2_X1 U579 ( .A(n516), .B(n515), .Z(G1328GAT) );
  NOR2_X1 U580 ( .A1(n520), .A2(n536), .ZN(n518) );
  XNOR2_X1 U581 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U583 ( .A(G36GAT), .B(n519), .ZN(G1329GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n542), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(G1331GAT) );
  NOR2_X1 U587 ( .A1(n584), .A2(n567), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n533), .A2(n523), .ZN(n530) );
  NOR2_X1 U589 ( .A1(n560), .A2(n530), .ZN(n524) );
  XOR2_X1 U590 ( .A(n524), .B(KEYINPUT42), .Z(n525) );
  XNOR2_X1 U591 ( .A(G57GAT), .B(n525), .ZN(G1332GAT) );
  NOR2_X1 U592 ( .A1(n536), .A2(n530), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT108), .B(n526), .Z(n527) );
  XNOR2_X1 U594 ( .A(G64GAT), .B(n527), .ZN(G1333GAT) );
  NOR2_X1 U595 ( .A1(n538), .A2(n530), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(G1334GAT) );
  NOR2_X1 U598 ( .A1(n542), .A2(n530), .ZN(n532) );
  XNOR2_X1 U599 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n531) );
  XNOR2_X1 U600 ( .A(n532), .B(n531), .ZN(G1335GAT) );
  NAND2_X1 U601 ( .A1(n534), .A2(n533), .ZN(n541) );
  NOR2_X1 U602 ( .A1(n560), .A2(n541), .ZN(n535) );
  XOR2_X1 U603 ( .A(G85GAT), .B(n535), .Z(G1336GAT) );
  NOR2_X1 U604 ( .A1(n536), .A2(n541), .ZN(n537) );
  XOR2_X1 U605 ( .A(G92GAT), .B(n537), .Z(G1337GAT) );
  NOR2_X1 U606 ( .A1(n538), .A2(n541), .ZN(n539) );
  XOR2_X1 U607 ( .A(KEYINPUT110), .B(n539), .Z(n540) );
  XNOR2_X1 U608 ( .A(G99GAT), .B(n540), .ZN(G1338GAT) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U610 ( .A(KEYINPUT44), .B(n543), .Z(n544) );
  XNOR2_X1 U611 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  NOR2_X1 U612 ( .A1(n559), .A2(n545), .ZN(n546) );
  NAND2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n548), .B(KEYINPUT113), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n556), .A2(n584), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n551) );
  NAND2_X1 U618 ( .A1(n556), .A2(n451), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G120GAT), .B(n552), .ZN(G1341GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n554) );
  NAND2_X1 U622 ( .A1(n556), .A2(n592), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U624 ( .A(G127GAT), .B(n555), .ZN(G1342GAT) );
  XOR2_X1 U625 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U626 ( .A1(n556), .A2(n578), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  NOR2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n574) );
  NOR2_X1 U630 ( .A1(n563), .A2(n574), .ZN(n564) );
  XOR2_X1 U631 ( .A(G141GAT), .B(n564), .Z(G1344GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n566) );
  XNOR2_X1 U633 ( .A(KEYINPUT116), .B(KEYINPUT53), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n571) );
  NOR2_X1 U635 ( .A1(n567), .A2(n574), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1345GAT) );
  NOR2_X1 U639 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U640 ( .A(G155GAT), .B(n573), .Z(G1346GAT) );
  NOR2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(G162GAT), .B(n576), .Z(G1347GAT) );
  AND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n582) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n579), .B(KEYINPUT123), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT124), .B(n580), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1351GAT) );
  INV_X1 U648 ( .A(n583), .ZN(n593) );
  NAND2_X1 U649 ( .A1(n593), .A2(n584), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT126), .B(KEYINPUT59), .Z(n586) );
  XNOR2_X1 U651 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1352GAT) );
  XOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT61), .Z(n591) );
  NAND2_X1 U655 ( .A1(n593), .A2(n589), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n591), .B(n590), .ZN(G1353GAT) );
  XOR2_X1 U657 ( .A(G211GAT), .B(KEYINPUT127), .Z(n595) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(G1354GAT) );
endmodule

