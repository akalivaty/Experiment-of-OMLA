//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n828,
    new_n829, new_n831, new_n832, new_n833, new_n834, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G15gat), .B(G22gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT92), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G8gat), .ZN(new_n210));
  INV_X1    g009(.A(G8gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n208), .A2(KEYINPUT92), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n213), .B1(G1gat), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(G1gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n217), .A2(new_n210), .A3(new_n212), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT89), .ZN(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G29gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G43gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT15), .B1(new_n228), .B2(G50gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(G50gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n220), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g032(.A1(new_n225), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT14), .B(G29gat), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(new_n221), .ZN(new_n236));
  INV_X1    g035(.A(G50gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G43gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n229), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(KEYINPUT89), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT90), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n228), .B2(G50gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n237), .A2(KEYINPUT90), .A3(G43gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n231), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n224), .A2(new_n226), .B1(new_n230), .B2(new_n231), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n233), .A2(new_n240), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n219), .B(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G229gat), .A2(G233gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT13), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n219), .A2(new_n248), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT91), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(new_n248), .B2(KEYINPUT17), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n247), .A2(new_n246), .ZN(new_n256));
  AOI21_X1  g055(.A(KEYINPUT89), .B1(new_n236), .B2(new_n239), .ZN(new_n257));
  AND4_X1   g056(.A1(KEYINPUT89), .A2(new_n239), .A3(new_n224), .A4(new_n226), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT17), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(KEYINPUT91), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n248), .A2(KEYINPUT17), .B1(new_n216), .B2(new_n218), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n253), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT93), .B1(new_n264), .B2(new_n250), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT18), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n252), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n250), .ZN(new_n268));
  AOI211_X1 g067(.A(new_n268), .B(new_n253), .C1(new_n262), .C2(new_n263), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n269), .A2(KEYINPUT93), .A3(KEYINPUT18), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n207), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n265), .A2(new_n266), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT18), .B1(new_n269), .B2(KEYINPUT93), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n272), .A2(new_n273), .A3(new_n206), .A4(new_n252), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  XOR2_X1   g075(.A(G1gat), .B(G29gat), .Z(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT84), .ZN(new_n278));
  XOR2_X1   g077(.A(G57gat), .B(G85gat), .Z(new_n279));
  XNOR2_X1  g078(.A(new_n278), .B(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n283));
  XNOR2_X1  g082(.A(G141gat), .B(G148gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT2), .ZN(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G162gat), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G141gat), .B(G148gat), .Z(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT79), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT79), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT2), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT80), .B(G155gat), .Z(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT81), .B(G162gat), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n287), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT1), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n297), .B(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n283), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n287), .B(new_n307), .C1(new_n292), .C2(new_n296), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  OR3_X1    g109(.A1(new_n297), .A2(new_n310), .A3(new_n301), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT82), .B(KEYINPUT4), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n312), .B1(new_n297), .B2(new_n301), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n309), .A2(new_n311), .A3(new_n303), .A4(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n305), .A2(new_n314), .ZN(new_n315));
  OR3_X1    g114(.A1(new_n297), .A2(new_n301), .A3(new_n312), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n310), .B1(new_n297), .B2(new_n301), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n316), .A2(new_n283), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n309), .A2(new_n303), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n282), .B1(new_n315), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n314), .A2(new_n305), .B1(new_n318), .B2(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n282), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NOR4_X1   g125(.A1(new_n323), .A2(KEYINPUT85), .A3(new_n325), .A4(new_n282), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT85), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(new_n321), .B2(KEYINPUT6), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT35), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n333));
  XOR2_X1   g132(.A(KEYINPUT73), .B(G211gat), .Z(new_n334));
  INV_X1    g133(.A(G218gat), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n333), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G197gat), .B(G204gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n338), .A3(new_n337), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n338), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n336), .A2(new_n339), .A3(new_n343), .A4(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n307), .B1(new_n345), .B2(KEYINPUT29), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n297), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT29), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n308), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G228gat), .A2(G233gat), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n349), .A2(new_n345), .B1(KEYINPUT86), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n350), .A2(KEYINPUT86), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n353), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n347), .A2(new_n355), .A3(new_n351), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(G22gat), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT31), .B(G50gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G22gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n356), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n355), .B1(new_n347), .B2(new_n351), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n359), .A2(new_n362), .B1(new_n366), .B2(new_n357), .ZN(new_n367));
  AND4_X1   g166(.A1(KEYINPUT87), .A2(new_n366), .A3(new_n357), .A4(new_n362), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n332), .A2(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT27), .B(G183gat), .ZN(new_n371));
  INV_X1    g170(.A(G190gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G183gat), .A2(G190gat), .ZN(new_n376));
  AND2_X1   g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  OR3_X1    g177(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT26), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(KEYINPUT26), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n375), .A2(new_n376), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT25), .ZN(new_n382));
  INV_X1    g181(.A(new_n378), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT23), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n377), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT64), .B(G169gat), .ZN(new_n386));
  INV_X1    g185(.A(G176gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT23), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n390), .B1(G183gat), .B2(G190gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n376), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n382), .B1(new_n389), .B2(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n395));
  NOR2_X1   g194(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n376), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT66), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT66), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(new_n376), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n391), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n385), .B(KEYINPUT25), .C1(G169gat), .C2(new_n388), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n394), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n381), .A2(new_n403), .A3(KEYINPUT75), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(G226gat), .ZN(new_n406));
  INV_X1    g205(.A(G233gat), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT75), .B1(new_n381), .B2(new_n403), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n405), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n381), .A2(new_n403), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n408), .A2(KEYINPUT29), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n411), .A2(new_n345), .A3(new_n414), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n412), .A2(new_n406), .A3(new_n407), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n413), .B1(new_n404), .B2(new_n409), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n345), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G8gat), .B(G36gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(G64gat), .B(G92gat), .ZN(new_n421));
  XOR2_X1   g220(.A(new_n420), .B(new_n421), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n415), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT77), .A3(KEYINPUT30), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT76), .B1(new_n415), .B2(new_n419), .ZN(new_n426));
  INV_X1    g225(.A(new_n345), .ZN(new_n427));
  INV_X1    g226(.A(new_n418), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n416), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT76), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n345), .A3(new_n414), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n426), .A2(new_n432), .A3(new_n423), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT77), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n429), .A2(new_n431), .A3(new_n422), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n436), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n425), .A2(new_n433), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n412), .A2(new_n301), .ZN(new_n441));
  INV_X1    g240(.A(new_n301), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n381), .A2(new_n403), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT67), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT67), .ZN(new_n448));
  AOI211_X1 g247(.A(new_n448), .B(new_n445), .C1(new_n441), .C2(new_n443), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT32), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT33), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n451), .B1(new_n447), .B2(new_n449), .ZN(new_n452));
  XOR2_X1   g251(.A(G15gat), .B(G43gat), .Z(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT68), .ZN(new_n454));
  XOR2_X1   g253(.A(G71gat), .B(G99gat), .Z(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT69), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n451), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n459), .B1(new_n458), .B2(new_n456), .ZN(new_n460));
  OAI211_X1 g259(.A(KEYINPUT32), .B(new_n460), .C1(new_n447), .C2(new_n449), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n444), .A2(new_n446), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n463), .B1(KEYINPUT70), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n444), .B2(new_n446), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n457), .A2(new_n470), .A3(new_n461), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n469), .B1(KEYINPUT71), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(KEYINPUT71), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n457), .B2(new_n461), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n370), .B(new_n440), .C1(new_n472), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT88), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n473), .B(new_n474), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n440), .A4(new_n370), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n425), .A2(new_n433), .A3(new_n437), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n425), .A2(new_n433), .A3(new_n437), .A4(KEYINPUT78), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n483), .A2(new_n330), .A3(new_n484), .A4(new_n438), .ZN(new_n485));
  INV_X1    g284(.A(new_n369), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n469), .A3(new_n471), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT35), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n477), .A2(new_n480), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT36), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n478), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n369), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n309), .A2(new_n316), .A3(new_n317), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n304), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n494), .B(KEYINPUT39), .C1(new_n304), .C2(new_n302), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n282), .C1(KEYINPUT39), .C2(new_n494), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g297(.A1(new_n496), .A2(new_n497), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n439), .A2(new_n322), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  OR3_X1    g299(.A1(new_n415), .A2(new_n419), .A3(KEYINPUT37), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n501), .A2(KEYINPUT38), .A3(new_n423), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n426), .A2(new_n432), .A3(KEYINPUT37), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n345), .B1(new_n428), .B2(new_n416), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n411), .A2(new_n427), .A3(new_n414), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT37), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n501), .A2(new_n506), .A3(new_n423), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT38), .ZN(new_n508));
  AOI22_X1  g307(.A1(new_n502), .A2(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n330), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(new_n435), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n500), .B(new_n486), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n469), .A2(new_n471), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT36), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n491), .A2(new_n492), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n276), .B1(new_n489), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(G99gat), .B(G106gat), .Z(new_n519));
  AND2_X1   g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT98), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n520), .A2(KEYINPUT97), .A3(new_n521), .A4(KEYINPUT7), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n521), .A2(G85gat), .A3(G92gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT97), .B1(G85gat), .B2(G92gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n522), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT99), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT99), .B1(G99gat), .B2(G106gat), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n519), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n534), .A2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(new_n531), .B2(new_n530), .ZN(new_n538));
  INV_X1    g337(.A(new_n519), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n523), .A2(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n522), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n543), .B1(KEYINPUT17), .B2(new_n248), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n262), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n543), .A2(new_n259), .B1(KEYINPUT41), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n518), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n545), .A2(new_n518), .A3(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n546), .A2(KEYINPUT41), .ZN(new_n552));
  INV_X1    g351(.A(G134gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G162gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n548), .B2(KEYINPUT100), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(KEYINPUT100), .A3(new_n550), .A4(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G57gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G64gat), .ZN(new_n561));
  INV_X1    g360(.A(G64gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(G57gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G71gat), .B(G78gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT94), .B1(G71gat), .B2(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR3_X1   g371(.A1(KEYINPUT94), .A2(G71gat), .A3(G78gat), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n566), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n561), .A2(new_n563), .B1(new_n567), .B2(new_n566), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n574), .A2(new_n575), .A3(KEYINPUT95), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n578));
  INV_X1    g377(.A(G71gat), .ZN(new_n579));
  INV_X1    g378(.A(G78gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n581), .A2(new_n571), .B1(G71gat), .B2(G78gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n562), .A2(G57gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n560), .A2(G64gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n568), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n577), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n570), .B1(new_n576), .B2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT95), .B1(new_n574), .B2(new_n575), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n585), .A3(new_n577), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n569), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT96), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G127gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n598), .B1(new_n597), .B2(new_n599), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n594), .A2(KEYINPUT21), .B1(new_n218), .B2(new_n216), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n600), .B2(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n609), .B1(new_n603), .B2(new_n604), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n559), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(G230gat), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(new_n407), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT101), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n620), .B1(new_n587), .B2(new_n542), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n592), .A2(KEYINPUT101), .A3(new_n541), .A4(new_n536), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n589), .A2(new_n593), .A3(new_n542), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT102), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n623), .A2(new_n625), .A3(new_n628), .A4(new_n624), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n542), .A2(new_n624), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n594), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n619), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n590), .A2(new_n591), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT96), .B1(new_n634), .B2(new_n570), .ZN(new_n635));
  AOI211_X1 g434(.A(new_n588), .B(new_n569), .C1(new_n590), .C2(new_n591), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n637), .A2(new_n542), .B1(new_n621), .B2(new_n622), .ZN(new_n638));
  INV_X1    g437(.A(new_n619), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n617), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n627), .A2(new_n629), .B1(new_n594), .B2(new_n631), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n642), .B(new_n616), .C1(new_n643), .C2(new_n619), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n613), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n516), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n647), .A2(new_n330), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT103), .B(G1gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(G1324gat));
  NOR2_X1   g449(.A1(new_n647), .A2(new_n440), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n211), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT104), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G8gat), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n647), .A2(new_n440), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT42), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n656), .B1(KEYINPUT42), .B2(new_n655), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n491), .A2(new_n514), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(G15gat), .B1(new_n647), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n478), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n661), .A2(G15gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n660), .B1(new_n647), .B2(new_n662), .ZN(G1326gat));
  OR3_X1    g462(.A1(new_n647), .A2(KEYINPUT105), .A3(new_n486), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT105), .B1(new_n647), .B2(new_n486), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT43), .B(G22gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1327gat));
  INV_X1    g467(.A(new_n559), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n611), .A2(new_n612), .ZN(new_n670));
  INV_X1    g469(.A(new_n645), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n516), .A2(new_n669), .A3(new_n670), .A4(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n225), .A3(new_n510), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n489), .A2(new_n515), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n669), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n676), .A2(KEYINPUT44), .A3(new_n669), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n670), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n682), .A2(new_n276), .A3(new_n645), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(G29gat), .B1(new_n684), .B2(new_n330), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n675), .A2(new_n685), .ZN(G1328gat));
  NOR3_X1   g485(.A1(new_n672), .A2(G36gat), .A3(new_n440), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT46), .ZN(new_n688));
  OAI21_X1  g487(.A(G36gat), .B1(new_n684), .B2(new_n440), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(G1329gat));
  NAND4_X1  g489(.A1(new_n679), .A2(new_n658), .A3(new_n680), .A4(new_n683), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(G43gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n673), .A2(new_n228), .A3(new_n478), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1330gat));
  OR2_X1    g495(.A1(new_n672), .A2(KEYINPUT106), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n486), .B1(new_n672), .B2(KEYINPUT106), .ZN(new_n698));
  AOI21_X1  g497(.A(G50gat), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT48), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n486), .A2(new_n237), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n681), .A2(new_n683), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n703), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT48), .B1(new_n705), .B2(new_n699), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(new_n706), .ZN(G1331gat));
  NOR3_X1   g506(.A1(new_n613), .A2(new_n275), .A3(new_n671), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n676), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n330), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(new_n560), .ZN(G1332gat));
  INV_X1    g510(.A(new_n709), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n440), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT107), .Z(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(new_n716), .Z(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n709), .B2(new_n659), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n478), .A2(new_n579), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n709), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1334gat));
  NOR2_X1   g521(.A1(new_n709), .A2(new_n486), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n580), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n670), .A2(new_n276), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(new_n671), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n679), .A2(new_n510), .A3(new_n680), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G85gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n725), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT109), .B(KEYINPUT51), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n676), .A2(new_n669), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  AOI211_X1 g530(.A(new_n559), .B(new_n725), .C1(new_n489), .C2(new_n515), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT51), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n731), .B(new_n645), .C1(new_n732), .C2(new_n734), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n330), .A2(G85gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n728), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT110), .ZN(G1336gat));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  INV_X1    g538(.A(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(G92gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n740), .A2(new_n741), .A3(new_n439), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n679), .A2(new_n439), .A3(new_n680), .A4(new_n726), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(KEYINPUT111), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n739), .B(new_n742), .C1(new_n745), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(G92gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n742), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT52), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(G1337gat));
  AOI21_X1  g550(.A(G99gat), .B1(new_n740), .B2(new_n478), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n681), .A2(new_n726), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n658), .A2(G99gat), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(G1338gat));
  NOR2_X1   g554(.A1(new_n486), .A2(G106gat), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n679), .A2(new_n369), .A3(new_n680), .A4(new_n726), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT112), .B(G106gat), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n740), .A2(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT113), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n733), .B(KEYINPUT51), .C1(new_n677), .C2(new_n725), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n762), .A2(new_n645), .A3(new_n731), .A4(new_n756), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(KEYINPUT114), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n740), .A2(new_n765), .A3(new_n756), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n757), .A2(new_n758), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n764), .A2(new_n766), .A3(new_n760), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n763), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n770), .A3(KEYINPUT53), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n761), .A2(new_n768), .A3(new_n771), .ZN(G1339gat));
  AOI21_X1  g571(.A(new_n639), .B1(new_n594), .B2(new_n631), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n628), .B1(new_n638), .B2(new_n624), .ZN(new_n774));
  INV_X1    g573(.A(new_n629), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT54), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT55), .B1(new_n777), .B2(new_n633), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n632), .B1(new_n774), .B2(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n779), .A2(new_n780), .A3(new_n639), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n617), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n644), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n616), .B1(new_n633), .B2(new_n780), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n776), .B(KEYINPUT54), .C1(new_n643), .C2(new_n619), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT55), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n264), .A2(new_n250), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n249), .A2(new_n251), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n205), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n274), .A2(new_n557), .A3(new_n558), .A4(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n783), .A2(new_n786), .A3(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n274), .A2(new_n789), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n645), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n785), .A2(KEYINPUT55), .A3(new_n617), .A4(new_n781), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(new_n275), .A3(new_n644), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n786), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n791), .B1(new_n796), .B2(new_n559), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n784), .A2(new_n785), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n644), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n779), .A2(new_n639), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n780), .B1(new_n630), .B2(new_n773), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n801), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n803), .B1(new_n806), .B2(new_n784), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n807), .A3(new_n275), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n669), .B1(new_n808), .B2(new_n793), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT115), .B1(new_n809), .B2(new_n791), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n799), .A2(new_n810), .A3(new_n670), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n613), .A2(new_n275), .A3(new_n645), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n369), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n510), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n513), .A2(new_n439), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818), .B2(new_n275), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n815), .A2(new_n478), .A3(new_n440), .ZN(new_n820));
  INV_X1    g619(.A(G113gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n820), .A2(new_n821), .A3(new_n276), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(G1340gat));
  AOI21_X1  g622(.A(G120gat), .B1(new_n818), .B2(new_n645), .ZN(new_n824));
  INV_X1    g623(.A(G120gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n820), .A2(new_n825), .A3(new_n671), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(G1341gat));
  NAND3_X1  g626(.A1(new_n818), .A2(new_n598), .A3(new_n682), .ZN(new_n828));
  OAI21_X1  g627(.A(G127gat), .B1(new_n820), .B2(new_n670), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1342gat));
  NAND2_X1  g629(.A1(new_n669), .A2(new_n553), .ZN(new_n831));
  OR3_X1    g630(.A1(new_n817), .A2(KEYINPUT56), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G134gat), .B1(new_n820), .B2(new_n559), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT56), .B1(new_n817), .B2(new_n831), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(G1343gat));
  INV_X1    g634(.A(G141gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n440), .A2(new_n510), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n658), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n791), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n800), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n784), .A2(KEYINPUT118), .A3(new_n785), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n801), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n795), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n844), .A2(new_n845), .B1(new_n645), .B2(new_n792), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(new_n669), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n812), .B1(new_n847), .B2(new_n670), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n848), .A2(new_n849), .A3(new_n486), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n670), .B1(new_n797), .B2(new_n798), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n809), .A2(KEYINPUT115), .A3(new_n791), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n813), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n852), .B1(new_n855), .B2(new_n369), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n850), .B1(new_n856), .B2(KEYINPUT117), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n486), .B1(new_n811), .B2(new_n813), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n858), .B1(new_n859), .B2(new_n852), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n839), .B1(new_n857), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n836), .B1(new_n861), .B2(new_n275), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n855), .A2(new_n369), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n839), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n864), .A2(new_n836), .A3(new_n275), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT58), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n863), .A2(KEYINPUT117), .A3(new_n851), .ZN(new_n868));
  INV_X1    g667(.A(new_n850), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n860), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n275), .A3(new_n838), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G141gat), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(new_n865), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n867), .A2(new_n874), .ZN(G1344gat));
  INV_X1    g674(.A(G148gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n864), .A2(new_n876), .A3(new_n645), .ZN(new_n877));
  XOR2_X1   g676(.A(new_n877), .B(KEYINPUT119), .Z(new_n878));
  AOI211_X1 g677(.A(KEYINPUT59), .B(new_n876), .C1(new_n861), .C2(new_n645), .ZN(new_n879));
  XNOR2_X1  g678(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n849), .B1(new_n848), .B2(new_n486), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n863), .B2(new_n851), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n645), .B1(new_n838), .B2(KEYINPUT121), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n883), .B1(KEYINPUT121), .B2(new_n838), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n878), .B1(new_n879), .B2(new_n886), .ZN(G1345gat));
  AOI21_X1  g686(.A(new_n294), .B1(new_n864), .B2(new_n682), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n682), .A2(new_n294), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n889), .B(KEYINPUT122), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n861), .B2(new_n890), .ZN(G1346gat));
  INV_X1    g690(.A(new_n295), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n864), .A2(new_n892), .A3(new_n669), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n861), .A2(new_n669), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n892), .ZN(G1347gat));
  NAND2_X1  g694(.A1(new_n439), .A2(new_n330), .ZN(new_n896));
  INV_X1    g695(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n478), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n898), .B(KEYINPUT123), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n814), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(G169gat), .B1(new_n900), .B2(new_n276), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n487), .B(new_n896), .C1(new_n811), .C2(new_n813), .ZN(new_n902));
  INV_X1    g701(.A(new_n386), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n275), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n901), .A2(new_n904), .ZN(G1348gat));
  OAI21_X1  g704(.A(G176gat), .B1(new_n900), .B2(new_n671), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n387), .A3(new_n645), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1349gat));
  OAI21_X1  g707(.A(G183gat), .B1(new_n900), .B2(new_n670), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n902), .A2(new_n371), .A3(new_n682), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n902), .A2(new_n372), .A3(new_n669), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n814), .A2(new_n669), .A3(new_n899), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n914), .A2(new_n915), .A3(G190gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n915), .B1(new_n914), .B2(G190gat), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT124), .ZN(G1351gat));
  INV_X1    g718(.A(G197gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n659), .A2(new_n897), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT125), .Z(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n275), .A3(new_n882), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n920), .B1(new_n923), .B2(KEYINPUT126), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n924), .B1(KEYINPUT126), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n863), .A2(new_n921), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n920), .A3(new_n275), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(G1352gat));
  INV_X1    g727(.A(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(new_n929), .A3(new_n645), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT62), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n922), .A2(new_n882), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(new_n645), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n931), .A2(new_n933), .ZN(G1353gat));
  NAND3_X1  g733(.A1(new_n926), .A2(new_n334), .A3(new_n682), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n882), .A2(new_n659), .A3(new_n682), .A4(new_n897), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n936), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT63), .B1(new_n936), .B2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n935), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(new_n669), .B1(new_n932), .B2(KEYINPUT127), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n922), .A2(KEYINPUT127), .A3(new_n882), .ZN(new_n941));
  OAI21_X1  g740(.A(G218gat), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n926), .A2(new_n335), .A3(new_n669), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(G1355gat));
endmodule


