//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:05 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(G143), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  OR2_X1    g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT0), .A3(G128), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  INV_X1    g012(.A(G134), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G137), .ZN(new_n200));
  INV_X1    g014(.A(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT11), .A3(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n199), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G131), .ZN(new_n205));
  INV_X1    g019(.A(G131), .ZN(new_n206));
  NAND4_X1  g020(.A1(new_n200), .A2(new_n202), .A3(new_n206), .A4(new_n203), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n197), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n195), .A2(new_n210), .A3(G128), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(KEYINPUT65), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n189), .B(G146), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n191), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n211), .A2(new_n215), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n199), .A2(G137), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n201), .A2(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n207), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n209), .A2(new_n223), .A3(KEYINPUT30), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G116), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G119), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT2), .B(G113), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT2), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G113), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n224), .A2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n207), .A2(new_n221), .A3(KEYINPUT64), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT64), .B1(new_n207), .B2(new_n221), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n218), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT66), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n245), .B(new_n218), .C1(new_n241), .C2(new_n242), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n246), .A3(new_n209), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n240), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n239), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n209), .A2(new_n250), .A3(new_n223), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NOR2_X1   g066(.A1(G237), .A2(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G210), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT67), .B1(new_n249), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT67), .ZN(new_n260));
  INV_X1    g074(.A(new_n257), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n251), .A2(new_n261), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n243), .A2(KEYINPUT66), .B1(new_n208), .B2(new_n197), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT30), .B1(new_n263), .B2(new_n246), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n260), .B(new_n262), .C1(new_n264), .C2(new_n240), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n259), .A2(KEYINPUT31), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n252), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n251), .B1(new_n247), .B2(new_n239), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(new_n267), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n261), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n247), .A2(new_n248), .ZN(new_n272));
  INV_X1    g086(.A(new_n240), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n258), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n266), .A2(new_n271), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(G472), .ZN(new_n278));
  INV_X1    g092(.A(G902), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT32), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(G472), .A2(G902), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(new_n281), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n261), .B1(new_n252), .B2(new_n267), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n269), .B2(new_n267), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n261), .B1(new_n249), .B2(new_n251), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n209), .A2(new_n223), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(new_n239), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n289), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n293));
  AOI21_X1  g107(.A(G902), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n277), .A2(new_n285), .B1(new_n295), .B2(G472), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n282), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G469), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n189), .A2(KEYINPUT1), .A3(G146), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n211), .A2(new_n217), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G104), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT3), .B1(new_n301), .B2(G107), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n303));
  INV_X1    g117(.A(G107), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(G104), .ZN(new_n305));
  INV_X1    g119(.A(G101), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n301), .A2(G107), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n302), .A2(new_n305), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n301), .A2(G107), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n304), .A2(G104), .ZN(new_n310));
  OAI21_X1  g124(.A(G101), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AND2_X1   g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n300), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT10), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n308), .A2(new_n311), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n315), .A2(new_n314), .ZN(new_n316));
  AOI22_X1  g130(.A1(new_n313), .A2(new_n314), .B1(new_n316), .B2(new_n218), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n302), .A2(new_n305), .A3(new_n307), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G101), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n308), .A2(KEYINPUT4), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(KEYINPUT71), .A3(G101), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT4), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n325), .A3(G101), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n197), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n208), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G110), .B(G140), .ZN(new_n330));
  INV_X1    g144(.A(G953), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n331), .A2(G227), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT12), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n315), .A2(new_n217), .A3(new_n211), .A4(new_n215), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n336), .B(new_n328), .C1(new_n313), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n313), .A2(new_n337), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT12), .B1(new_n339), .B2(new_n208), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n335), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n317), .A2(new_n327), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n208), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n334), .B1(new_n344), .B2(new_n329), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n298), .B(new_n279), .C1(new_n342), .C2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n329), .B1(new_n338), .B2(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n333), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n334), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n344), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT72), .B1(new_n329), .B2(new_n334), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n348), .B(G469), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(G469), .A2(G902), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n346), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G140), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G125), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G140), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT16), .ZN(new_n359));
  OR3_X1    g173(.A1(new_n357), .A2(KEYINPUT16), .A3(G140), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n187), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n360), .A3(G146), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n225), .A2(G128), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n216), .A2(KEYINPUT23), .A3(G119), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n225), .A2(G128), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n365), .B(new_n366), .C1(new_n367), .C2(KEYINPUT23), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT24), .B(G110), .Z(new_n369));
  XNOR2_X1  g183(.A(G119), .B(G128), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n368), .A2(G110), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT69), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n356), .A2(new_n358), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(G146), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n356), .A2(new_n358), .A3(KEYINPUT69), .A4(new_n187), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT68), .B(G110), .ZN(new_n378));
  OAI22_X1  g192(.A1(new_n368), .A2(new_n378), .B1(new_n369), .B2(new_n370), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(new_n379), .A3(new_n363), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT22), .B(G137), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n331), .A2(G221), .A3(G234), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n372), .A2(new_n380), .A3(new_n384), .ZN(new_n387));
  INV_X1    g201(.A(G234), .ZN(new_n388));
  AOI21_X1  g202(.A(G902), .B1(new_n388), .B2(G217), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT70), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n386), .A2(new_n279), .A3(new_n387), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n392), .A2(KEYINPUT25), .ZN(new_n393));
  OAI21_X1  g207(.A(G217), .B1(new_n388), .B2(G902), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n394), .B1(new_n392), .B2(KEYINPUT25), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT9), .B(G234), .ZN(new_n397));
  OAI21_X1  g211(.A(G221), .B1(new_n397), .B2(G902), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n354), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(G214), .B1(G237), .B2(G902), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT73), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n197), .A2(new_n357), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n218), .A2(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g218(.A(KEYINPUT78), .B(G224), .Z(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n331), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT77), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n404), .B(new_n407), .ZN(new_n408));
  AND3_X1   g222(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT5), .ZN(new_n409));
  OAI21_X1  g223(.A(G113), .B1(new_n226), .B2(KEYINPUT5), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n238), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(new_n315), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G122), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n318), .A2(KEYINPUT71), .A3(G101), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT71), .B1(new_n318), .B2(G101), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n308), .A2(KEYINPUT4), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n239), .A2(new_n326), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n413), .B(new_n414), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT75), .ZN(new_n421));
  INV_X1    g235(.A(new_n414), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n239), .A2(new_n326), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n412), .B1(new_n324), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g240(.A(KEYINPUT74), .B(new_n412), .C1(new_n324), .C2(new_n423), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n421), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT74), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n424), .A2(new_n425), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT75), .A4(new_n422), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(KEYINPUT6), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n426), .A2(new_n427), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT6), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT76), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT76), .ZN(new_n437));
  NOR4_X1   g251(.A1(new_n426), .A2(new_n427), .A3(new_n437), .A4(KEYINPUT6), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n408), .B(new_n433), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n402), .A2(new_n403), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT80), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(new_n406), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n441), .B2(new_n406), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT81), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n312), .A2(KEYINPUT79), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n446), .A2(new_n411), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n414), .B(KEYINPUT8), .Z(new_n448));
  AOI21_X1  g262(.A(new_n448), .B1(new_n446), .B2(new_n411), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n406), .A2(KEYINPUT7), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n447), .A2(new_n449), .B1(new_n404), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n440), .A2(new_n452), .A3(new_n443), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n445), .A2(new_n420), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n454), .A2(new_n279), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n439), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n439), .A2(new_n457), .A3(new_n455), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n401), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G113), .B(G122), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(new_n301), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n331), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n189), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n253), .A2(G143), .A3(G214), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n206), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT83), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n467), .A2(new_n189), .ZN(new_n472));
  AOI21_X1  g286(.A(G143), .B1(new_n253), .B2(G214), .ZN(new_n473));
  OAI21_X1  g287(.A(G131), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT83), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n468), .A2(new_n475), .A3(new_n206), .A4(new_n469), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(new_n374), .B(KEYINPUT19), .Z(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(new_n187), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n477), .A2(new_n363), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n374), .A2(G146), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n377), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n468), .A2(new_n469), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n468), .B2(new_n469), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n465), .B1(new_n480), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT17), .B(G131), .C1(new_n472), .C2(new_n473), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n362), .A2(new_n489), .A3(new_n363), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n471), .A2(new_n474), .A3(new_n491), .A4(new_n476), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n493), .A2(new_n487), .A3(new_n465), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(KEYINPUT84), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n490), .A2(new_n492), .B1(new_n482), .B2(new_n486), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n465), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n488), .B1(new_n495), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g313(.A1(G475), .A2(G902), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n500), .B(KEYINPUT85), .Z(new_n501));
  OAI21_X1  g315(.A(new_n463), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n480), .A2(new_n487), .ZN(new_n503));
  INV_X1    g317(.A(new_n465), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND4_X1   g319(.A1(new_n497), .A2(new_n493), .A3(new_n487), .A4(new_n465), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n497), .B1(new_n496), .B2(new_n465), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  INV_X1    g323(.A(new_n501), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OR2_X1    g325(.A1(new_n496), .A2(new_n465), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n512), .B1(new_n506), .B2(new_n507), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n279), .ZN(new_n514));
  AOI22_X1  g328(.A1(new_n502), .A2(new_n511), .B1(new_n514), .B2(G475), .ZN(new_n515));
  INV_X1    g329(.A(G217), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n397), .A2(new_n516), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n227), .B2(G122), .ZN(new_n520));
  INV_X1    g334(.A(G122), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(KEYINPUT86), .A3(G116), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n521), .A2(G116), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n304), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n189), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n216), .A2(G143), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n199), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n530), .A2(G134), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n526), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT14), .B1(new_n521), .B2(G116), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n521), .A2(KEYINPUT86), .A3(G116), .ZN(new_n534));
  AOI21_X1  g348(.A(KEYINPUT86), .B1(new_n521), .B2(G116), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT87), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT87), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n523), .A2(new_n538), .A3(new_n533), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT14), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n524), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n532), .B1(new_n542), .B2(G107), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT13), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n528), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n530), .A2(new_n545), .A3(G134), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n527), .B(new_n528), .C1(new_n544), .C2(new_n199), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n523), .A2(new_n525), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(G107), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n548), .B1(new_n550), .B2(new_n526), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n518), .B1(new_n543), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT88), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n526), .ZN(new_n554));
  INV_X1    g368(.A(new_n548), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n536), .A2(KEYINPUT87), .B1(new_n540), .B2(new_n524), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n304), .B1(new_n557), .B2(new_n539), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n556), .B(new_n517), .C1(new_n558), .C2(new_n532), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n553), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT88), .B(new_n518), .C1(new_n543), .C2(new_n551), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n279), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(G478), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT89), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT89), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n567), .A3(new_n564), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n564), .B(KEYINPUT90), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n560), .A2(new_n279), .A3(new_n561), .A4(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT91), .ZN(new_n572));
  NOR2_X1   g386(.A1(KEYINPUT92), .A2(G952), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(KEYINPUT92), .A2(G952), .ZN(new_n575));
  AOI21_X1  g389(.A(G953), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n388), .B2(new_n466), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT21), .B(G898), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n279), .B(new_n331), .C1(G234), .C2(G237), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  AND4_X1   g396(.A1(new_n515), .A2(new_n569), .A3(new_n572), .A4(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n297), .A2(new_n399), .A3(new_n461), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT93), .B(G101), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n584), .B(new_n585), .ZN(G3));
  AND3_X1   g400(.A1(new_n439), .A2(new_n457), .A3(new_n455), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n457), .B1(new_n439), .B2(new_n455), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n400), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT94), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n459), .A2(new_n460), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n592), .A3(new_n400), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n560), .A2(new_n595), .A3(new_n561), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n552), .A2(KEYINPUT33), .A3(new_n559), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n596), .A2(G478), .A3(new_n279), .A4(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n562), .A2(new_n563), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n599), .B1(new_n598), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(new_n515), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n582), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n270), .A2(new_n261), .B1(new_n274), .B2(new_n275), .ZN(new_n607));
  AOI211_X1 g421(.A(G472), .B(G902), .C1(new_n607), .C2(new_n266), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n278), .B1(new_n277), .B2(new_n279), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n354), .A2(new_n396), .A3(new_n398), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n594), .A2(new_n606), .A3(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(new_n612), .B(KEYINPUT96), .Z(new_n613));
  XOR2_X1   g427(.A(KEYINPUT34), .B(G104), .Z(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n568), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n567), .B1(new_n562), .B2(new_n564), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n571), .A2(KEYINPUT91), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n571), .A2(KEYINPUT91), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n616), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n514), .A2(G475), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n508), .A2(new_n462), .A3(new_n510), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n502), .A2(new_n622), .A3(KEYINPUT97), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n499), .A2(new_n463), .A3(new_n501), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n462), .B1(new_n508), .B2(new_n510), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n620), .A2(new_n621), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  OAI21_X1  g442(.A(KEYINPUT98), .B1(new_n628), .B2(new_n581), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n623), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n569), .A2(new_n572), .B1(G475), .B2(new_n514), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .A4(new_n582), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n594), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n611), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NOR2_X1   g453(.A1(new_n608), .A2(new_n609), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n393), .A2(new_n395), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n385), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n381), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n389), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n354), .A2(new_n398), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n640), .A2(new_n461), .A3(new_n583), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  INV_X1    g464(.A(G900), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n578), .B1(new_n651), .B2(new_n580), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n628), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n590), .A2(new_n593), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n354), .A2(new_n398), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(G902), .B1(new_n607), .B2(new_n266), .ZN(new_n657));
  AOI21_X1  g471(.A(KEYINPUT32), .B1(new_n657), .B2(new_n278), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n277), .A2(new_n285), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n295), .A2(G472), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(new_n656), .B(new_n645), .C1(new_n658), .C2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n216), .ZN(G30));
  XOR2_X1   g478(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n591), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n652), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n656), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  INV_X1    g483(.A(new_n620), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n515), .ZN(new_n671));
  INV_X1    g485(.A(new_n400), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n645), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n259), .A2(new_n265), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n261), .B2(new_n292), .ZN(new_n676));
  OAI21_X1  g490(.A(G472), .B1(new_n676), .B2(G902), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n282), .A2(new_n659), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n666), .A2(new_n674), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n189), .ZN(G45));
  NAND2_X1  g496(.A1(new_n502), .A2(new_n511), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n621), .ZN(new_n684));
  INV_X1    g498(.A(new_n652), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n684), .B(new_n685), .C1(new_n601), .C2(new_n602), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n590), .A2(new_n593), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n688), .A2(new_n662), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT101), .B(G146), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G48));
  OAI21_X1  g505(.A(new_n396), .B1(new_n658), .B2(new_n661), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n342), .A2(new_n345), .ZN(new_n693));
  OAI21_X1  g507(.A(G469), .B1(new_n693), .B2(G902), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n398), .A3(new_n346), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n594), .A2(new_n696), .A3(new_n606), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT41), .B(G113), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G15));
  NAND2_X1  g513(.A1(new_n636), .A2(new_n696), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  INV_X1    g515(.A(new_n645), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n282), .B2(new_n296), .ZN(new_n703));
  INV_X1    g517(.A(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n594), .A2(new_n583), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G119), .ZN(G21));
  NOR2_X1   g520(.A1(new_n695), .A2(new_n581), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n593), .A2(new_n590), .A3(new_n671), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n292), .A2(KEYINPUT28), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n257), .B1(new_n709), .B2(new_n268), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n710), .B1(new_n275), .B2(new_n274), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n284), .B1(new_n711), .B2(new_n266), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n277), .A2(new_n279), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(KEYINPUT102), .A3(G472), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n657), .B2(new_n278), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n712), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT103), .B1(new_n717), .B2(new_n396), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n716), .ZN(new_n719));
  INV_X1    g533(.A(new_n712), .ZN(new_n720));
  AND4_X1   g534(.A1(KEYINPUT103), .A2(new_n719), .A3(new_n396), .A4(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n708), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT104), .B(G122), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G24));
  NAND4_X1  g538(.A1(new_n590), .A2(new_n593), .A3(new_n687), .A4(new_n704), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n609), .A2(KEYINPUT102), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n657), .A2(new_n715), .A3(new_n278), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n645), .B(new_n720), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT105), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT105), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n717), .A2(new_n730), .A3(new_n645), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n725), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT106), .B(G125), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G27));
  XOR2_X1   g548(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n587), .A2(new_n588), .A3(new_n672), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT108), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n352), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT72), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n335), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(new_n344), .A3(new_n349), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n742), .A2(KEYINPUT108), .A3(G469), .A4(new_n348), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n353), .B(KEYINPUT107), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n739), .A2(new_n743), .A3(new_n346), .A4(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n745), .A2(new_n398), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n737), .A2(new_n687), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n736), .B1(new_n747), .B2(new_n692), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n459), .A2(new_n460), .A3(new_n400), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n745), .A2(new_n398), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n686), .ZN(new_n751));
  INV_X1    g565(.A(new_n396), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n752), .B1(new_n282), .B2(new_n296), .ZN(new_n753));
  NOR2_X1   g567(.A1(KEYINPUT109), .A2(KEYINPUT42), .ZN(new_n754));
  INV_X1    g568(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n751), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n748), .A2(new_n756), .A3(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n757), .B1(new_n748), .B2(new_n756), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XOR2_X1   g575(.A(KEYINPUT111), .B(G131), .Z(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G33));
  NAND3_X1  g577(.A1(new_n653), .A2(new_n737), .A3(new_n746), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n692), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n199), .ZN(G36));
  NAND2_X1  g580(.A1(new_n742), .A2(new_n348), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n298), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n768), .B2(new_n767), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n744), .ZN(new_n771));
  OR2_X1    g585(.A1(new_n771), .A2(KEYINPUT46), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(KEYINPUT46), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n346), .A3(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n398), .A3(new_n667), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n684), .B1(new_n603), .B2(KEYINPUT113), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(KEYINPUT113), .B2(new_n603), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n603), .B1(new_n780), .B2(new_n684), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n780), .B2(new_n684), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n779), .A2(KEYINPUT43), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT43), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n640), .A2(new_n702), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  AOI211_X1 g603(.A(new_n749), .B(new_n775), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NAND2_X1  g607(.A1(new_n774), .A2(new_n398), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n774), .A2(KEYINPUT47), .A3(new_n398), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n297), .A2(new_n749), .A3(new_n396), .A4(new_n686), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NAND2_X1  g615(.A1(new_n694), .A2(new_n346), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n802), .A2(KEYINPUT49), .ZN(new_n804));
  INV_X1    g618(.A(new_n401), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n396), .A2(new_n398), .A3(new_n805), .ZN(new_n806));
  NOR4_X1   g620(.A1(new_n782), .A2(new_n803), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(new_n679), .A3(new_n666), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n594), .B(new_n696), .C1(new_n635), .C2(new_n606), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n705), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n590), .A2(new_n593), .A3(new_n671), .A4(new_n707), .ZN(new_n812));
  INV_X1    g626(.A(new_n718), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n717), .A2(KEYINPUT103), .A3(new_n396), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT115), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  AND4_X1   g630(.A1(new_n730), .A2(new_n719), .A3(new_n645), .A4(new_n720), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n730), .B1(new_n717), .B2(new_n645), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n751), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n749), .A2(new_n628), .A3(new_n750), .A4(new_n652), .ZN(new_n820));
  INV_X1    g634(.A(new_n662), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n569), .A2(new_n572), .A3(new_n621), .A4(new_n685), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n630), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n737), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n820), .A2(new_n753), .B1(new_n821), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n713), .A2(G472), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n399), .A3(new_n280), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n805), .B(new_n582), .C1(new_n587), .C2(new_n588), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n620), .A2(new_n515), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n591), .A2(new_n805), .A3(new_n583), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n646), .A3(new_n280), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n828), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n830), .A2(new_n831), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n603), .B2(new_n515), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT116), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n684), .B(new_n840), .C1(new_n601), .C2(new_n602), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n805), .B1(new_n587), .B2(new_n588), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n515), .A2(new_n569), .A3(new_n572), .A4(new_n582), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n610), .A3(new_n844), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n838), .A2(new_n842), .B1(new_n845), .B2(new_n297), .ZN(new_n846));
  INV_X1    g660(.A(new_n832), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n611), .A2(new_n461), .A3(new_n582), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(KEYINPUT117), .A3(new_n647), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n837), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n827), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n722), .A2(new_n852), .A3(new_n810), .A4(new_n705), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n816), .A2(new_n851), .A3(new_n761), .A4(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n594), .B(new_n821), .C1(new_n653), .C2(new_n687), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n750), .A2(new_n645), .A3(new_n652), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n594), .A2(new_n678), .A3(new_n671), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n817), .A2(new_n818), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n855), .B(new_n857), .C1(new_n858), .C2(new_n725), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT52), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n662), .B1(new_n688), .B2(new_n654), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n732), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n863), .A3(new_n857), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n809), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n809), .B1(new_n748), .B2(new_n756), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n722), .A2(new_n868), .A3(new_n705), .A4(new_n810), .ZN(new_n869));
  OAI22_X1  g683(.A1(new_n764), .A2(new_n692), .B1(new_n662), .B2(new_n824), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n729), .A2(new_n731), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n870), .B1(new_n871), .B2(new_n751), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT117), .B1(new_n848), .B2(new_n647), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n611), .A2(new_n461), .A3(new_n582), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n839), .A2(new_n841), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n584), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n872), .A2(new_n877), .A3(new_n849), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n869), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT118), .A4(new_n849), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n880), .A2(new_n860), .A3(new_n864), .A4(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n866), .A2(new_n867), .A3(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n860), .A2(new_n864), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n816), .A2(new_n853), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n759), .A2(new_n760), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n878), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT53), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n883), .B1(new_n889), .B2(new_n867), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n783), .A2(new_n578), .A3(new_n786), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n594), .A2(new_n704), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n813), .A2(new_n814), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n749), .A2(new_n695), .ZN(new_n895));
  AND4_X1   g709(.A1(new_n396), .A2(new_n679), .A3(new_n578), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n604), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n894), .A2(new_n576), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n891), .A2(new_n895), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n899), .A2(KEYINPUT48), .A3(new_n692), .ZN(new_n900));
  OAI21_X1  g714(.A(KEYINPUT48), .B1(new_n899), .B2(new_n692), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n695), .A2(new_n400), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n891), .A2(new_n666), .A3(new_n893), .A4(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT50), .Z(new_n905));
  OAI211_X1 g719(.A(new_n796), .B(new_n797), .C1(new_n398), .C2(new_n802), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(new_n893), .A3(new_n737), .A4(new_n891), .ZN(new_n907));
  AND3_X1   g721(.A1(new_n896), .A2(new_n515), .A3(new_n603), .ZN(new_n908));
  INV_X1    g722(.A(new_n899), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n871), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n905), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n902), .B1(new_n911), .B2(KEYINPUT51), .ZN(new_n912));
  AND4_X1   g726(.A1(KEYINPUT51), .A2(new_n905), .A3(new_n907), .A4(new_n910), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n890), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(G952), .A2(G953), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n808), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n331), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n879), .B1(new_n827), .B2(new_n850), .ZN(new_n919));
  AND4_X1   g733(.A1(new_n705), .A2(new_n722), .A3(new_n868), .A4(new_n810), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n920), .A3(new_n881), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(new_n865), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n888), .B2(new_n809), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n279), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n433), .B1(new_n436), .B2(new_n438), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n408), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n918), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n924), .A2(G210), .ZN(new_n930));
  XOR2_X1   g744(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(KEYINPUT120), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT120), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n930), .A2(new_n934), .A3(new_n931), .A4(new_n928), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n929), .B1(new_n933), .B2(new_n935), .ZN(G51));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n937));
  NOR3_X1   g751(.A1(new_n923), .A2(new_n279), .A3(new_n770), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n744), .B(KEYINPUT57), .Z(new_n939));
  AND3_X1   g753(.A1(new_n866), .A2(new_n867), .A3(new_n882), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n867), .B1(new_n866), .B2(new_n882), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(new_n693), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n938), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n937), .B1(new_n944), .B2(new_n917), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n866), .A2(new_n882), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT54), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n883), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n693), .B1(new_n948), .B2(new_n939), .ZN(new_n949));
  OAI211_X1 g763(.A(KEYINPUT121), .B(new_n918), .C1(new_n949), .C2(new_n938), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n945), .A2(new_n950), .ZN(G54));
  NAND3_X1  g765(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n952), .A2(new_n499), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n499), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n917), .ZN(G60));
  NAND2_X1  g769(.A1(new_n596), .A2(new_n597), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT122), .Z(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT59), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n957), .B1(new_n890), .B2(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n948), .A2(new_n957), .A3(new_n959), .ZN(new_n961));
  NOR3_X1   g775(.A1(new_n960), .A2(new_n917), .A3(new_n961), .ZN(G63));
  NAND2_X1  g776(.A1(G217), .A2(G902), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT60), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT123), .B1(new_n923), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT123), .ZN(new_n966));
  INV_X1    g780(.A(new_n964), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n946), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n386), .A2(new_n387), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT124), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n965), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n966), .B1(new_n946), .B2(new_n967), .ZN(new_n972));
  AOI211_X1 g786(.A(KEYINPUT123), .B(new_n964), .C1(new_n866), .C2(new_n882), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n643), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n971), .A2(new_n974), .A3(new_n918), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n971), .A2(new_n974), .A3(KEYINPUT61), .A4(new_n918), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(G66));
  INV_X1    g793(.A(new_n579), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n331), .B1(new_n980), .B2(new_n405), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n885), .A2(new_n849), .A3(new_n877), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n331), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n926), .B1(G898), .B2(new_n331), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n983), .B(new_n984), .Z(G69));
  AOI22_X1  g799(.A1(new_n790), .A2(new_n791), .B1(new_n798), .B2(new_n799), .ZN(new_n986));
  INV_X1    g800(.A(new_n681), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n862), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NOR3_X1   g803(.A1(new_n692), .A2(new_n668), .A3(new_n749), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n990), .B1(new_n847), .B2(new_n842), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n986), .A2(new_n989), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n331), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n272), .A2(new_n224), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(new_n478), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(new_n996), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n331), .A2(G900), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n594), .A2(new_n671), .A3(new_n753), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n775), .A2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n1001), .A2(new_n886), .A3(new_n765), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n986), .A2(new_n1002), .A3(new_n862), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n999), .B1(new_n1003), .B2(new_n331), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n998), .B1(new_n1004), .B2(KEYINPUT125), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT125), .ZN(new_n1006));
  AOI211_X1 g820(.A(new_n1006), .B(new_n999), .C1(new_n1003), .C2(new_n331), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n997), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n331), .B1(G227), .B2(G900), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1009), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1011), .B(new_n997), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1010), .A2(new_n1012), .ZN(G72));
  NAND2_X1  g827(.A1(G472), .A2(G902), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT63), .Z(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n993), .B2(new_n982), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1016), .B(new_n257), .C1(new_n249), .C2(new_n251), .ZN(new_n1017));
  INV_X1    g831(.A(new_n288), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n675), .B1(KEYINPUT127), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(KEYINPUT127), .B2(new_n1018), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1015), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1017), .B1(new_n889), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1003), .A2(new_n982), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1015), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n252), .B(new_n261), .C1(new_n264), .C2(new_n240), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n918), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1027), .A2(KEYINPUT126), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT126), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1029), .B(new_n918), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1022), .B1(new_n1028), .B2(new_n1030), .ZN(G57));
endmodule


