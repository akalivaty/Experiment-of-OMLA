//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:09 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n565, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n455), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  OAI211_X1 g043(.A(new_n467), .B(G2104), .C1(new_n468), .C2(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n470), .B(KEYINPUT3), .C1(new_n462), .C2(KEYINPUT70), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT69), .B1(new_n468), .B2(G2104), .ZN(new_n472));
  AND3_X1   g047(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(G2104), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT67), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g056(.A(G125), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(KEYINPUT68), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G125), .C1(new_n480), .C2(new_n481), .ZN(new_n485));
  NAND2_X1  g060(.A1(G113), .A2(G2104), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n477), .B1(new_n487), .B2(G2105), .ZN(G160));
  NAND2_X1  g063(.A1(new_n473), .A2(G2105), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT72), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  INV_X1    g066(.A(new_n475), .ZN(new_n492));
  MUX2_X1   g067(.A(G100), .B(G112), .S(G2105), .Z(new_n493));
  AOI22_X1  g068(.A1(new_n492), .A2(G136), .B1(G2104), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n491), .A2(new_n494), .ZN(G162));
  OAI211_X1 g070(.A(G138), .B(new_n474), .C1(new_n480), .C2(new_n481), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT4), .A2(G138), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(G102), .A2(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(new_n474), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n469), .A2(new_n471), .A3(G126), .A4(new_n472), .ZN(new_n504));
  NAND2_X1  g079(.A1(G114), .A2(G2104), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G2105), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n498), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n512), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n515), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n519), .A2(KEYINPUT73), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(new_n526), .A3(new_n518), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n519), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n532));
  INV_X1    g107(.A(new_n512), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n529), .A2(new_n531), .A3(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(G168));
  AND2_X1   g111(.A1(new_n528), .A2(G52), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n512), .A2(new_n519), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n538), .A2(new_n514), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n528), .A2(G43), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n514), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n510), .A2(new_n511), .B1(new_n517), .B2(new_n518), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G81), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  AOI22_X1  g130(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  OAI22_X1  g132(.A1(new_n556), .A2(new_n514), .B1(new_n539), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n528), .A2(G53), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  OR2_X1    g139(.A1(G168), .A2(KEYINPUT74), .ZN(new_n565));
  NAND2_X1  g140(.A1(G168), .A2(KEYINPUT74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G286));
  INV_X1    g143(.A(new_n527), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n526), .B1(new_n517), .B2(new_n518), .ZN(new_n570));
  OAI211_X1 g145(.A(G49), .B(G543), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n510), .A2(new_n572), .A3(new_n511), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n546), .A2(G87), .B1(G651), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n571), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  NAND3_X1  g155(.A1(new_n519), .A2(G48), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n539), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n512), .A2(G61), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n514), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G305));
  NAND2_X1  g163(.A1(G72), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n533), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G85), .B2(new_n546), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n528), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  NOR2_X1   g170(.A1(G301), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n528), .B(KEYINPUT76), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(G54), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n539), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n546), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n533), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n601), .A2(new_n602), .B1(new_n605), .B2(G651), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(new_n595), .ZN(G284));
  AOI21_X1  g183(.A(new_n596), .B1(new_n607), .B2(new_n595), .ZN(G321));
  NAND2_X1  g184(.A1(G299), .A2(new_n595), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n567), .B2(new_n595), .ZN(G297));
  XNOR2_X1  g186(.A(G297), .B(KEYINPUT77), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n607), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n613), .A3(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n549), .A2(new_n595), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT11), .Z(G282));
  INV_X1    g193(.A(new_n617), .ZN(G323));
  INV_X1    g194(.A(KEYINPUT67), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n468), .A2(G2104), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n478), .A2(new_n479), .A3(KEYINPUT67), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n625), .A2(G2104), .A3(new_n474), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(G2100), .ZN(new_n631));
  MUX2_X1   g206(.A(G99), .B(G111), .S(G2105), .Z(new_n632));
  AOI22_X1  g207(.A1(new_n492), .A2(G135), .B1(G2104), .B2(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n634), .B1(new_n490), .B2(G123), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT15), .B(G2435), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2427), .ZN(new_n641));
  INV_X1    g216(.A(G2430), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n644), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n644), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2084), .B(G2090), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT78), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g232(.A1(G2072), .A2(G2078), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n442), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n657), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT81), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n659), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n656), .B(new_n665), .C1(new_n660), .C2(new_n662), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT80), .ZN(new_n667));
  NOR3_X1   g242(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT79), .B(KEYINPUT18), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n664), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2096), .B(G2100), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT82), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(G227));
  XOR2_X1   g249(.A(G1971), .B(G1976), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1956), .B(G2474), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1961), .B(G1966), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT20), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n677), .A2(new_n678), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n676), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(new_n676), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT83), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n685), .B(new_n687), .Z(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G5), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G171), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G1961), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT31), .B(G11), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT30), .B(G28), .Z(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G29), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(new_n635), .B2(G29), .ZN(new_n702));
  INV_X1    g277(.A(G1966), .ZN(new_n703));
  NOR2_X1   g278(.A1(G168), .A2(new_n694), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n694), .B2(G21), .ZN(new_n705));
  OAI211_X1 g280(.A(new_n698), .B(new_n702), .C1(new_n703), .C2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G29), .B2(G32), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n490), .A2(G129), .ZN(new_n709));
  NAND3_X1  g284(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT86), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n712));
  AOI22_X1  g287(.A1(new_n711), .A2(new_n712), .B1(G105), .B2(new_n463), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n712), .B2(new_n711), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G141), .B2(new_n492), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  MUX2_X1   g293(.A(new_n708), .B(new_n707), .S(new_n718), .Z(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT27), .B(G1996), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT24), .B(G34), .Z(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(G29), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G160), .B2(G29), .ZN(new_n723));
  OAI22_X1  g298(.A1(new_n719), .A2(new_n720), .B1(G2084), .B2(new_n723), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n706), .B(new_n724), .C1(G2084), .C2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(new_n720), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT88), .Z(new_n727));
  NAND2_X1  g302(.A1(new_n705), .A2(new_n703), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT89), .Z(new_n729));
  NOR2_X1   g304(.A1(G27), .A2(G29), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G164), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2078), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n717), .A2(G33), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n625), .A2(G127), .ZN(new_n734));
  AND2_X1   g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  OAI21_X1  g310(.A(G2105), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n463), .A2(G103), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT25), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(new_n492), .B2(G139), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(new_n717), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G2072), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n729), .A2(new_n732), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n725), .A2(new_n727), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT90), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT84), .B(G16), .Z(new_n747));
  MUX2_X1   g322(.A(G24), .B(G290), .S(new_n747), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1986), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n747), .A2(G22), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G166), .B2(new_n747), .ZN(new_n751));
  INV_X1    g326(.A(G1971), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  MUX2_X1   g328(.A(G23), .B(new_n575), .S(G16), .Z(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT33), .B(G1976), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(G6), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n587), .B2(G16), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT32), .B(G1981), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n753), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n749), .B1(new_n761), .B2(KEYINPUT34), .ZN(new_n762));
  NOR2_X1   g337(.A1(G25), .A2(G29), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n490), .A2(G119), .ZN(new_n764));
  MUX2_X1   g339(.A(G95), .B(G107), .S(G2105), .Z(new_n765));
  AOI22_X1  g340(.A1(new_n492), .A2(G131), .B1(G2104), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT35), .B(G1991), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n762), .B(new_n771), .C1(KEYINPUT34), .C2(new_n761), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT36), .ZN(new_n773));
  NOR2_X1   g348(.A1(G29), .A2(G35), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G162), .B2(G29), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT92), .Z(new_n776));
  XOR2_X1   g351(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G2090), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n778), .A2(G2090), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n607), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G4), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1348), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n747), .A2(G19), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n549), .B2(new_n747), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G1341), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n782), .B2(new_n783), .ZN(new_n788));
  INV_X1    g363(.A(G20), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n747), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n562), .B2(new_n694), .ZN(new_n792));
  INV_X1    g367(.A(G1956), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n717), .A2(G26), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT28), .Z(new_n796));
  NAND2_X1  g371(.A1(new_n490), .A2(G128), .ZN(new_n797));
  MUX2_X1   g372(.A(G104), .B(G116), .S(G2105), .Z(new_n798));
  AOI22_X1  g373(.A1(new_n492), .A2(G140), .B1(G2104), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n796), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT85), .B(G2067), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n784), .A2(new_n788), .A3(new_n794), .A4(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n779), .A2(new_n780), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g380(.A1(new_n746), .A2(new_n773), .A3(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n598), .A2(new_n606), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n613), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT93), .B(G55), .ZN(new_n811));
  AOI211_X1 g386(.A(new_n524), .B(new_n811), .C1(new_n525), .C2(new_n527), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n813));
  INV_X1    g388(.A(G93), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n813), .A2(new_n514), .B1(new_n539), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n548), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n548), .A2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n810), .B(new_n820), .Z(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n822));
  INV_X1    g397(.A(G860), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(KEYINPUT39), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n817), .A2(new_n823), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(G145));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n741), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n767), .A2(new_n627), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n767), .A2(new_n627), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n490), .A2(G130), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT97), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n490), .A2(new_n837), .A3(G130), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  MUX2_X1   g414(.A(G106), .B(G118), .S(G2105), .Z(new_n840));
  AOI22_X1  g415(.A1(new_n492), .A2(G142), .B1(G2104), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n834), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n843), .A2(new_n833), .A3(new_n832), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n800), .A2(new_n716), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n797), .A2(new_n709), .A3(new_n799), .A4(new_n715), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n508), .B(KEYINPUT95), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n848), .B(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n741), .A2(new_n829), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n845), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n845), .B1(new_n851), .B2(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n831), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G162), .B(G160), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n635), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n851), .A2(new_n852), .ZN(new_n859));
  AND2_X1   g434(.A1(new_n842), .A2(new_n844), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n861), .A2(new_n830), .A3(new_n853), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n856), .A2(new_n858), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT98), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n856), .A2(new_n865), .A3(new_n858), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n858), .B1(new_n856), .B2(new_n862), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n868), .A2(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n607), .A2(new_n613), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n820), .B(new_n873), .Z(new_n874));
  OAI21_X1  g449(.A(KEYINPUT99), .B1(new_n607), .B2(G299), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n808), .A2(new_n876), .A3(new_n562), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n607), .A2(G299), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT100), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n879), .A2(KEYINPUT41), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n881), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G303), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(new_n575), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n888), .B(new_n889), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n891), .A2(KEYINPUT101), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT42), .Z(new_n893));
  NOR2_X1   g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n887), .A2(new_n893), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n595), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n817), .A2(new_n595), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n872), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n896), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n894), .ZN(new_n902));
  OAI211_X1 g477(.A(KEYINPUT102), .B(new_n898), .C1(new_n902), .C2(new_n595), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(G295));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n897), .B2(new_n899), .ZN(new_n906));
  OAI211_X1 g481(.A(KEYINPUT103), .B(new_n898), .C1(new_n902), .C2(new_n595), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G331));
  NOR2_X1   g483(.A1(G171), .A2(new_n535), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n565), .A2(G171), .A3(new_n566), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n820), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n911), .A2(new_n818), .A3(new_n819), .A4(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT105), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT105), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n820), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n914), .A2(new_n915), .ZN(new_n920));
  OAI22_X1  g495(.A1(new_n919), .A2(new_n886), .B1(new_n882), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n890), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n879), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n884), .A3(new_n885), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n891), .A3(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n926));
  INV_X1    g501(.A(G37), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n922), .A2(new_n925), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT106), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n884), .A2(new_n885), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n930), .A2(new_n920), .B1(new_n919), .B2(new_n879), .ZN(new_n931));
  AOI21_X1  g506(.A(G37), .B1(new_n931), .B2(new_n891), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n933), .A3(new_n926), .A4(new_n922), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n931), .A2(new_n891), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n932), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n939), .A2(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n922), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n926), .A3(new_n932), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(KEYINPUT44), .B2(new_n944), .ZN(G397));
  XOR2_X1   g520(.A(KEYINPUT107), .B(G1384), .Z(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n508), .A2(KEYINPUT108), .A3(KEYINPUT45), .A4(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n485), .A2(new_n486), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n484), .B1(new_n625), .B2(G125), .ZN(new_n954));
  OAI21_X1  g529(.A(G2105), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n477), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(G40), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n508), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT56), .B(G2072), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n952), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n955), .A2(G40), .A3(new_n956), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  AOI21_X1  g539(.A(G2105), .B1(new_n500), .B2(new_n501), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n474), .B1(new_n504), .B2(new_n505), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n964), .B(G1384), .C1(new_n967), .C2(new_n498), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT50), .B1(new_n508), .B2(new_n958), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n793), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n562), .B(KEYINPUT57), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G2067), .ZN(new_n976));
  NAND4_X1  g551(.A1(G160), .A2(G40), .A3(new_n958), .A4(new_n508), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  AOI22_X1  g553(.A1(new_n976), .A2(new_n978), .B1(new_n970), .B2(new_n783), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n975), .B1(new_n808), .B2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n973), .A2(new_n962), .A3(new_n971), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(new_n981), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT61), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n975), .A2(KEYINPUT61), .A3(new_n981), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n963), .A2(new_n958), .A3(new_n976), .A4(new_n508), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n508), .A2(new_n958), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n964), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n508), .A2(KEYINPUT50), .A3(new_n958), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n957), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n987), .B(KEYINPUT60), .C1(new_n991), .C2(G1348), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n992), .A2(KEYINPUT118), .A3(new_n607), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT118), .B1(new_n992), .B2(new_n607), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n992), .A2(new_n607), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n979), .A2(KEYINPUT60), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n985), .B(new_n986), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n999), .A2(KEYINPUT59), .ZN(new_n1000));
  INV_X1    g575(.A(G1996), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n952), .A2(new_n1001), .A3(new_n960), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  XOR2_X1   g578(.A(KEYINPUT58), .B(G1341), .Z(new_n1004));
  NAND2_X1  g579(.A1(new_n977), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n549), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n999), .A2(KEYINPUT59), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI221_X1 g585(.A(new_n549), .B1(new_n999), .B2(KEYINPUT59), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1000), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n982), .B1(new_n998), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2084), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n963), .B(new_n1014), .C1(new_n968), .C2(new_n969), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  AOI211_X1 g591(.A(new_n1016), .B(G1384), .C1(new_n967), .C2(new_n498), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1017), .A2(new_n957), .A3(new_n959), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1018), .B2(G1966), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n535), .A2(G8), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT119), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI211_X1 g598(.A(KEYINPUT51), .B(new_n1021), .C1(new_n1019), .C2(G8), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n988), .A2(new_n1016), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n963), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n703), .B1(new_n1027), .B2(new_n1017), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1025), .B1(new_n1028), .B2(new_n1015), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT51), .B1(new_n1029), .B2(new_n1021), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1024), .B1(KEYINPUT120), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(KEYINPUT51), .C1(new_n1029), .C2(new_n1021), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1023), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT121), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n946), .B1(new_n967), .B2(new_n498), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT108), .B1(new_n1037), .B2(KEYINPUT45), .ZN(new_n1038));
  INV_X1    g613(.A(new_n951), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n508), .A2(new_n947), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1016), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n963), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1036), .B1(new_n1040), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT45), .B1(new_n508), .B2(new_n947), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1044), .ZN(new_n1048));
  NOR3_X1   g623(.A1(new_n957), .A2(new_n1047), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT121), .A3(new_n952), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2078), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n952), .A2(new_n1052), .A3(new_n960), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1053), .A2(new_n1043), .B1(new_n697), .B2(new_n970), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1051), .A2(new_n1054), .A3(G301), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1018), .A2(new_n1044), .ZN(new_n1056));
  AOI21_X1  g631(.A(G301), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1035), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT113), .B(G86), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n581), .B1(new_n539), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(G1981), .B1(new_n1060), .B2(new_n586), .ZN(new_n1061));
  INV_X1    g636(.A(G1981), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT112), .B1(new_n587), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT112), .ZN(new_n1064));
  NOR4_X1   g639(.A1(new_n583), .A2(new_n586), .A3(new_n1064), .A4(G1981), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1061), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI211_X1 g643(.A(KEYINPUT49), .B(new_n1061), .C1(new_n1063), .C2(new_n1065), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1068), .A2(G8), .A3(new_n977), .A4(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n571), .A2(new_n574), .A3(G1976), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1071), .B(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(G8), .C1(new_n957), .C2(new_n988), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  INV_X1    g650(.A(G1976), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n576), .A2(new_n578), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(new_n977), .A3(G8), .A4(new_n1073), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1070), .A2(new_n1075), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1971), .B1(new_n952), .B2(new_n960), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n970), .A2(G2090), .ZN(new_n1083));
  OAI21_X1  g658(.A(G8), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(G303), .A2(G8), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT55), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1081), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n752), .B1(new_n1040), .B2(new_n1027), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT109), .ZN(new_n1089));
  INV_X1    g664(.A(G2090), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n991), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT109), .B1(new_n970), .B2(G2090), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n1086), .B(KEYINPUT110), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(G8), .A3(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1058), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1034), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(G171), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1054), .A2(G301), .A3(new_n1056), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(KEYINPUT54), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(KEYINPUT122), .A3(KEYINPUT54), .A4(new_n1101), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1013), .A2(new_n1098), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1021), .B1(new_n1019), .B2(G8), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT120), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1033), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n1022), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1087), .A2(new_n1095), .A3(new_n1057), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1112), .B2(new_n1022), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT123), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1112), .A2(new_n1022), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT62), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1114), .A4(new_n1115), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n579), .A2(new_n1076), .ZN(new_n1123));
  XNOR2_X1  g698(.A(new_n1123), .B(KEYINPUT114), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1070), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1126), .ZN(new_n1127));
  OAI211_X1 g702(.A(G8), .B(new_n977), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1095), .B2(new_n1081), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1086), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1093), .B2(G8), .ZN(new_n1131));
  OR3_X1    g706(.A1(new_n1131), .A2(KEYINPUT115), .A3(new_n1081), .ZN(new_n1132));
  AND4_X1   g707(.A1(KEYINPUT63), .A2(new_n1095), .A3(new_n567), .A4(new_n1029), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT115), .B1(new_n1131), .B2(new_n1081), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT63), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1029), .A2(new_n567), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1129), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1107), .A2(new_n1118), .A3(new_n1122), .A4(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1042), .A2(new_n957), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n800), .B(new_n976), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n716), .B(new_n1001), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n768), .A2(new_n770), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n768), .A2(new_n770), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  XNOR2_X1  g722(.A(G290), .B(G1986), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1142), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1141), .A2(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1143), .A2(new_n709), .A3(new_n715), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1142), .A2(new_n1001), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1152), .A2(KEYINPUT46), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(KEYINPUT46), .ZN(new_n1154));
  AOI22_X1  g729(.A1(new_n1142), .A2(new_n1151), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT47), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1157));
  OAI22_X1  g732(.A1(new_n1157), .A2(new_n1146), .B1(G2067), .B2(new_n800), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1158), .A2(new_n1142), .ZN(new_n1159));
  NOR2_X1   g734(.A1(G290), .A2(G1986), .ZN(new_n1160));
  AOI21_X1  g735(.A(KEYINPUT48), .B1(new_n1142), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1142), .A2(KEYINPUT48), .A3(new_n1160), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1156), .A2(new_n1159), .A3(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1165), .B(KEYINPUT124), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1150), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT125), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT125), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1150), .A2(new_n1169), .A3(new_n1166), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g746(.A(G227), .ZN(new_n1173));
  NAND4_X1  g747(.A1(new_n692), .A2(G319), .A3(new_n653), .A4(new_n1173), .ZN(new_n1174));
  XOR2_X1   g748(.A(new_n1174), .B(KEYINPUT126), .Z(new_n1175));
  AOI21_X1  g749(.A(new_n1175), .B1(new_n867), .B2(new_n869), .ZN(new_n1176));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  AND3_X1   g751(.A1(new_n939), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n1177), .B1(new_n939), .B2(new_n1176), .ZN(new_n1179));
  NOR2_X1   g753(.A1(new_n1178), .A2(new_n1179), .ZN(G308));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n1176), .ZN(G225));
endmodule


