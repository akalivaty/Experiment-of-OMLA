//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n452, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1137;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT66), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(new_n458), .B(KEYINPUT70), .Z(G261));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2106), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n457), .A2(new_n449), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OR2_X1    g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT71), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT71), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G113), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2104), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(KEYINPUT72), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n477), .A2(KEYINPUT72), .ZN(new_n479));
  OAI21_X1  g054(.A(G101), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n467), .A2(new_n468), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n481), .A2(G137), .A3(new_n476), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(G160));
  AND2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G136), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT73), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT74), .B1(new_n486), .B2(new_n476), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT74), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n481), .A2(new_n491), .A3(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G124), .ZN(new_n495));
  OR2_X1    g070(.A1(G100), .A2(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n496), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  INV_X1    g074(.A(KEYINPUT75), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n476), .B2(G114), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT75), .A3(G2105), .ZN(new_n503));
  INV_X1    g078(.A(G102), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n476), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n501), .A2(new_n503), .A3(G2104), .A4(new_n505), .ZN(new_n506));
  OAI211_X1 g081(.A(G126), .B(G2105), .C1(new_n484), .C2(new_n485), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n476), .A2(G138), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT4), .B1(new_n486), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n511));
  INV_X1    g086(.A(new_n509), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n481), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n508), .B1(new_n510), .B2(new_n513), .ZN(G164));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n525), .B1(new_n526), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n520), .A2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n515), .A2(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n539));
  INV_X1    g114(.A(new_n524), .ZN(new_n540));
  INV_X1    g115(.A(G51), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n536), .B(new_n538), .C1(new_n542), .C2(KEYINPUT76), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n542), .A2(KEYINPUT76), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n543), .A2(new_n544), .ZN(G168));
  AOI22_X1  g120(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n546), .A2(new_n519), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n524), .A2(G52), .ZN(new_n548));
  INV_X1    g123(.A(G90), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n531), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n547), .A2(new_n550), .ZN(G171));
  AOI22_X1  g126(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n519), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n524), .A2(G43), .ZN(new_n554));
  INV_X1    g129(.A(G81), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n555), .B2(new_n531), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n524), .A2(G53), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G91), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n566), .A2(new_n519), .B1(new_n567), .B2(new_n531), .ZN(new_n568));
  NOR2_X1   g143(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G299));
  INV_X1    g145(.A(G171), .ZN(G301));
  OR2_X1    g146(.A1(new_n543), .A2(new_n544), .ZN(G286));
  NAND2_X1  g147(.A1(new_n537), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n524), .A2(G49), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  OAI211_X1 g151(.A(G48), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n531), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n515), .B2(new_n516), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n537), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n519), .B2(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n531), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n517), .A2(G66), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n519), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G54), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n597), .B1(new_n540), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n524), .A2(KEYINPUT77), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n590), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  OR3_X1    g181(.A1(G168), .A2(KEYINPUT78), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT78), .B1(G168), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n569), .ZN(G297));
  OAI211_X1 g184(.A(new_n607), .B(new_n608), .C1(G868), .C2(new_n569), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n603), .B1(new_n611), .B2(G860), .ZN(G148));
  NOR2_X1   g187(.A1(new_n557), .A2(G868), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n603), .A2(new_n611), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G868), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g192(.A(new_n481), .B1(new_n478), .B2(new_n479), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT13), .Z(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n487), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n476), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI221_X1 g202(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n493), .C2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G2096), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n622), .A2(new_n623), .A3(new_n630), .ZN(G156));
  INV_X1    g206(.A(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n636), .B1(new_n635), .B2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n643), .ZN(new_n645));
  AND3_X1   g220(.A1(new_n644), .A2(G14), .A3(new_n645), .ZN(G401));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n621), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n629), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n654), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1956), .B(G2474), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1961), .B(G1966), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n660), .A2(new_n663), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT20), .Z(new_n667));
  AOI211_X1 g242(.A(new_n665), .B(new_n667), .C1(new_n660), .C2(new_n664), .ZN(new_n668));
  XOR2_X1   g243(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  MUX2_X1   g249(.A(G24), .B(G290), .S(G16), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1986), .ZN(new_n676));
  MUX2_X1   g251(.A(G6), .B(G305), .S(G16), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT82), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT32), .B(G1981), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n678), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G22), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(G166), .B2(new_n683), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1971), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n683), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n683), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT33), .B(G1976), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  NOR4_X1   g266(.A1(new_n681), .A2(new_n682), .A3(new_n686), .A4(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT34), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n676), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G25), .A2(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n487), .A2(G131), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n476), .A2(G107), .ZN(new_n697));
  OAI21_X1  g272(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n698));
  INV_X1    g273(.A(G119), .ZN(new_n699));
  OAI221_X1 g274(.A(new_n696), .B1(new_n697), .B2(new_n698), .C1(new_n493), .C2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n695), .B1(new_n702), .B2(G29), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT81), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT35), .B(G1991), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n694), .B(new_n706), .C1(new_n693), .C2(new_n692), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT83), .B(KEYINPUT36), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n683), .A2(G19), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT87), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n557), .B2(new_n683), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1341), .ZN(new_n713));
  NOR2_X1   g288(.A1(G171), .A2(new_n683), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G5), .B2(new_n683), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n713), .B1(new_n717), .B2(KEYINPUT93), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G32), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n487), .A2(G141), .ZN(new_n721));
  OAI21_X1  g296(.A(G105), .B1(new_n478), .B2(new_n479), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT26), .Z(new_n724));
  NAND3_X1  g299(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G129), .B2(new_n494), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n720), .B1(new_n726), .B2(new_n719), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT89), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT27), .B(G1996), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n718), .B1(KEYINPUT93), .B2(new_n717), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT25), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n487), .A2(G139), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n735), .A2(new_n476), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n734), .A2(new_n736), .A3(new_n719), .ZN(new_n737));
  INV_X1    g312(.A(G33), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n719), .B2(new_n738), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G2072), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n715), .A2(new_n716), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(G2072), .ZN(new_n742));
  NAND2_X1  g317(.A1(G160), .A2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT24), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(KEYINPUT24), .B2(new_n744), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(G2084), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n740), .A2(new_n741), .A3(new_n742), .A4(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT31), .B(G11), .Z(new_n751));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n719), .B1(new_n752), .B2(G28), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n753), .A2(KEYINPUT92), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(new_n752), .B2(G28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n753), .A2(KEYINPUT92), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n628), .A2(new_n719), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n751), .B(new_n757), .C1(new_n758), .C2(KEYINPUT91), .ZN(new_n759));
  OAI221_X1 g334(.A(new_n759), .B1(KEYINPUT91), .B2(new_n758), .C1(new_n748), .C2(new_n747), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n719), .A2(G26), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT28), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n494), .A2(G128), .ZN(new_n763));
  OAI21_X1  g338(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n764));
  INV_X1    g339(.A(G116), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G2105), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(new_n487), .B2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT88), .B(G2067), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n683), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n683), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n771), .B1(G1966), .B2(new_n773), .ZN(new_n774));
  NOR4_X1   g349(.A1(new_n730), .A2(new_n750), .A3(new_n760), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n683), .A2(G20), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT95), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT23), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G299), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT96), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G1956), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n719), .A2(G27), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n719), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT94), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G2078), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G1966), .B2(new_n773), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n775), .A2(new_n781), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n719), .A2(G35), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G162), .B2(new_n719), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT29), .Z(new_n790));
  INV_X1    g365(.A(G2090), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G4), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT84), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n602), .B2(new_n683), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT86), .Z(new_n796));
  XOR2_X1   g371(.A(KEYINPUT85), .B(G1348), .Z(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n790), .A2(new_n791), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n798), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n792), .A2(new_n799), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n728), .A2(new_n729), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT90), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n787), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n709), .A2(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n603), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(new_n519), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n524), .A2(G55), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n813), .B2(new_n531), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n557), .A2(new_n815), .ZN(new_n816));
  OAI22_X1  g391(.A1(new_n553), .A2(new_n556), .B1(new_n811), .B2(new_n814), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n809), .B(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  INV_X1    g395(.A(G860), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n815), .A2(new_n821), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT37), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(G145));
  XNOR2_X1  g401(.A(new_n702), .B(KEYINPUT98), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(new_n619), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n702), .A2(KEYINPUT98), .ZN(new_n829));
  INV_X1    g404(.A(new_n619), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n702), .A2(KEYINPUT98), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n494), .A2(G130), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  INV_X1    g410(.A(G118), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(G2105), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n487), .B2(G142), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n833), .B(new_n839), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n734), .A2(new_n736), .A3(KEYINPUT97), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n726), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n768), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n510), .A2(new_n513), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n506), .A2(new_n507), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n843), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n628), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n498), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT100), .Z(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(new_n840), .B2(new_n847), .ZN(new_n853));
  AOI21_X1  g428(.A(G37), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n833), .A2(new_n839), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n833), .A2(new_n839), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n847), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT99), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n840), .A2(new_n859), .A3(new_n847), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n848), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n854), .B1(new_n861), .B2(new_n851), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(G395));
  OR3_X1    g439(.A1(new_n602), .A2(new_n569), .A3(KEYINPUT102), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT102), .B1(new_n602), .B2(new_n569), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(KEYINPUT103), .A3(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(G299), .B2(new_n603), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT103), .B1(new_n865), .B2(new_n866), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT41), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n614), .B(new_n818), .ZN(new_n871));
  AOI22_X1  g446(.A1(new_n865), .A2(new_n866), .B1(new_n569), .B2(new_n602), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n868), .A2(new_n869), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n875), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G303), .B(new_n688), .ZN(new_n878));
  XOR2_X1   g453(.A(G290), .B(G305), .Z(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT42), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n877), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n882), .A2(G868), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n883), .B1(G868), .B2(new_n815), .ZN(G295));
  OAI21_X1  g459(.A(new_n883), .B1(G868), .B2(new_n815), .ZN(G331));
  XNOR2_X1  g460(.A(new_n880), .B(KEYINPUT106), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n873), .B1(new_n868), .B2(new_n869), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT107), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n872), .A2(KEYINPUT107), .A3(KEYINPUT41), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G286), .A2(G301), .ZN(new_n894));
  NAND2_X1  g469(.A1(G168), .A2(G171), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n894), .A2(new_n818), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n818), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n896), .B2(new_n897), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n901), .B2(new_n896), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n876), .ZN(new_n904));
  OAI211_X1 g479(.A(KEYINPUT108), .B(new_n887), .C1(new_n900), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n899), .B2(new_n893), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n886), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n870), .A2(new_n903), .A3(new_n874), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n898), .B1(new_n868), .B2(new_n869), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n870), .A2(new_n903), .A3(new_n913), .A4(new_n874), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n911), .A2(new_n880), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G37), .ZN(new_n916));
  AND2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n909), .A2(new_n917), .A3(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT43), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n915), .A2(new_n916), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n914), .A2(new_n912), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n886), .B1(new_n921), .B2(new_n911), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT44), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n909), .A2(new_n917), .A3(new_n919), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT43), .B1(new_n920), .B2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n925), .A2(new_n930), .ZN(G397));
  INV_X1    g506(.A(G2067), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n768), .B(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n726), .B(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n702), .A2(new_n705), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n702), .A2(new_n705), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n846), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n475), .A2(new_n480), .A3(G40), .A4(new_n482), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(G290), .A2(G1986), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT48), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n946), .A2(new_n935), .ZN(new_n952));
  OR2_X1    g527(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(KEYINPUT46), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n933), .A2(new_n726), .ZN(new_n955));
  AOI22_X1  g530(.A1(new_n953), .A2(new_n954), .B1(new_n946), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  INV_X1    g532(.A(new_n937), .ZN(new_n958));
  OAI22_X1  g533(.A1(new_n958), .A2(new_n938), .B1(G2067), .B2(new_n768), .ZN(new_n959));
  AOI211_X1 g534(.A(new_n951), .B(new_n957), .C1(new_n946), .C2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n960), .B(KEYINPUT127), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT117), .ZN(new_n962));
  AOI21_X1  g537(.A(G1384), .B1(new_n844), .B2(new_n845), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT109), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n965), .B(new_n943), .C1(G164), .C2(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n945), .B1(new_n963), .B2(KEYINPUT45), .ZN(new_n968));
  AOI21_X1  g543(.A(G1971), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AND4_X1   g544(.A1(G40), .A2(new_n475), .A3(new_n480), .A4(new_n482), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT50), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n970), .B1(new_n963), .B2(new_n971), .ZN(new_n972));
  AOI211_X1 g547(.A(KEYINPUT50), .B(G1384), .C1(new_n844), .C2(new_n845), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n972), .A2(G2090), .A3(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(G8), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n970), .A2(new_n963), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n688), .A2(G1976), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(G8), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT52), .ZN(new_n982));
  XNOR2_X1  g557(.A(KEYINPUT112), .B(G1976), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n979), .A2(new_n980), .A3(G8), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G1981), .ZN(new_n987));
  OAI221_X1 g562(.A(G86), .B1(new_n528), .B2(new_n527), .C1(new_n530), .C2(new_n529), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n585), .A2(new_n987), .A3(new_n988), .A4(new_n577), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n580), .A2(KEYINPUT113), .A3(new_n987), .A4(new_n585), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n579), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n988), .A2(KEYINPUT114), .A3(new_n577), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n994), .A2(new_n585), .A3(new_n995), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n991), .A2(new_n992), .B1(new_n996), .B2(G1981), .ZN(new_n997));
  XOR2_X1   g572(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n998));
  OAI21_X1  g573(.A(KEYINPUT116), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n1000));
  INV_X1    g575(.A(new_n998), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n991), .A2(new_n992), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n517), .A2(G61), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n519), .B1(new_n1003), .B2(new_n583), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n993), .B2(new_n579), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n987), .B1(new_n1005), .B2(new_n995), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1000), .B(new_n1001), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n999), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n979), .A2(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n997), .B2(KEYINPUT49), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n986), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n978), .A2(new_n1011), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n972), .A2(G2084), .A3(new_n973), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1966), .B1(new_n968), .B2(new_n944), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(G286), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n977), .ZN(new_n1018));
  INV_X1    g593(.A(new_n974), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n969), .B2(KEYINPUT110), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  AOI211_X1 g596(.A(new_n1021), .B(G1971), .C1(new_n967), .C2(new_n968), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n1018), .C1(new_n1020), .C2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n970), .B1(new_n942), .B2(new_n943), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n964), .B2(new_n966), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1021), .B1(new_n1027), .B2(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1028), .A2(new_n1029), .A3(new_n1019), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1030), .A2(KEYINPUT111), .A3(G8), .A4(new_n1018), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1012), .B(new_n1017), .C1(new_n1025), .C2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n962), .B1(new_n1032), .B2(KEYINPUT63), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(new_n1031), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1012), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n1016), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT63), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT117), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1018), .B1(new_n1030), .B2(G8), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1011), .ZN(new_n1040));
  NOR4_X1   g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n1037), .A4(new_n1017), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1034), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1033), .A2(new_n1038), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n963), .A2(KEYINPUT45), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1044), .B1(new_n1026), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n942), .A2(KEYINPUT50), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n963), .A2(new_n971), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1047), .A2(new_n748), .A3(new_n970), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(G8), .A3(G286), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1052), .B(G8), .C1(new_n1050), .C2(G286), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT122), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(KEYINPUT51), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G286), .A2(G8), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1015), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT122), .B1(new_n1057), .B2(new_n1052), .ZN(new_n1058));
  OAI211_X1 g633(.A(KEYINPUT122), .B(G8), .C1(new_n1050), .C2(G286), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1051), .B(new_n1055), .C1(new_n1058), .C2(new_n1061), .ZN(new_n1062));
  XOR2_X1   g637(.A(G171), .B(KEYINPUT54), .Z(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n967), .A2(new_n968), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(G2078), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1047), .A2(new_n970), .A3(new_n1048), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n716), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1064), .A2(G2078), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n968), .A2(new_n944), .A3(new_n1070), .ZN(new_n1071));
  AND3_X1   g646(.A1(new_n1068), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1069), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1063), .B(new_n1066), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1068), .B(KEYINPUT124), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(new_n1063), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1034), .A2(new_n1062), .A3(new_n1035), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT125), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1012), .B1(new_n1025), .B2(new_n1031), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT125), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(new_n1062), .A4(new_n1078), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n1084));
  XNOR2_X1  g659(.A(new_n569), .B(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n972), .A2(new_n973), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n1086), .B2(G1956), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1067), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1027), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1085), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1085), .A3(new_n1093), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n942), .A2(new_n945), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1096), .A2(KEYINPUT120), .A3(new_n932), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n979), .B2(G2067), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1097), .B(new_n1099), .C1(new_n1086), .C2(G1348), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(new_n603), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1094), .B1(new_n1095), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1095), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1094), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1100), .A2(KEYINPUT60), .A3(new_n602), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1100), .B(new_n603), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1107), .B1(new_n1108), .B2(KEYINPUT60), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT58), .B(G1341), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1065), .A2(G1996), .B1(new_n1096), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n557), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT59), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1106), .A2(new_n1109), .A3(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1105), .A2(new_n1104), .A3(new_n1094), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1103), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1080), .A2(new_n1083), .A3(new_n1116), .ZN(new_n1117));
  AOI211_X1 g692(.A(G1976), .B(G288), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(new_n1002), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1034), .A2(new_n1040), .B1(new_n1009), .B2(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1121), .A2(KEYINPUT62), .A3(new_n1051), .A4(new_n1055), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1062), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1066), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1126));
  AND4_X1   g701(.A1(G171), .A2(new_n1034), .A3(new_n1035), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1043), .A2(new_n1117), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n1130));
  XNOR2_X1  g705(.A(G290), .B(G1986), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n946), .B1(new_n940), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1130), .B1(new_n1129), .B2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n961), .B1(new_n1133), .B2(new_n1134), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g710(.A1(G229), .A2(new_n464), .A3(G401), .A4(G227), .ZN(new_n1137));
  NAND3_X1  g711(.A1(new_n1137), .A2(new_n928), .A3(new_n862), .ZN(G225));
  INV_X1    g712(.A(G225), .ZN(G308));
endmodule


