//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  OR2_X1    g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G112), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G2105), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(new_n468), .B2(new_n469), .ZN(new_n482));
  AOI211_X1 g057(.A(new_n478), .B(new_n480), .C1(G124), .C2(new_n482), .ZN(G162));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(G2105), .B1(KEYINPUT64), .B2(G114), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT64), .A2(G114), .ZN(new_n486));
  OAI211_X1 g061(.A(G2104), .B(new_n484), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n463), .C2(new_n462), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(G651), .ZN(new_n497));
  AND3_X1   g072(.A1(KEYINPUT65), .A2(KEYINPUT5), .A3(G543), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT5), .B1(KEYINPUT65), .B2(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(G62), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT66), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n499), .ZN(new_n505));
  NAND3_X1  g080(.A1(KEYINPUT65), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n507), .A2(G88), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n508), .A2(G50), .A3(G543), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n509), .B(new_n510), .C1(new_n502), .C2(KEYINPUT66), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT67), .B1(new_n504), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n502), .A2(KEYINPUT66), .ZN(new_n513));
  AND2_X1   g088(.A1(new_n509), .A2(new_n510), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n513), .A2(new_n514), .A3(new_n515), .A4(new_n503), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n512), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT68), .ZN(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT7), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n508), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n507), .A2(new_n508), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI221_X1 g101(.A(new_n522), .B1(new_n523), .B2(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n520), .A2(new_n527), .ZN(G168));
  AOI22_X1  g103(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n497), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n525), .A2(new_n531), .B1(new_n532), .B2(new_n523), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n530), .A2(new_n533), .ZN(G171));
  AND2_X1   g109(.A1(new_n508), .A2(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT69), .B(G43), .Z(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n537), .B1(new_n538), .B2(new_n525), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n497), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT70), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g120(.A(KEYINPUT71), .B(KEYINPUT8), .Z(new_n546));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  OAI21_X1  g124(.A(G65), .B1(new_n498), .B2(new_n499), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G651), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT74), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT74), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n555), .A3(G651), .ZN(new_n556));
  INV_X1    g131(.A(new_n508), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n498), .A2(new_n499), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g134(.A1(new_n554), .A2(new_n556), .B1(G91), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT72), .B(KEYINPUT9), .Z(new_n562));
  NOR3_X1   g137(.A1(new_n561), .A2(KEYINPUT73), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT73), .B1(new_n561), .B2(new_n562), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n560), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  INV_X1    g146(.A(G49), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n525), .A2(new_n571), .B1(new_n572), .B2(new_n523), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n558), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(KEYINPUT75), .A3(G651), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n559), .A2(G86), .B1(new_n535), .B2(G48), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G305));
  XOR2_X1   g161(.A(KEYINPUT76), .B(G47), .Z(new_n587));
  AOI22_X1  g162(.A1(new_n559), .A2(G85), .B1(new_n535), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI211_X1 g164(.A(new_n588), .B(KEYINPUT77), .C1(new_n497), .C2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT77), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n589), .A2(new_n497), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  INV_X1    g168(.A(new_n587), .ZN(new_n594));
  OAI22_X1  g169(.A1(new_n525), .A2(new_n593), .B1(new_n594), .B2(new_n523), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n591), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n590), .A2(new_n596), .ZN(G290));
  INV_X1    g172(.A(G54), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n523), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n599), .B2(new_n523), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n558), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(G651), .ZN(new_n605));
  AOI21_X1  g180(.A(KEYINPUT10), .B1(new_n559), .B2(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  INV_X1    g182(.A(G92), .ZN(new_n608));
  NOR3_X1   g183(.A1(new_n525), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n601), .B(new_n605), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(new_n611), .B2(G171), .ZN(G284));
  OAI21_X1  g188(.A(new_n612), .B1(new_n611), .B2(G171), .ZN(G321));
  NAND2_X1  g189(.A1(G299), .A2(new_n611), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n611), .B2(G168), .ZN(G297));
  OAI21_X1  g191(.A(new_n615), .B1(new_n611), .B2(G168), .ZN(G280));
  INV_X1    g192(.A(new_n610), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR3_X1   g199(.A1(new_n464), .A2(new_n471), .A3(G2105), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT13), .Z(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n482), .A2(G123), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n633));
  INV_X1    g208(.A(G111), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G2105), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(G135), .B2(new_n470), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n638), .A2(G2096), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n628), .A2(new_n629), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(G2096), .ZN(new_n641));
  NAND4_X1  g216(.A1(new_n630), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2427), .B(G2430), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT82), .Z(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n644), .B2(new_n645), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT84), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  OAI21_X1  g239(.A(KEYINPUT17), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI22_X1  g241(.A1(new_n665), .A2(new_n666), .B1(new_n664), .B2(new_n663), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  INV_X1    g243(.A(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n664), .A3(new_n662), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n629), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT85), .B(G2096), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n684));
  XOR2_X1   g259(.A(new_n683), .B(new_n684), .Z(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT87), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n679), .A2(new_n682), .A3(new_n686), .ZN(new_n689));
  NOR3_X1   g264(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1981), .B(G1986), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(G229));
  INV_X1    g271(.A(KEYINPUT36), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G23), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n576), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT33), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(G1976), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(G1976), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n698), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n698), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G1971), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(G1971), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n709), .A2(G16), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n710), .B1(G6), .B2(G16), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT32), .B(G1981), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND4_X1  g288(.A1(new_n704), .A2(new_n707), .A3(new_n708), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT92), .B(KEYINPUT34), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n712), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n711), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n703), .B2(new_n702), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n720), .A2(new_n715), .A3(new_n707), .A4(new_n708), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n698), .A2(G24), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT91), .Z(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G290), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(G1986), .Z(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G25), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n482), .A2(G119), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT88), .ZN(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G107), .B2(new_n481), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT89), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n470), .A2(G131), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n730), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT90), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n728), .B1(new_n738), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT35), .B(G1991), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n739), .A2(new_n741), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n725), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n717), .A2(new_n721), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n697), .B1(new_n745), .B2(KEYINPUT93), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n717), .A2(new_n721), .A3(new_n748), .A4(new_n744), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G168), .A2(new_n698), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n698), .B2(G21), .ZN(new_n752));
  INV_X1    g327(.A(G1966), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AND2_X1   g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  NOR2_X1   g331(.A1(G171), .A2(new_n698), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G5), .B2(new_n698), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n754), .B(new_n755), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n726), .A2(G32), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n470), .A2(G141), .B1(G105), .B2(new_n472), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n482), .A2(G129), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT26), .Z(new_n764));
  NAND3_X1  g339(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n760), .B1(new_n766), .B2(new_n726), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT27), .B(G1996), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(G16), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n542), .B2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G34), .ZN(new_n772));
  AOI21_X1  g347(.A(G29), .B1(new_n772), .B2(KEYINPUT24), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(KEYINPUT24), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n474), .B2(new_n726), .ZN(new_n775));
  INV_X1    g350(.A(G2084), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI22_X1  g352(.A1(new_n771), .A2(G1341), .B1(new_n777), .B2(KEYINPUT99), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n758), .A2(new_n756), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n778), .B(new_n779), .C1(KEYINPUT99), .C2(new_n777), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n759), .A2(new_n769), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n726), .A2(G35), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT100), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G162), .B2(new_n726), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT29), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2090), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n726), .A2(G33), .ZN(new_n787));
  NAND2_X1  g362(.A1(G115), .A2(G2104), .ZN(new_n788));
  INV_X1    g363(.A(G127), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n464), .B2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n481), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n791), .B2(new_n790), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n794));
  NAND3_X1  g369(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n796), .A2(new_n797), .B1(G139), .B2(new_n470), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n787), .B1(new_n800), .B2(new_n726), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G2072), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n726), .A2(G26), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT28), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n470), .A2(G140), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n482), .A2(G128), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n481), .A2(G116), .ZN(new_n807));
  OAI21_X1  g382(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n805), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n804), .B1(new_n809), .B2(G29), .ZN(new_n810));
  XOR2_X1   g385(.A(KEYINPUT95), .B(G2067), .Z(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT31), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(G11), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(G11), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT30), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n816), .A2(G28), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n726), .B1(new_n816), .B2(G28), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n814), .B(new_n815), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n637), .B2(G29), .ZN(new_n820));
  INV_X1    g395(.A(new_n775), .ZN(new_n821));
  NOR2_X1   g396(.A1(G27), .A2(G29), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G164), .B2(G29), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n821), .A2(G2084), .B1(G2078), .B2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n820), .B(new_n824), .C1(G2078), .C2(new_n823), .ZN(new_n825));
  AOI211_X1 g400(.A(new_n812), .B(new_n825), .C1(G1341), .C2(new_n771), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n698), .A2(G4), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n618), .B2(new_n698), .ZN(new_n828));
  INV_X1    g403(.A(G1348), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n786), .A2(new_n802), .A3(new_n826), .A4(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT101), .B(KEYINPUT23), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n698), .A2(G20), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT102), .B(G1956), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR3_X1   g412(.A1(new_n781), .A2(new_n831), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n750), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(KEYINPUT94), .B1(new_n745), .B2(KEYINPUT36), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n749), .B2(new_n746), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n839), .A2(new_n841), .ZN(G311));
  AND2_X1   g417(.A1(new_n746), .A2(new_n749), .ZN(new_n843));
  OAI211_X1 g418(.A(new_n750), .B(new_n838), .C1(new_n843), .C2(new_n840), .ZN(G150));
  AOI22_X1  g419(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n845), .A2(new_n497), .ZN(new_n846));
  INV_X1    g421(.A(G93), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  OAI22_X1  g423(.A1(new_n525), .A2(new_n847), .B1(new_n848), .B2(new_n523), .ZN(new_n849));
  OAI21_X1  g424(.A(G860), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  AOI22_X1  g426(.A1(new_n559), .A2(G93), .B1(new_n535), .B2(G55), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(KEYINPUT103), .C1(new_n497), .C2(new_n845), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(new_n846), .B2(new_n849), .ZN(new_n855));
  OAI221_X1 g430(.A(new_n537), .B1(new_n525), .B2(new_n538), .C1(new_n540), .C2(new_n497), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n846), .A2(new_n849), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n542), .A2(KEYINPUT103), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n618), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT104), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  AOI21_X1  g442(.A(G860), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n851), .B1(new_n869), .B2(new_n870), .ZN(G145));
  XNOR2_X1  g446(.A(G162), .B(G160), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n638), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n737), .B(new_n627), .Z(new_n874));
  XNOR2_X1  g449(.A(G164), .B(new_n809), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n482), .A2(G130), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n481), .A2(G118), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G142), .B2(new_n470), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n875), .B(new_n880), .Z(new_n881));
  OR2_X1    g456(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n874), .A2(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n799), .A2(new_n765), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n766), .B(KEYINPUT106), .Z(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n799), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n882), .B2(new_n883), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n873), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n882), .A2(new_n883), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(new_n886), .ZN(new_n893));
  INV_X1    g468(.A(new_n873), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n888), .ZN(new_n895));
  INV_X1    g470(.A(G37), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n897), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g473(.A(KEYINPUT109), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n573), .B2(new_n575), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n559), .A2(G87), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n535), .A2(G49), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT109), .A4(new_n574), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(new_n709), .ZN(new_n905));
  NOR2_X1   g480(.A1(G303), .A2(G290), .ZN(new_n906));
  AND3_X1   g481(.A1(G290), .A2(new_n516), .A3(new_n512), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n904), .B(G305), .ZN(new_n909));
  NAND2_X1  g484(.A1(G303), .A2(G290), .ZN(new_n910));
  INV_X1    g485(.A(new_n512), .ZN(new_n911));
  INV_X1    g486(.A(new_n516), .ZN(new_n912));
  OAI211_X1 g487(.A(new_n596), .B(new_n590), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT42), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n860), .B(new_n621), .ZN(new_n917));
  NAND2_X1  g492(.A1(G299), .A2(new_n618), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n610), .A2(new_n560), .A3(new_n567), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT107), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n917), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n610), .A2(new_n560), .A3(KEYINPUT108), .A4(new_n567), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n918), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT41), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(G299), .B2(new_n618), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n928), .A2(new_n929), .B1(new_n919), .B2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n922), .B(new_n924), .C1(new_n917), .C2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n916), .B1(new_n932), .B2(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(KEYINPUT110), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(G868), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(G868), .B2(new_n858), .ZN(G295));
  OAI21_X1  g513(.A(new_n937), .B1(G868), .B2(new_n858), .ZN(G331));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT43), .ZN(new_n941));
  INV_X1    g516(.A(new_n527), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT68), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n519), .B(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(G171), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n520), .A2(new_n527), .B1(new_n530), .B2(new_n533), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n860), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n857), .A2(new_n859), .A3(new_n946), .A4(new_n945), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n920), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n931), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n915), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n896), .B1(new_n953), .B2(new_n915), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n941), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n950), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n928), .A2(new_n929), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n930), .A2(new_n919), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n961), .B2(new_n951), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n908), .A2(new_n914), .ZN(new_n963));
  AOI21_X1  g538(.A(G37), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n950), .A2(KEYINPUT111), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n920), .A2(new_n929), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n930), .A2(new_n926), .A3(new_n927), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n966), .A2(new_n967), .B1(new_n949), .B2(new_n948), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n950), .A2(KEYINPUT111), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n965), .B(new_n915), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n964), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n940), .B1(new_n957), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT43), .B1(new_n955), .B2(new_n956), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n964), .A2(new_n941), .A3(new_n970), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT44), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n972), .A2(new_n975), .A3(KEYINPUT112), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n957), .A2(new_n971), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT44), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n963), .B(new_n950), .C1(new_n931), .C2(new_n952), .ZN(new_n980));
  AND4_X1   g555(.A1(new_n941), .A2(new_n980), .A3(new_n970), .A4(new_n896), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n941), .B1(new_n964), .B2(new_n954), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n940), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n977), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n976), .A2(new_n984), .ZN(G397));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G164), .B2(G1384), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n493), .A2(new_n495), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n487), .A2(new_n488), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1384), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(KEYINPUT115), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n988), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT113), .B(G40), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n467), .A2(new_n473), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n992), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(KEYINPUT50), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT116), .B(G2090), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(G1384), .B1(new_n989), .B2(new_n990), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n997), .B1(new_n1002), .B2(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT45), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(G164), .B2(G1384), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G1971), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n986), .B1(new_n1001), .B2(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n512), .A2(new_n516), .A3(G8), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n512), .A2(new_n516), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n988), .B2(new_n993), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n991), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n1019));
  INV_X1    g594(.A(new_n997), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1017), .B(new_n753), .C1(new_n1018), .C2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n995), .A2(new_n776), .A3(new_n999), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1002), .A2(KEYINPUT115), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n987), .B(G1384), .C1(new_n989), .C2(new_n990), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1004), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n1003), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1017), .B1(new_n1028), .B2(new_n753), .ZN(new_n1029));
  OAI211_X1 g604(.A(G8), .B(G168), .C1(new_n1024), .C2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT63), .ZN(new_n1031));
  OAI21_X1  g606(.A(KEYINPUT50), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n997), .B1(new_n1002), .B2(new_n994), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1032), .A2(new_n1000), .A3(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n986), .B1(new_n1034), .B2(new_n1008), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1035), .B2(new_n1014), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1016), .B1(new_n1030), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G305), .A2(G1981), .ZN(new_n1038));
  INV_X1    g613(.A(G1981), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n583), .A2(new_n1039), .A3(new_n585), .A4(new_n584), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT49), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n988), .A2(new_n993), .A3(new_n1020), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1038), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n576), .A2(G1976), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1042), .A2(G8), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT52), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT117), .B(G1976), .Z(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1054), .A2(G8), .A3(new_n1042), .A4(new_n1050), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1037), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1049), .B(new_n1056), .C1(new_n1014), .C2(new_n1009), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT63), .B1(new_n1059), .B2(new_n1030), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1043), .ZN(new_n1061));
  NOR2_X1   g636(.A1(G288), .A2(G1976), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1049), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1040), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1058), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1005), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1067));
  XNOR2_X1  g642(.A(KEYINPUT56), .B(G2072), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1020), .B1(new_n998), .B2(KEYINPUT50), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n988), .A2(new_n993), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1071), .B1(new_n1072), .B2(KEYINPUT50), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT120), .B1(new_n1073), .B2(G1956), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  INV_X1    g651(.A(G1956), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1070), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n560), .A2(new_n1080), .A3(new_n567), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n559), .A2(G91), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n555), .B1(new_n552), .B2(G651), .ZN(new_n1083));
  AOI211_X1 g658(.A(KEYINPUT74), .B(new_n497), .C1(new_n550), .C2(new_n551), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT73), .ZN(new_n1086));
  INV_X1    g661(.A(new_n562), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n535), .A2(new_n1086), .A3(G53), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n566), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n564), .ZN(new_n1090));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n1085), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1081), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1090), .B2(KEYINPUT121), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT123), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT57), .B1(new_n567), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1081), .A2(new_n1098), .A3(new_n1091), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1095), .A2(new_n1096), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1096), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1079), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1348), .B1(new_n995), .B2(new_n999), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1042), .A2(G2067), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n618), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1079), .B2(new_n1106), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1102), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  INV_X1    g684(.A(G1996), .ZN(new_n1110));
  XOR2_X1   g685(.A(KEYINPUT58), .B(G1341), .Z(new_n1111));
  AOI22_X1  g686(.A1(new_n1067), .A2(new_n1110), .B1(new_n1042), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1109), .B1(new_n1112), .B2(new_n856), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1042), .A2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(G1996), .B2(new_n1006), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(KEYINPUT59), .A3(new_n542), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n995), .A2(new_n999), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n829), .ZN(new_n1118));
  OR2_X1    g693(.A1(new_n1042), .A2(G2067), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n618), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1113), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1118), .A2(new_n610), .A3(new_n1119), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1120), .B1(new_n1123), .B2(new_n1105), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1076), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1126));
  AOI211_X1 g701(.A(KEYINPUT120), .B(G1956), .C1(new_n1032), .C2(new_n1033), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1106), .B(new_n1069), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT61), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1125), .B1(new_n1102), .B2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1069), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(new_n1099), .A3(new_n1095), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1128), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1108), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1021), .B1(new_n1072), .B2(new_n1004), .ZN(new_n1135));
  OAI21_X1  g710(.A(KEYINPUT119), .B1(new_n1135), .B2(G1966), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1136), .A2(G168), .A3(new_n1023), .A4(new_n1022), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1137), .A2(new_n1138), .A3(G8), .ZN(new_n1139));
  OAI21_X1  g714(.A(G286), .B1(new_n1024), .B2(new_n1029), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(G8), .A3(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(KEYINPUT51), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n1143));
  INV_X1    g718(.A(G2078), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT53), .B1(new_n1067), .B2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1961), .B1(new_n995), .B2(new_n999), .ZN(new_n1146));
  INV_X1    g721(.A(G40), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT124), .B1(new_n474), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT124), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n467), .A2(new_n1149), .A3(new_n473), .A4(G40), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1005), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1019), .A2(KEYINPUT53), .A3(new_n1144), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NOR4_X1   g728(.A1(new_n1145), .A2(new_n1146), .A3(new_n1153), .A4(G171), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1003), .A2(new_n1144), .A3(new_n1005), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT53), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1117), .A2(new_n756), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1135), .A2(KEYINPUT53), .A3(new_n1144), .ZN(new_n1158));
  AOI21_X1  g733(.A(G301), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1143), .B1(new_n1154), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1034), .A2(new_n1008), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1014), .B1(new_n1161), .B2(G8), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1015), .A2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1157), .A2(new_n1158), .A3(G301), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1145), .A2(new_n1146), .A3(new_n1153), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1164), .B(KEYINPUT54), .C1(new_n1165), .C2(G301), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1160), .A2(new_n1163), .A3(new_n1057), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1142), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1066), .B1(new_n1134), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1141), .A2(KEYINPUT51), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT62), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1137), .A2(new_n1138), .A3(G8), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1163), .A2(new_n1057), .A3(new_n1159), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1173), .A2(KEYINPUT125), .A3(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(KEYINPUT62), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT125), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1169), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n766), .A2(new_n1110), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n809), .B(G2067), .Z(new_n1182));
  INV_X1    g757(.A(new_n765), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1181), .B(new_n1182), .C1(new_n1110), .C2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1005), .A2(new_n997), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT114), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n738), .A2(new_n741), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n737), .A2(new_n740), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1185), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G290), .B(G1986), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1191), .B1(new_n1185), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1180), .A2(new_n1193), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1185), .ZN(new_n1196));
  NOR3_X1   g771(.A1(new_n1196), .A2(G1986), .A3(G290), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT48), .Z(new_n1198));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1191), .B2(KEYINPUT127), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n809), .A2(G2067), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1196), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  OAI22_X1  g777(.A1(new_n1195), .A2(new_n1199), .B1(new_n1202), .B2(KEYINPUT126), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1202), .A2(KEYINPUT126), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1196), .B1(new_n1183), .B2(new_n1182), .ZN(new_n1205));
  OR3_X1    g780(.A1(new_n1196), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1206));
  OAI21_X1  g781(.A(KEYINPUT46), .B1(new_n1196), .B2(G1996), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1203), .A2(new_n1204), .A3(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1194), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g786(.A1(G229), .A2(new_n459), .A3(G227), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n974), .ZN(new_n1214));
  NAND4_X1  g788(.A1(new_n1213), .A2(new_n897), .A3(new_n660), .A4(new_n1214), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


