//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1297,
    new_n1298, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XOR2_X1   g0014(.A(KEYINPUT64), .B(G244), .Z(new_n215));
  INV_X1    g0015(.A(G77), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(G226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n230), .B(new_n234), .Z(G358));
  XNOR2_X1  g0035(.A(G50), .B(G68), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT67), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G97), .ZN(new_n245));
  NOR2_X1   g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G232), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n244), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n246), .B1(new_n251), .B2(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT74), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n249), .A2(new_n250), .ZN(new_n254));
  INV_X1    g0054(.A(G226), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n255), .A2(G1698), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n253), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(KEYINPUT3), .A2(G33), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  OAI211_X1 g0059(.A(new_n256), .B(new_n253), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n252), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT75), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT75), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n252), .B(new_n264), .C1(new_n257), .C2(new_n261), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(G1), .A3(G13), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(new_n267), .A3(G274), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n267), .A2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(KEYINPUT76), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT76), .ZN(new_n277));
  OAI21_X1  g0077(.A(G238), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n273), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT13), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT13), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n269), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n282), .A2(G190), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n267), .B1(new_n262), .B2(KEYINPUT75), .ZN(new_n286));
  AOI211_X1 g0086(.A(KEYINPUT13), .B(new_n279), .C1(new_n286), .C2(new_n265), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n283), .B1(new_n269), .B2(new_n280), .ZN(new_n288));
  OAI21_X1  g0088(.A(G200), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G20), .A2(G33), .ZN(new_n290));
  INV_X1    g0090(.A(G68), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(G50), .B1(G20), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n212), .A2(G33), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT69), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n294), .B2(new_n216), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n211), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n295), .A2(KEYINPUT11), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n291), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n301), .B(KEYINPUT12), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(new_n297), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n270), .A2(G20), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n303), .A2(G68), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n298), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT11), .B1(new_n295), .B2(new_n297), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n285), .A2(new_n289), .A3(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT77), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n285), .A2(new_n289), .A3(KEYINPUT77), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n270), .B2(G20), .ZN(new_n315));
  AOI22_X1  g0115(.A1(new_n315), .A2(new_n303), .B1(new_n300), .B2(new_n314), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT16), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT7), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n254), .B2(G20), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n259), .A2(new_n258), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n291), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g0123(.A1(G58), .A2(G68), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n201), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n290), .A2(G159), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n318), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT7), .B1(new_n321), .B2(new_n212), .ZN(new_n329));
  NOR4_X1   g0129(.A1(new_n259), .A2(new_n258), .A3(new_n319), .A4(G20), .ZN(new_n330));
  OAI21_X1  g0130(.A(G68), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n327), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(KEYINPUT16), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n297), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT78), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT78), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n328), .A2(new_n333), .A3(new_n336), .A4(new_n297), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n317), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT80), .ZN(new_n339));
  INV_X1    g0139(.A(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(G223), .B(new_n340), .C1(new_n259), .C2(new_n258), .ZN(new_n341));
  OAI211_X1 g0141(.A(G226), .B(G1698), .C1(new_n259), .C2(new_n258), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G87), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n344), .A2(KEYINPUT79), .A3(new_n268), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT79), .B1(new_n344), .B2(new_n268), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n267), .A2(G232), .A3(new_n271), .ZN(new_n347));
  AND2_X1   g0147(.A1(KEYINPUT71), .A2(G179), .ZN(new_n348));
  NOR2_X1   g0148(.A1(KEYINPUT71), .A2(G179), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n273), .A2(new_n347), .A3(new_n350), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n345), .A2(new_n346), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n344), .A2(new_n268), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n273), .A2(new_n347), .ZN(new_n354));
  AOI21_X1  g0154(.A(G169), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n339), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT79), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n344), .A2(KEYINPUT79), .A3(new_n268), .ZN(new_n359));
  INV_X1    g0159(.A(new_n351), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n353), .A2(new_n354), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n361), .A2(KEYINPUT80), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT18), .B1(new_n338), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n297), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n331), .A2(new_n332), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(new_n318), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n336), .B1(new_n370), .B2(new_n333), .ZN(new_n371));
  AND4_X1   g0171(.A1(new_n336), .A2(new_n328), .A3(new_n297), .A4(new_n333), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n316), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n361), .A2(KEYINPUT80), .A3(new_n364), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT80), .B1(new_n361), .B2(new_n364), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n367), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n358), .A2(new_n380), .A3(new_n359), .A4(new_n354), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n362), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n316), .B(new_n384), .C1(new_n371), .C2(new_n372), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT17), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n338), .A2(KEYINPUT17), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n313), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT14), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(G169), .C1(new_n287), .C2(new_n288), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n282), .A2(G179), .A3(new_n284), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n282), .A2(new_n284), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n396), .B2(G169), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n395), .A2(new_n397), .B1(new_n307), .B2(new_n306), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G50), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n212), .B1(new_n201), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT70), .ZN(new_n402));
  XNOR2_X1  g0202(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(G150), .ZN(new_n404));
  INV_X1    g0204(.A(new_n290), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n403), .B1(new_n404), .B2(new_n405), .C1(new_n294), .C2(new_n314), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n297), .ZN(new_n407));
  INV_X1    g0207(.A(new_n303), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n304), .A2(G50), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n408), .A2(new_n409), .B1(G50), .B2(new_n299), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT9), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n254), .A2(G222), .A3(new_n340), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n216), .B2(new_n254), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n254), .A2(G1698), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT68), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n418), .B2(G223), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n419), .A2(new_n267), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n273), .B1(new_n255), .B2(new_n274), .ZN(new_n421));
  OAI21_X1  g0221(.A(G200), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n421), .ZN(new_n423));
  OAI211_X1 g0223(.A(G190), .B(new_n423), .C1(new_n419), .C2(new_n267), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n407), .A2(KEYINPUT9), .A3(new_n411), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n414), .A2(new_n422), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT10), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT9), .B1(new_n407), .B2(new_n411), .ZN(new_n428));
  AOI211_X1 g0228(.A(new_n413), .B(new_n410), .C1(new_n406), .C2(new_n297), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT10), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n424), .A4(new_n422), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n420), .A2(new_n421), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n350), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n412), .C1(G169), .C2(new_n434), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n215), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n267), .A2(G274), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n438), .A2(new_n275), .B1(new_n439), .B2(new_n272), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n251), .A2(new_n340), .ZN(new_n441));
  XNOR2_X1  g0241(.A(KEYINPUT72), .B(G107), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n441), .B1(new_n254), .B2(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n418), .B2(G238), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n440), .B1(new_n444), .B2(new_n267), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G200), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n303), .A2(G77), .A3(new_n304), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G77), .B2(new_n299), .ZN(new_n448));
  INV_X1    g0248(.A(new_n314), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n449), .A2(new_n290), .B1(G20), .B2(G77), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT15), .B(G87), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT73), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(new_n293), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n448), .B1(new_n453), .B2(new_n297), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n446), .B(new_n454), .C1(new_n380), .C2(new_n445), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n454), .B1(new_n445), .B2(new_n363), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n350), .B(new_n440), .C1(new_n444), .C2(new_n267), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(new_n458), .ZN(new_n459));
  NOR4_X1   g0259(.A1(new_n391), .A2(new_n399), .A3(new_n437), .A4(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(G107), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT72), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT72), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G107), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT23), .B1(new_n465), .B2(new_n212), .ZN(new_n466));
  INV_X1    g0266(.A(G116), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT84), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G116), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(new_n212), .A3(G33), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n212), .A2(G107), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT23), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n466), .A2(new_n472), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n254), .A2(new_n212), .A3(G87), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT22), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n479), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n254), .A2(new_n481), .A3(new_n212), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT24), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n476), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n476), .B2(new_n483), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n297), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(G13), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G1), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n473), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT25), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n270), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n299), .A2(new_n493), .A3(new_n211), .A4(new_n296), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n461), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(G257), .B(G1698), .C1(new_n259), .C2(new_n258), .ZN(new_n497));
  OAI211_X1 g0297(.A(G250), .B(new_n340), .C1(new_n259), .C2(new_n258), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n268), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n270), .A2(G45), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g0303(.A(G41), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT5), .A2(G41), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(new_n268), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G264), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(G274), .A3(new_n267), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n501), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n268), .A2(new_n500), .B1(new_n508), .B2(G264), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT87), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n510), .ZN(new_n515));
  AOI21_X1  g0315(.A(G190), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(G200), .B1(new_n513), .B2(new_n510), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n488), .B(new_n496), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n512), .A2(new_n515), .A3(G169), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n501), .A2(new_n509), .A3(G179), .A4(new_n510), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT88), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT88), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n513), .A2(new_n523), .A3(G179), .A4(new_n510), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n520), .A2(new_n525), .B1(new_n488), .B2(new_n496), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(G20), .B1(new_n246), .B2(KEYINPUT19), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT85), .ZN(new_n529));
  INV_X1    g0329(.A(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n245), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n529), .B1(new_n465), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n442), .A2(KEYINPUT85), .A3(new_n530), .A4(new_n245), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n254), .A2(new_n212), .A3(G68), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n293), .A2(new_n245), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(KEYINPUT19), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n297), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n452), .A2(new_n300), .ZN(new_n539));
  INV_X1    g0339(.A(new_n494), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G87), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n267), .A2(G250), .A3(new_n502), .ZN(new_n543));
  INV_X1    g0343(.A(G45), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G1), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n267), .A2(G274), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(G244), .B(G1698), .C1(new_n259), .C2(new_n258), .ZN(new_n548));
  OAI211_X1 g0348(.A(G238), .B(new_n340), .C1(new_n259), .C2(new_n258), .ZN(new_n549));
  XNOR2_X1  g0349(.A(KEYINPUT84), .B(G116), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n548), .B(new_n549), .C1(new_n244), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n547), .B1(new_n551), .B2(new_n268), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n380), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G200), .B2(new_n552), .ZN(new_n554));
  INV_X1    g0354(.A(new_n350), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n555), .B(new_n547), .C1(new_n268), .C2(new_n551), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n268), .ZN(new_n557));
  INV_X1    g0357(.A(new_n547), .ZN(new_n558));
  AOI21_X1  g0358(.A(G169), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n452), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n540), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n538), .A2(new_n539), .A3(new_n562), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n542), .A2(new_n554), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G250), .A2(G1698), .ZN(new_n566));
  NAND2_X1  g0366(.A1(KEYINPUT4), .A2(G244), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(G1698), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n254), .A2(new_n568), .B1(G33), .B2(G283), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(new_n340), .C1(new_n259), .C2(new_n258), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n268), .ZN(new_n574));
  INV_X1    g0374(.A(new_n506), .ZN(new_n575));
  NOR2_X1   g0375(.A1(KEYINPUT5), .A2(G41), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n545), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(G257), .A3(new_n267), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n510), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n579), .A3(new_n350), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n267), .B1(new_n569), .B2(new_n572), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n510), .A2(new_n578), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n363), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n299), .A2(G97), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n585), .B1(new_n540), .B2(G97), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n465), .B1(new_n329), .B2(new_n330), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n245), .A2(new_n461), .A3(KEYINPUT6), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT6), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G97), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n461), .A2(KEYINPUT81), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G107), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n589), .A2(new_n591), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n589), .A2(new_n591), .B1(new_n592), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g0396(.A(G20), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n290), .A2(G77), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n588), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n587), .B1(new_n599), .B2(new_n297), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n565), .B1(new_n584), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n297), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n586), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n603), .A2(KEYINPUT83), .A3(new_n580), .A4(new_n583), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n574), .A2(new_n579), .A3(KEYINPUT82), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT82), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n581), .B2(new_n582), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n605), .A2(new_n607), .A3(G200), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n574), .A2(new_n579), .A3(G190), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n600), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n564), .A2(new_n601), .A3(new_n604), .A4(new_n610), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n508), .A2(G270), .B1(new_n439), .B2(new_n507), .ZN(new_n612));
  OAI211_X1 g0412(.A(G264), .B(G1698), .C1(new_n259), .C2(new_n258), .ZN(new_n613));
  OAI211_X1 g0413(.A(G257), .B(new_n340), .C1(new_n259), .C2(new_n258), .ZN(new_n614));
  INV_X1    g0414(.A(G303), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n254), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n268), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  OAI22_X1  g0418(.A1(new_n494), .A2(new_n467), .B1(new_n299), .B2(new_n471), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G33), .A2(G283), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n621), .B(new_n212), .C1(G33), .C2(new_n245), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n297), .B(new_n622), .C1(new_n471), .C2(new_n212), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT20), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n620), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n618), .A2(G179), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n363), .B1(new_n612), .B2(new_n617), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(new_n627), .A3(KEYINPUT21), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT21), .B1(new_n629), .B2(new_n627), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n612), .A2(new_n617), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n627), .B1(G200), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n380), .B2(new_n634), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n611), .A2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n460), .A2(new_n527), .A3(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n436), .ZN(new_n640));
  INV_X1    g0440(.A(new_n379), .ZN(new_n641));
  INV_X1    g0441(.A(new_n458), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n399), .B1(new_n642), .B2(new_n309), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n641), .B1(new_n643), .B2(new_n389), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n640), .B1(new_n644), .B2(new_n433), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n512), .A2(new_n515), .A3(G169), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n522), .A2(new_n524), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n476), .A2(new_n483), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(KEYINPUT24), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n368), .B1(new_n649), .B2(new_n485), .ZN(new_n650));
  INV_X1    g0450(.A(new_n496), .ZN(new_n651));
  OAI22_X1  g0451(.A1(new_n646), .A2(new_n647), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(KEYINPUT89), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT89), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n525), .A2(new_n520), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n488), .A2(new_n496), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n633), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n611), .A2(new_n519), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT26), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n604), .A2(new_n601), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n662), .B2(new_n564), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n560), .A2(new_n563), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n542), .A2(new_n554), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n584), .A2(new_n600), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n664), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n664), .B1(new_n667), .B2(KEYINPUT26), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n660), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n460), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n645), .A2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n490), .A2(new_n212), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT90), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT27), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n673), .B(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n675), .A2(new_n679), .A3(G213), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n656), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n527), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT92), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT92), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n527), .A2(new_n686), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n526), .A2(new_n682), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n629), .A2(new_n627), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT21), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n628), .A3(new_n630), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n682), .A2(new_n627), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n637), .B2(new_n696), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  XOR2_X1   g0499(.A(KEYINPUT91), .B(G330), .Z(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n633), .A2(new_n682), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n685), .A2(new_n687), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n653), .A2(new_n657), .A3(new_n682), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n707), .B1(new_n706), .B2(new_n708), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n704), .B1(new_n710), .B2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(KEYINPUT94), .ZN(new_n713));
  INV_X1    g0513(.A(new_n206), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(G41), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n206), .A2(KEYINPUT94), .A3(new_n504), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G1), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n532), .A2(new_n533), .A3(new_n467), .ZN(new_n719));
  OAI22_X1  g0519(.A1(new_n718), .A2(new_n719), .B1(new_n209), .B2(new_n717), .ZN(new_n720));
  XOR2_X1   g0520(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n721));
  XNOR2_X1  g0521(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XOR2_X1   g0522(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n680), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G343), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n724), .B1(new_n670), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n695), .B1(new_n656), .B2(new_n655), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n728), .A2(new_n611), .A3(new_n519), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT98), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n560), .A2(new_n731), .A3(new_n563), .ZN(new_n732));
  AOI22_X1  g0532(.A1(new_n667), .A2(KEYINPUT26), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n662), .A2(new_n661), .A3(new_n564), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n726), .B1(new_n729), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT99), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n652), .A2(new_n633), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n604), .A2(new_n601), .A3(new_n610), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n738), .A2(new_n739), .A3(new_n518), .A4(new_n564), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(new_n734), .A3(new_n733), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT99), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n742), .A3(new_n726), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n727), .B1(new_n744), .B2(KEYINPUT29), .ZN(new_n745));
  XOR2_X1   g0545(.A(KEYINPUT96), .B(KEYINPUT31), .Z(new_n746));
  INV_X1    g0546(.A(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n618), .A2(G179), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n513), .A2(new_n552), .A3(new_n574), .A4(new_n579), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n574), .A2(new_n579), .ZN(new_n751));
  INV_X1    g0551(.A(new_n552), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G179), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n634), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n753), .A2(new_n755), .A3(KEYINPUT30), .A4(new_n513), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n555), .B1(new_n612), .B2(new_n617), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n757), .A2(new_n511), .A3(new_n751), .A4(new_n752), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n750), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n682), .ZN(new_n760));
  MUX2_X1   g0560(.A(new_n746), .B(KEYINPUT31), .S(new_n760), .Z(new_n761));
  NAND3_X1  g0561(.A1(new_n638), .A2(new_n527), .A3(new_n726), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n700), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n745), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n722), .B1(new_n764), .B2(G1), .ZN(G364));
  NOR2_X1   g0565(.A1(G13), .A2(G33), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT101), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n699), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n717), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n489), .A2(G20), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G45), .ZN(new_n772));
  OR2_X1    g0572(.A1(new_n772), .A2(KEYINPUT100), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n270), .B1(new_n772), .B2(KEYINPUT100), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n714), .A2(new_n321), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G355), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n778), .B1(G116), .B2(new_n206), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n239), .A2(G45), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n714), .A2(new_n254), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(new_n544), .B2(new_n210), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n779), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n211), .B1(G20), .B2(new_n363), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n768), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n776), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n212), .A2(G190), .ZN(new_n789));
  NAND3_X1  g0589(.A1(new_n789), .A2(new_n754), .A3(G200), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT102), .ZN(new_n791));
  NOR2_X1   g0591(.A1(G179), .A2(G200), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT103), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n791), .A2(G283), .B1(new_n794), .B2(G329), .ZN(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT104), .Z(new_n796));
  NAND3_X1  g0596(.A1(new_n555), .A2(new_n382), .A3(new_n789), .ZN(new_n797));
  INV_X1    g0597(.A(G311), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n212), .A2(new_n380), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n800), .A2(new_n754), .A3(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n792), .A2(G190), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI221_X1 g0605(.A(new_n321), .B1(new_n801), .B2(new_n615), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n212), .A2(new_n382), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n555), .A2(G190), .A3(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G326), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n555), .A2(new_n382), .A3(new_n800), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n555), .A2(new_n380), .A3(new_n807), .ZN(new_n813));
  XNOR2_X1  g0613(.A(KEYINPUT105), .B(KEYINPUT33), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(G317), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n810), .B1(new_n811), .B2(new_n812), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  NOR4_X1   g0616(.A1(new_n796), .A2(new_n799), .A3(new_n806), .A4(new_n816), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(KEYINPUT106), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(KEYINPUT106), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n254), .B1(new_n801), .B2(new_n530), .ZN(new_n820));
  INV_X1    g0620(.A(new_n793), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(G159), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT32), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n820), .B(new_n823), .C1(G97), .C2(new_n803), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n791), .A2(G107), .ZN(new_n825));
  INV_X1    g0625(.A(new_n812), .ZN(new_n826));
  INV_X1    g0626(.A(new_n797), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G58), .A2(new_n826), .B1(new_n827), .B2(G77), .ZN(new_n828));
  INV_X1    g0628(.A(new_n813), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G50), .A2(new_n809), .B1(new_n829), .B2(G68), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n824), .A2(new_n825), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n818), .A2(new_n819), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n788), .B1(new_n832), .B2(new_n785), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n701), .A2(new_n776), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n699), .A2(new_n700), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n769), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G396));
  NAND2_X1  g0637(.A1(new_n670), .A2(new_n726), .ZN(new_n838));
  INV_X1    g0638(.A(new_n446), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n454), .B1(new_n445), .B2(new_n380), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n839), .A2(new_n840), .B1(new_n454), .B2(new_n726), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n458), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n642), .A2(new_n726), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n682), .B1(new_n660), .B2(new_n669), .ZN(new_n846));
  INV_X1    g0646(.A(new_n844), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n763), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT107), .Z(new_n852));
  AOI21_X1  g0652(.A(new_n776), .B1(new_n849), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n776), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n785), .A2(new_n766), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n216), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n785), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n791), .A2(G87), .ZN(new_n859));
  INV_X1    g0659(.A(new_n794), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n859), .B1(new_n805), .B2(new_n812), .C1(new_n798), .C2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(G283), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n813), .A2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n321), .B1(new_n801), .B2(new_n461), .C1(new_n804), .C2(new_n245), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n615), .A2(new_n808), .B1(new_n797), .B2(new_n550), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n861), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G137), .A2(new_n809), .B1(new_n829), .B2(G150), .ZN(new_n867));
  INV_X1    g0667(.A(G143), .ZN(new_n868));
  INV_X1    g0668(.A(G159), .ZN(new_n869));
  OAI221_X1 g0669(.A(new_n867), .B1(new_n868), .B2(new_n812), .C1(new_n869), .C2(new_n797), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT34), .ZN(new_n871));
  OR2_X1    g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n791), .A2(G68), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n254), .B1(new_n801), .B2(new_n400), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(G58), .B2(new_n803), .ZN(new_n875));
  INV_X1    g0675(.A(G132), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n873), .B(new_n875), .C1(new_n876), .C2(new_n860), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n870), .B2(new_n871), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n866), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n857), .B1(new_n858), .B2(new_n879), .C1(new_n847), .C2(new_n767), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n854), .A2(new_n880), .ZN(G384));
  NOR2_X1   g0681(.A1(new_n771), .A2(new_n270), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n682), .B1(new_n307), .B2(new_n306), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT109), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n884), .A2(new_n309), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n398), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(G169), .B1(new_n287), .B2(new_n288), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT14), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(new_n394), .A3(new_n393), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n311), .B2(new_n312), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n886), .B1(new_n890), .B2(new_n883), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n334), .A2(new_n316), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n725), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n379), .B2(new_n389), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n356), .A2(new_n365), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n385), .A2(new_n896), .A3(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(KEYINPUT37), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT110), .B1(new_n338), .B2(new_n366), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT110), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n373), .A2(new_n376), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(KEYINPUT111), .B(KEYINPUT37), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n385), .B(new_n903), .C1(new_n338), .C2(new_n680), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n898), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n895), .A2(new_n905), .A3(KEYINPUT38), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n895), .B2(new_n905), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n682), .B(new_n844), .C1(new_n660), .C2(new_n669), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n843), .B(KEYINPUT108), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n891), .B1(new_n906), .B2(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  INV_X1    g0711(.A(new_n903), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n385), .B1(new_n366), .B2(new_n338), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n338), .A2(new_n680), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n912), .B1(new_n338), .B2(new_n384), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n373), .A2(new_n725), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n916), .A2(new_n899), .A3(new_n901), .A4(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n914), .B1(new_n379), .B2(new_n389), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n911), .B1(new_n906), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n895), .A2(new_n905), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT38), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n895), .A2(new_n905), .A3(KEYINPUT38), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n399), .A2(new_n726), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n922), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n641), .A2(new_n725), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n910), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT112), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT112), .ZN(new_n935));
  NAND4_X1  g0735(.A1(new_n910), .A2(new_n930), .A3(new_n935), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n745), .A2(KEYINPUT113), .A3(new_n460), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n733), .A2(new_n734), .ZN(new_n939));
  AOI211_X1 g0739(.A(KEYINPUT99), .B(new_n682), .C1(new_n939), .C2(new_n740), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n742), .B1(new_n741), .B2(new_n726), .ZN(new_n941));
  OAI21_X1  g0741(.A(KEYINPUT29), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n838), .A2(new_n723), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n942), .A2(new_n460), .A3(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT113), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n938), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n645), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n937), .B(new_n948), .Z(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n906), .A2(new_n907), .ZN(new_n951));
  INV_X1    g0751(.A(new_n746), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(new_n759), .B2(new_n682), .ZN(new_n953));
  INV_X1    g0753(.A(new_n760), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(KEYINPUT31), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n844), .B1(new_n762), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n889), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n883), .B1(new_n313), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n398), .A2(new_n885), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n950), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT114), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n891), .B(new_n956), .C1(new_n906), .C2(new_n907), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n964), .A2(KEYINPUT114), .A3(new_n950), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n956), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n921), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n926), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n966), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n762), .A2(new_n955), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n460), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n700), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n972), .B2(new_n974), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n882), .B1(new_n949), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n949), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n595), .A2(new_n596), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT35), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(KEYINPUT35), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n981), .A2(G116), .A3(new_n213), .A4(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT36), .ZN(new_n984));
  NOR3_X1   g0784(.A1(new_n209), .A2(new_n216), .A3(new_n324), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n291), .A2(G50), .ZN(new_n986));
  OAI211_X1 g0786(.A(G1), .B(new_n489), .C1(new_n985), .C2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n978), .A2(new_n984), .A3(new_n987), .ZN(G367));
  NOR2_X1   g0788(.A1(new_n234), .A2(new_n782), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n786), .B1(new_n206), .B2(new_n452), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n776), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(KEYINPUT46), .A2(G116), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n801), .A2(new_n992), .B1(new_n790), .B2(new_n245), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n254), .B(new_n993), .C1(G317), .C2(new_n821), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n801), .A2(new_n550), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n994), .B1(KEYINPUT46), .B2(new_n995), .C1(new_n442), .C2(new_n804), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G294), .A2(new_n829), .B1(new_n809), .B2(G311), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n862), .B2(new_n797), .C1(new_n615), .C2(new_n812), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G150), .A2(new_n826), .B1(new_n829), .B2(G159), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n400), .B2(new_n797), .C1(new_n868), .C2(new_n808), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n804), .A2(new_n291), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n801), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n790), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G58), .A2(new_n1003), .B1(new_n1004), .B2(G77), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n321), .B1(new_n821), .B2(G137), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI22_X1  g0807(.A1(new_n996), .A2(new_n998), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT47), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n991), .B1(new_n1009), .B2(new_n785), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n564), .B1(new_n542), .B2(new_n726), .ZN(new_n1011));
  OR3_X1    g0811(.A1(new_n664), .A2(new_n542), .A3(new_n726), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1011), .A2(new_n1012), .A3(new_n768), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n739), .B1(new_n600), .B2(new_n726), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n666), .A2(new_n682), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n710), .B2(new_n711), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT45), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g0820(.A(KEYINPUT45), .B(new_n1017), .C1(new_n710), .C2(new_n711), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n711), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1017), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1023), .A2(new_n709), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT44), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(KEYINPUT44), .A3(new_n709), .A4(new_n1024), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1022), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n703), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n1020), .A2(new_n1021), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n704), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n706), .B1(new_n690), .B2(new_n705), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(new_n701), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n764), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1031), .A2(new_n1033), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n764), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n717), .B(KEYINPUT41), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n775), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1043));
  AOI21_X1  g0843(.A(KEYINPUT43), .B1(new_n1043), .B2(KEYINPUT115), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(KEYINPUT115), .B2(new_n1043), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(KEYINPUT43), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT42), .ZN(new_n1048));
  OR3_X1    g0848(.A1(new_n706), .A2(new_n1048), .A3(new_n1024), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1048), .B1(new_n706), .B2(new_n1024), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n601), .B(new_n604), .C1(new_n1024), .C2(new_n652), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1049), .A2(new_n1050), .B1(new_n726), .B2(new_n1051), .ZN(new_n1052));
  MUX2_X1   g0852(.A(new_n1047), .B(new_n1045), .S(new_n1052), .Z(new_n1053));
  NOR2_X1   g0853(.A1(new_n704), .A2(new_n1024), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1014), .B1(new_n1042), .B2(new_n1055), .ZN(G387));
  NAND2_X1  g0856(.A1(new_n1035), .A2(new_n775), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1003), .A2(G77), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n254), .C1(new_n404), .C2(new_n793), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G50), .B2(new_n826), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n291), .A2(new_n797), .B1(new_n808), .B2(new_n869), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n449), .B2(new_n829), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n791), .A2(G97), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n561), .A2(new_n803), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1060), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n254), .B1(new_n821), .B2(G326), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n804), .A2(new_n862), .B1(new_n801), .B2(new_n805), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(G311), .A2(new_n829), .B1(new_n809), .B2(G322), .ZN(new_n1068));
  INV_X1    g0868(.A(G317), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1068), .B1(new_n615), .B2(new_n797), .C1(new_n1069), .C2(new_n812), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1067), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT49), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1066), .B1(new_n550), .B2(new_n790), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1065), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n785), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n782), .B1(new_n230), .B2(G45), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n719), .B2(new_n777), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n314), .A2(G50), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT50), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n544), .B1(new_n291), .B2(new_n216), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n719), .B(new_n1083), .C1(new_n1082), .C2(new_n1081), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n1080), .A2(new_n1084), .B1(G107), .B2(new_n206), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n855), .B1(new_n1085), .B2(new_n786), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n768), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1078), .B(new_n1086), .C1(new_n690), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1036), .A2(new_n770), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1035), .A2(new_n764), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1057), .B(new_n1088), .C1(new_n1089), .C2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1024), .A2(new_n768), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n786), .B1(new_n245), .B2(new_n206), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n242), .B2(new_n781), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n404), .A2(new_n808), .B1(new_n812), .B2(new_n869), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT51), .Z(new_n1097));
  AOI22_X1  g0897(.A1(new_n1003), .A2(G68), .B1(new_n821), .B2(G143), .ZN(new_n1098));
  INV_X1    g0898(.A(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1099), .A2(KEYINPUT117), .B1(new_n829), .B2(G50), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n321), .B1(new_n803), .B2(G77), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n1098), .A2(new_n1102), .B1(new_n827), .B2(new_n449), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1100), .A2(new_n859), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n798), .A2(new_n812), .B1(new_n808), .B2(new_n1069), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT52), .Z(new_n1106));
  OAI221_X1 g0906(.A(new_n321), .B1(new_n793), .B2(new_n811), .C1(new_n801), .C2(new_n862), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(new_n471), .B2(new_n803), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n829), .A2(G303), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n827), .A2(G294), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1108), .A2(new_n825), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n1097), .A2(new_n1104), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n855), .B(new_n1095), .C1(new_n1112), .C2(new_n785), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1093), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT116), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT116), .B1(new_n1032), .B2(new_n704), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n775), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1114), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1038), .A2(new_n770), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(new_n1119), .B2(new_n1036), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1092), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1117), .B1(new_n1115), .B2(KEYINPUT116), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n770), .B(new_n1038), .C1(new_n1125), .C2(new_n1037), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1125), .A2(new_n775), .B1(new_n1093), .B2(new_n1113), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(KEYINPUT118), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(G390));
  NAND3_X1  g0929(.A1(new_n460), .A2(G330), .A3(new_n973), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT113), .B1(new_n745), .B2(new_n460), .ZN(new_n1131));
  AND4_X1   g0931(.A1(KEYINPUT113), .A2(new_n942), .A3(new_n460), .A4(new_n943), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n645), .B(new_n1130), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n909), .B1(new_n744), .B2(new_n847), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n763), .A2(new_n847), .A3(new_n891), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n891), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n956), .A2(G330), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1135), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n891), .B1(new_n763), .B2(new_n847), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1140), .A2(new_n1141), .B1(new_n908), .B2(new_n909), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(KEYINPUT120), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n928), .B1(new_n906), .B2(new_n921), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n909), .B1(new_n846), .B2(new_n847), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n928), .B1(new_n1149), .B2(new_n1136), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n922), .A2(new_n927), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1140), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT119), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1148), .A2(new_n1152), .A3(new_n1135), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n847), .B1(new_n940), .B2(new_n941), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n909), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1146), .B1(new_n1160), .B2(new_n891), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n891), .B1(new_n908), .B2(new_n909), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n1162), .A2(new_n928), .B1(new_n922), .B2(new_n927), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1157), .B(new_n1140), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1155), .A2(new_n1156), .A3(new_n1164), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1145), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1164), .A2(new_n1156), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1157), .B1(new_n1153), .B2(new_n1140), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n717), .B1(new_n1172), .B2(new_n1166), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n775), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n855), .B1(new_n314), .B2(new_n856), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n467), .A2(new_n812), .B1(new_n808), .B2(new_n862), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G97), .B2(new_n827), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n321), .B1(new_n801), .B2(new_n530), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G77), .B2(new_n803), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n465), .A2(new_n829), .B1(new_n794), .B2(G294), .ZN(new_n1181));
  AND4_X1   g0981(.A1(new_n873), .A2(new_n1178), .A3(new_n1180), .A4(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT54), .B(G143), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n827), .A2(new_n1184), .B1(G159), .B2(new_n803), .ZN(new_n1185));
  INV_X1    g0985(.A(G137), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1185), .B1(new_n1186), .B2(new_n813), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT121), .Z(new_n1188));
  NOR2_X1   g0988(.A1(new_n801), .A2(new_n404), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT53), .ZN(new_n1190));
  INV_X1    g0990(.A(G128), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1190), .B1(new_n1191), .B2(new_n808), .C1(new_n876), .C2(new_n812), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n794), .A2(G125), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n254), .C1(new_n400), .C2(new_n790), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1182), .B1(new_n1188), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1151), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1176), .B1(new_n858), .B2(new_n1196), .C1(new_n1197), .C2(new_n767), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1174), .A2(new_n1175), .A3(new_n1198), .ZN(G378));
  AOI21_X1  g0999(.A(new_n680), .B1(new_n407), .B2(new_n411), .ZN(new_n1200));
  AND2_X1   g1000(.A1(new_n437), .A2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n437), .A2(new_n1200), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OR3_X1    g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1204), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(G330), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n968), .B2(new_n970), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1207), .B1(new_n966), .B2(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n964), .A2(KEYINPUT114), .A3(new_n950), .ZN(new_n1211));
  AOI21_X1  g1011(.A(KEYINPUT114), .B1(new_n964), .B2(new_n950), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1209), .B(new_n1207), .C1(new_n1211), .C2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n937), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1209), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1207), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1218), .A2(new_n936), .A3(new_n934), .A4(new_n1213), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1215), .A2(KEYINPUT122), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT122), .B1(new_n1215), .B2(new_n1219), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n775), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n855), .B1(new_n400), .B2(new_n856), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n804), .A2(new_n404), .B1(new_n1183), .B2(new_n801), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G125), .A2(new_n809), .B1(new_n826), .B2(G128), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1186), .B2(new_n797), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G132), .C2(new_n829), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n244), .B(new_n504), .C1(new_n790), .C2(new_n869), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G124), .B2(new_n821), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1229), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n860), .A2(new_n862), .B1(new_n467), .B2(new_n808), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1004), .A2(G58), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n254), .A2(G41), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1002), .A2(new_n1058), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n452), .A2(new_n797), .ZN(new_n1238));
  OAI22_X1  g1038(.A1(new_n245), .A2(new_n813), .B1(new_n812), .B2(new_n461), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1234), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n1240), .A2(KEYINPUT58), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G50), .B(new_n1236), .C1(new_n244), .C2(new_n504), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1240), .A2(KEYINPUT58), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(new_n1233), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1223), .B1(new_n858), .B2(new_n1244), .C1(new_n1207), .C2(new_n767), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1222), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT123), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1133), .A2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n947), .A2(KEYINPUT123), .A3(new_n645), .A4(new_n1130), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1172), .B2(new_n1166), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT122), .ZN(new_n1252));
  NOR3_X1   g1052(.A1(new_n937), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1218), .A2(new_n1213), .B1(new_n936), .B2(new_n934), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1215), .A2(KEYINPUT122), .A3(new_n1219), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1251), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n770), .B1(new_n1257), .B2(KEYINPUT57), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1248), .B(new_n1249), .C1(new_n1165), .C2(new_n1144), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(KEYINPUT124), .A4(KEYINPUT57), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1219), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1251), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1261), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1246), .B1(new_n1258), .B2(new_n1265), .ZN(G375));
  NAND2_X1  g1066(.A1(new_n1133), .A2(new_n1143), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1145), .A2(new_n1041), .A3(new_n1168), .A4(new_n1267), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n891), .A2(G13), .A3(G33), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n855), .B1(new_n291), .B2(new_n856), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n801), .A2(new_n869), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1235), .A2(new_n254), .ZN(new_n1272));
  AOI211_X1 g1072(.A(new_n1271), .B(new_n1272), .C1(G50), .C2(new_n803), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1273), .B1(new_n1191), .B2(new_n860), .C1(new_n404), .C2(new_n797), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT127), .Z(new_n1275));
  OAI22_X1  g1075(.A1(new_n1186), .A2(new_n812), .B1(new_n813), .B2(new_n1183), .ZN(new_n1276));
  OR3_X1    g1076(.A1(new_n808), .A2(KEYINPUT126), .A3(new_n876), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT126), .B1(new_n808), .B2(new_n876), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n254), .B1(new_n791), .B2(G77), .ZN(new_n1280));
  XOR2_X1   g1080(.A(new_n1280), .B(KEYINPUT125), .Z(new_n1281));
  OAI22_X1  g1081(.A1(new_n860), .A2(new_n615), .B1(new_n805), .B2(new_n808), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G283), .A2(new_n826), .B1(new_n829), .B2(new_n471), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1064), .C1(new_n245), .C2(new_n801), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1282), .B(new_n1284), .C1(new_n465), .C2(new_n827), .ZN(new_n1285));
  AOI22_X1  g1085(.A1(new_n1275), .A2(new_n1279), .B1(new_n1281), .B2(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1270), .B1(new_n1286), .B2(new_n858), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n1143), .A2(new_n1120), .B1(new_n1269), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1268), .A2(new_n1289), .ZN(G381));
  INV_X1    g1090(.A(G387), .ZN(new_n1291));
  NOR4_X1   g1091(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1292));
  INV_X1    g1092(.A(G378), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  OR3_X1    g1094(.A1(new_n1294), .A2(G390), .A3(G375), .ZN(G407));
  NAND2_X1  g1095(.A1(new_n681), .A2(G213), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G407), .B(G213), .C1(G375), .C2(new_n1298), .ZN(G409));
  OAI211_X1 g1099(.A(G378), .B(new_n1246), .C1(new_n1258), .C2(new_n1265), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1260), .A2(new_n775), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1259), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1245), .B(new_n1301), .C1(new_n1302), .C2(new_n1040), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1293), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1296), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1144), .A2(KEYINPUT60), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(new_n1267), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n770), .B1(new_n1307), .B2(new_n1267), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1289), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(G384), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  OAI211_X1 g1112(.A(G384), .B(new_n1289), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1297), .A2(G2897), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT61), .B1(new_n1306), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1128), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT118), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1291), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(G393), .B(G396), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1124), .A2(new_n1128), .A3(G387), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1324), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1324), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT63), .ZN(new_n1331));
  OAI21_X1  g1131(.A(new_n1331), .B1(new_n1306), .B2(new_n1314), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1297), .B1(new_n1300), .B2(new_n1304), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1314), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1333), .A2(KEYINPUT63), .A3(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1321), .A2(new_n1330), .A3(new_n1332), .A4(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1333), .A2(new_n1337), .A3(new_n1334), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT61), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1339), .B1(new_n1333), .B2(new_n1319), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1337), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1341));
  NOR3_X1   g1141(.A1(new_n1338), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1336), .B1(new_n1342), .B2(new_n1330), .ZN(G405));
  NAND2_X1  g1143(.A1(G375), .A2(new_n1293), .ZN(new_n1344));
  AND3_X1   g1144(.A1(new_n1344), .A2(new_n1314), .A3(new_n1300), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1314), .B1(new_n1344), .B2(new_n1300), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(new_n1347), .B(new_n1330), .ZN(G402));
endmodule


