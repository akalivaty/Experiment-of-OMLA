//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT65), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT66), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND3_X1   g036(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n462));
  AND3_X1   g037(.A1(KEYINPUT67), .A2(G113), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT67), .B1(G113), .B2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OAI21_X1  g042(.A(G125), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n469), .B2(G2105), .ZN(new_n470));
  OAI211_X1 g045(.A(G137), .B(new_n461), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT3), .B(G2104), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n474), .A2(KEYINPUT68), .A3(G137), .A4(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n466), .A2(new_n467), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n466), .C2(new_n467), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n466), .B2(new_n467), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n491), .B(new_n494), .C1(new_n467), .C2(new_n466), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n497));
  OAI21_X1  g072(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT69), .A2(G114), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n501), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n503), .B(KEYINPUT70), .C1(new_n499), .C2(new_n498), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n512), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  XOR2_X1   g089(.A(new_n514), .B(KEYINPUT72), .Z(new_n515));
  OAI21_X1  g090(.A(G651), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(G651), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n523), .A2(G50), .A3(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n523), .A2(G88), .A3(new_n512), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(G166));
  NAND2_X1  g102(.A1(new_n523), .A2(new_n512), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n532), .A2(new_n533), .B1(new_n512), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n523), .A2(new_n537), .A3(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n537), .B1(new_n523), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n536), .B1(new_n540), .B2(G51), .ZN(G168));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  XOR2_X1   g117(.A(KEYINPUT74), .B(G52), .Z(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n528), .A2(new_n545), .B1(new_n546), .B2(new_n517), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  NAND2_X1  g123(.A1(new_n540), .A2(G43), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n512), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n529), .A2(G81), .B1(new_n553), .B2(G651), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n521), .A2(new_n522), .ZN(new_n561));
  INV_X1    g136(.A(new_n518), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n561), .A2(G543), .A3(new_n562), .A4(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n512), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n517), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n565), .A2(new_n566), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n523), .A2(G91), .A3(new_n512), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n567), .A2(new_n569), .A3(new_n570), .A4(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n526), .A2(KEYINPUT76), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n516), .A2(new_n576), .A3(new_n524), .A4(new_n525), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n575), .A2(new_n577), .ZN(G303));
  INV_X1    g153(.A(KEYINPUT77), .ZN(new_n579));
  AND2_X1   g154(.A1(G49), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n579), .B1(new_n523), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n523), .A2(new_n579), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n523), .A2(G87), .A3(new_n512), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n584), .A2(new_n588), .ZN(G288));
  NAND3_X1  g164(.A1(new_n523), .A2(G48), .A3(G543), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n523), .A2(G86), .A3(new_n512), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n510), .B2(new_n511), .ZN(new_n593));
  AND2_X1   g168(.A1(G73), .A2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n591), .A3(new_n595), .ZN(G305));
  AND2_X1   g171(.A1(new_n540), .A2(G47), .ZN(new_n597));
  XOR2_X1   g172(.A(KEYINPUT78), .B(G85), .Z(new_n598));
  AOI22_X1  g173(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  OAI22_X1  g174(.A1(new_n528), .A2(new_n598), .B1(new_n599), .B2(new_n517), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n603), .B(KEYINPUT79), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n512), .A2(G66), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n517), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND4_X1  g182(.A1(new_n561), .A2(G92), .A3(new_n562), .A4(new_n512), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .A4(new_n512), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(G54), .B1(new_n538), .B2(new_n539), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n604), .B1(G868), .B2(new_n618), .ZN(G284));
  OAI21_X1  g194(.A(new_n604), .B1(G868), .B2(new_n618), .ZN(G321));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(G299), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G168), .B2(new_n621), .ZN(G297));
  OAI21_X1  g198(.A(new_n622), .B1(G168), .B2(new_n621), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n549), .A2(new_n554), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n621), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n617), .A2(G559), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(new_n629), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n480), .A2(G135), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT82), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n482), .A2(G123), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT83), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n636), .A2(new_n637), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n637), .B2(new_n636), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n635), .A3(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n461), .A2(G2104), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n479), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n647), .B(new_n648), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT13), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT88), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(KEYINPUT14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2451), .B(G2454), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n667), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(G401));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  XNOR2_X1  g248(.A(G2067), .B(G2678), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT17), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n672), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(G2100), .ZN(new_n679));
  XOR2_X1   g254(.A(G2072), .B(G2078), .Z(new_n680));
  AOI21_X1  g255(.A(new_n680), .B1(new_n675), .B2(KEYINPUT18), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(G2096), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n679), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(KEYINPUT20), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n686), .A2(new_n687), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(new_n693), .B(new_n692), .S(new_n685), .Z(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n698), .A2(new_n700), .ZN(new_n703));
  AND3_X1   g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n702), .B1(new_n701), .B2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(G229));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n707));
  AND3_X1   g282(.A1(new_n523), .A2(new_n579), .A3(new_n580), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(new_n581), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n707), .B1(new_n709), .B2(new_n587), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n584), .A2(new_n588), .A3(KEYINPUT92), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G16), .B2(G23), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT33), .B(G1976), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n715), .A2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G22), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  MUX2_X1   g298(.A(G6), .B(G305), .S(G16), .Z(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT32), .B(G1981), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NAND4_X1  g301(.A1(new_n717), .A2(new_n718), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n719), .A2(G24), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n601), .B2(new_n719), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n733), .A2(G1986), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(G1986), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G25), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n480), .A2(G131), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n482), .A2(G119), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT89), .B1(G95), .B2(G2105), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(KEYINPUT89), .A2(G95), .A3(G2105), .ZN(new_n742));
  OAI221_X1 g317(.A(G2104), .B1(G107), .B2(new_n461), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n738), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n737), .B1(new_n745), .B2(new_n736), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT35), .B(G1991), .Z(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT90), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n746), .B(new_n748), .Z(new_n749));
  NOR3_X1   g324(.A1(new_n734), .A2(new_n735), .A3(new_n749), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n730), .A2(new_n731), .A3(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT93), .B(KEYINPUT36), .Z(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n730), .A2(new_n731), .A3(new_n750), .A4(new_n752), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n736), .A2(G33), .ZN(new_n757));
  INV_X1    g332(.A(G127), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n479), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  OAI21_X1  g335(.A(G2105), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT97), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(KEYINPUT97), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT25), .ZN(new_n764));
  NAND2_X1  g339(.A1(G103), .A2(G2104), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(G2105), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n461), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n480), .A2(G139), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n762), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n757), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT98), .Z(new_n771));
  OAI21_X1  g346(.A(KEYINPUT99), .B1(new_n771), .B2(G2072), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n770), .B(KEYINPUT98), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT99), .ZN(new_n774));
  INV_X1    g349(.A(G2072), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n736), .A2(G32), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n480), .A2(G141), .ZN(new_n779));
  INV_X1    g354(.A(G105), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n646), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n482), .A2(G129), .ZN(new_n782));
  NAND3_X1  g357(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT26), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n778), .B1(new_n786), .B2(new_n736), .ZN(new_n787));
  XOR2_X1   g362(.A(KEYINPUT27), .B(G1996), .Z(new_n788));
  INV_X1    g363(.A(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(G29), .B1(new_n789), .B2(KEYINPUT24), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT24), .B2(new_n789), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(new_n477), .B2(new_n736), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n787), .A2(new_n788), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n771), .B2(G2072), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n777), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(KEYINPUT100), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT100), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n777), .A2(new_n798), .A3(new_n795), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n641), .B(KEYINPUT85), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(G29), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT102), .ZN(new_n802));
  NOR2_X1   g377(.A1(G16), .A2(G21), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G168), .B2(G16), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT101), .B(G1966), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n804), .B(new_n805), .Z(new_n806));
  AND2_X1   g381(.A1(new_n802), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT104), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n719), .A2(G5), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G171), .B2(new_n719), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT103), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT31), .B(G11), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT30), .B(G28), .Z(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G29), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n801), .B2(KEYINPUT102), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n807), .A2(new_n808), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n802), .A2(new_n818), .A3(new_n806), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT104), .B1(new_n820), .B2(new_n813), .ZN(new_n821));
  AND4_X1   g396(.A1(new_n797), .A2(new_n799), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n719), .A2(G19), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(new_n555), .B2(new_n719), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G1341), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n736), .A2(G35), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G162), .B2(new_n736), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT29), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(G2090), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n787), .A2(new_n788), .B1(new_n792), .B2(new_n793), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n736), .A2(G27), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G164), .B2(new_n736), .ZN(new_n832));
  INV_X1    g407(.A(G2078), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n829), .A2(new_n830), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT96), .B(KEYINPUT28), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n736), .A2(G26), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n480), .A2(G140), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n482), .A2(G128), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n461), .A2(G116), .ZN(new_n841));
  OAI21_X1  g416(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n839), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT94), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NOR3_X1   g420(.A1(new_n845), .A2(KEYINPUT95), .A3(new_n736), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n847), .B1(new_n844), .B2(G29), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n838), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(G2067), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g426(.A(G2067), .B(new_n838), .C1(new_n846), .C2(new_n848), .ZN(new_n852));
  AOI211_X1 g427(.A(new_n825), .B(new_n835), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(G4), .A2(G16), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n618), .B2(G16), .ZN(new_n855));
  INV_X1    g430(.A(G1348), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n811), .A2(new_n812), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n828), .A2(G2090), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n719), .A2(G20), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT23), .Z(new_n861));
  AOI21_X1  g436(.A(new_n861), .B1(G299), .B2(G16), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G1956), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT105), .ZN(new_n865));
  NAND4_X1  g440(.A1(new_n853), .A2(new_n857), .A3(new_n858), .A4(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n822), .A2(KEYINPUT106), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n797), .A2(new_n819), .A3(new_n799), .A4(new_n821), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n866), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n756), .B1(new_n868), .B2(new_n871), .ZN(G311));
  INV_X1    g447(.A(new_n756), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT106), .B1(new_n822), .B2(new_n867), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n870), .A2(new_n866), .A3(new_n869), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(G150));
  AOI22_X1  g451(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n877), .A2(new_n517), .ZN(new_n878));
  INV_X1    g453(.A(G93), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n878), .B1(new_n879), .B2(new_n528), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n540), .B2(G55), .ZN(new_n881));
  INV_X1    g456(.A(G860), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT37), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n617), .A2(new_n625), .ZN(new_n885));
  XOR2_X1   g460(.A(KEYINPUT107), .B(KEYINPUT38), .Z(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n555), .A2(new_n881), .ZN(new_n888));
  INV_X1    g463(.A(G55), .ZN(new_n889));
  OAI221_X1 g464(.A(new_n878), .B1(new_n879), .B2(new_n528), .C1(new_n542), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n627), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n887), .B(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n894), .A2(KEYINPUT39), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n882), .B1(new_n894), .B2(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n884), .B1(new_n895), .B2(new_n896), .ZN(G145));
  NAND2_X1  g472(.A1(new_n643), .A2(G162), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n800), .A2(new_n486), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(G160), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n844), .B(G164), .ZN(new_n902));
  INV_X1    g477(.A(new_n649), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n844), .B(new_n506), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n649), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n769), .B(new_n786), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n482), .A2(G130), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n461), .A2(G118), .ZN(new_n910));
  OAI21_X1  g485(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(G142), .B2(new_n480), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(new_n744), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(new_n914), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n904), .A2(new_n906), .A3(new_n915), .A4(new_n916), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(G37), .B1(new_n901), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n901), .A2(new_n920), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT108), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n901), .A2(new_n920), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n921), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g502(.A(new_n526), .B(G305), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G290), .A2(new_n712), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n713), .A2(new_n601), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n929), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n930), .A2(new_n931), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT110), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(KEYINPUT110), .A3(new_n929), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n629), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n892), .B(new_n940), .ZN(new_n941));
  OR2_X1    g516(.A1(G299), .A2(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g517(.A1(G299), .A2(KEYINPUT109), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n942), .A2(new_n613), .A3(new_n612), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n612), .A2(new_n613), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(KEYINPUT109), .A3(G299), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n941), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(KEYINPUT41), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n939), .B(new_n949), .C1(new_n941), .C2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n949), .B1(new_n941), .B2(new_n953), .ZN(new_n955));
  INV_X1    g530(.A(new_n938), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n934), .B2(new_n936), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT111), .B(KEYINPUT42), .Z(new_n959));
  AND3_X1   g534(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n954), .B2(new_n958), .ZN(new_n961));
  OAI21_X1  g536(.A(G868), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n890), .A2(new_n621), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(G295));
  NAND2_X1  g539(.A1(new_n962), .A2(new_n963), .ZN(G331));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n888), .A2(G286), .A3(new_n891), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(G286), .B1(new_n888), .B2(new_n891), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n968), .A2(new_n969), .A3(G301), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n892), .A2(G168), .ZN(new_n971));
  AOI21_X1  g546(.A(G171), .B1(new_n971), .B2(new_n967), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n948), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(G301), .B1(new_n968), .B2(new_n969), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n971), .A2(G171), .A3(new_n967), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n950), .A4(new_n952), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n939), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n957), .A2(new_n973), .A3(new_n976), .ZN(new_n980));
  AND3_X1   g555(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n979), .B1(new_n978), .B2(new_n980), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n966), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n978), .A2(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n978), .A2(new_n979), .A3(new_n980), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(KEYINPUT44), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n987), .ZN(G397));
  INV_X1    g563(.A(G1384), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n502), .A2(new_n504), .ZN(new_n990));
  INV_X1    g565(.A(new_n495), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n494), .B1(new_n474), .B2(new_n491), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n488), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n989), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n998), .B(KEYINPUT114), .Z(new_n999));
  XNOR2_X1  g574(.A(new_n844), .B(G2067), .ZN(new_n1000));
  INV_X1    g575(.A(new_n786), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n1004), .B(KEYINPUT46), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT47), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n786), .A2(new_n1003), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n999), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  XOR2_X1   g586(.A(new_n744), .B(new_n748), .Z(new_n1012));
  NAND2_X1  g587(.A1(new_n999), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g589(.A1(G290), .A2(G1986), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1015), .A2(new_n996), .A3(new_n997), .ZN(new_n1016));
  XOR2_X1   g591(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1017));
  XNOR2_X1  g592(.A(new_n1016), .B(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1007), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n745), .A2(new_n748), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT125), .Z(new_n1021));
  OAI22_X1  g596(.A1(new_n1010), .A2(new_n1021), .B1(G2067), .B2(new_n844), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1019), .B1(new_n999), .B2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1384), .B1(new_n496), .B2(new_n505), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI211_X1 g602(.A(KEYINPUT50), .B(G1384), .C1(new_n496), .C2(new_n505), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n856), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1024), .A2(new_n1025), .A3(new_n850), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n617), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1032));
  XNOR2_X1  g607(.A(G299), .B(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1956), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n995), .A2(G1384), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n506), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1037), .ZN(new_n1039));
  AOI211_X1 g614(.A(KEYINPUT115), .B(new_n1039), .C1(new_n496), .C2(new_n505), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n996), .B(new_n1024), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(KEYINPUT119), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1035), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1033), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n997), .B1(new_n994), .B2(new_n995), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n1043), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT121), .A3(new_n1035), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1031), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1033), .B(new_n1035), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n1054));
  XNOR2_X1  g629(.A(new_n1053), .B(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1029), .A2(new_n617), .A3(new_n1030), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT60), .B1(new_n1057), .B2(new_n1031), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT60), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n618), .A2(new_n1059), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n1061));
  XOR2_X1   g636(.A(KEYINPUT122), .B(G1996), .Z(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1049), .B(new_n1063), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT58), .B(G1341), .Z(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n994), .B2(new_n997), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1061), .B1(new_n1067), .B2(new_n555), .ZN(new_n1068));
  AOI211_X1 g643(.A(KEYINPUT59), .B(new_n627), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1058), .B(new_n1060), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1053), .A2(KEYINPUT61), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1047), .B2(new_n1051), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1033), .B1(new_n1050), .B2(new_n1035), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1055), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1056), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1037), .B1(new_n990), .B2(new_n993), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1024), .C1(new_n1025), .C2(KEYINPUT45), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  INV_X1    g655(.A(G1966), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n997), .B1(new_n994), .B2(KEYINPUT50), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1028), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n793), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1080), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1087));
  OAI21_X1  g662(.A(G286), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT116), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1090), .A2(G168), .A3(new_n1085), .A4(new_n1082), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(G8), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT51), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(new_n1094), .A3(G8), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n710), .A2(new_n711), .A3(G1976), .ZN(new_n1097));
  INV_X1    g672(.A(G8), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1098), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(KEYINPUT52), .ZN(new_n1101));
  INV_X1    g676(.A(G1976), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT52), .B1(G288), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1097), .A2(new_n1103), .A3(new_n1099), .ZN(new_n1104));
  NAND2_X1  g679(.A1(G305), .A2(G1981), .ZN(new_n1105));
  INV_X1    g680(.A(G1981), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n590), .A2(new_n591), .A3(new_n595), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT49), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(KEYINPUT49), .A3(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1099), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1101), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1041), .A2(new_n722), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1115));
  INV_X1    g690(.A(G2090), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1098), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n575), .A2(G8), .A3(new_n577), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT55), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n575), .A2(KEYINPUT55), .A3(G8), .A4(new_n577), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1113), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1123), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1041), .A2(new_n722), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n1098), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1124), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1049), .B(new_n833), .C1(new_n1038), .C2(new_n1040), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1048), .A2(KEYINPUT53), .A3(new_n833), .A4(new_n1049), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n812), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(KEYINPUT124), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(new_n1137), .A3(new_n812), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .A4(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1130), .A2(new_n1131), .B1(new_n812), .B2(new_n1136), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1079), .B2(G2078), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1049), .A2(KEYINPUT123), .A3(new_n833), .A4(new_n1078), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(KEYINPUT53), .ZN(new_n1145));
  AOI21_X1  g720(.A(G301), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1129), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1139), .A2(G171), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1141), .A2(G301), .A3(new_n1145), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1148), .A2(KEYINPUT54), .A3(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1096), .A2(new_n1128), .A3(new_n1147), .A4(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(G1971), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1136), .A2(G2090), .ZN(new_n1153));
  OAI211_X1 g728(.A(G8), .B(new_n1123), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(new_n1099), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1107), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G288), .A2(G1976), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1112), .B2(new_n1157), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1154), .A2(new_n1113), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(G168), .A2(G8), .ZN(new_n1160));
  AND2_X1   g735(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1160), .B1(new_n1161), .B2(new_n1090), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1101), .A2(new_n1104), .A3(new_n1112), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1162), .A2(new_n1127), .A3(new_n1163), .A4(new_n1154), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1124), .A2(KEYINPUT63), .A3(new_n1127), .A4(new_n1162), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1159), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI22_X1  g743(.A1(new_n1077), .A2(new_n1151), .B1(new_n1168), .B2(KEYINPUT117), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1096), .A2(KEYINPUT62), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1128), .A2(new_n1146), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT62), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT117), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1175), .B(new_n1159), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1169), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(G290), .A2(G1986), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1015), .A2(KEYINPUT113), .A3(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1179), .B(new_n998), .C1(KEYINPUT113), .C2(new_n1178), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1011), .A2(new_n1180), .A3(new_n1013), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1023), .B1(new_n1177), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g757(.A(new_n459), .B(G227), .C1(new_n669), .C2(new_n670), .ZN(new_n1184));
  OAI21_X1  g758(.A(new_n1184), .B1(new_n704), .B2(new_n705), .ZN(new_n1185));
  INV_X1    g759(.A(KEYINPUT127), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OAI211_X1 g761(.A(new_n1184), .B(KEYINPUT127), .C1(new_n704), .C2(new_n705), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI211_X1 g763(.A(new_n926), .B(new_n1189), .C1(new_n981), .C2(new_n982), .ZN(G225));
  INV_X1    g764(.A(G225), .ZN(G308));
endmodule


