

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U552 ( .A(KEYINPUT95), .B(n599), .Z(n705) );
  NOR2_X1 U553 ( .A1(n526), .A2(G2104), .ZN(n908) );
  XNOR2_X1 U554 ( .A(n654), .B(n653), .ZN(n656) );
  XNOR2_X1 U555 ( .A(n683), .B(KEYINPUT103), .ZN(n684) );
  NOR2_X1 U556 ( .A1(G651), .A2(G543), .ZN(n805) );
  INV_X1 U557 ( .A(KEYINPUT85), .ZN(n533) );
  NOR2_X2 U558 ( .A1(n530), .A2(n529), .ZN(G160) );
  XOR2_X1 U559 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n518) );
  AND2_X1 U560 ( .A1(n656), .A2(n655), .ZN(n519) );
  NOR2_X1 U561 ( .A1(n667), .A2(n664), .ZN(n652) );
  XNOR2_X1 U562 ( .A(KEYINPUT99), .B(KEYINPUT30), .ZN(n653) );
  INV_X1 U563 ( .A(G168), .ZN(n655) );
  INV_X1 U564 ( .A(KEYINPUT100), .ZN(n658) );
  XNOR2_X1 U565 ( .A(n658), .B(KEYINPUT31), .ZN(n659) );
  BUF_X1 U566 ( .A(n600), .Z(n670) );
  INV_X1 U567 ( .A(KEYINPUT101), .ZN(n665) );
  NAND2_X1 U568 ( .A1(n600), .A2(G8), .ZN(n599) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n520) );
  NOR2_X1 U570 ( .A1(KEYINPUT88), .A2(n732), .ZN(n747) );
  AND2_X1 U571 ( .A1(G2104), .A2(n526), .ZN(n527) );
  AND2_X1 U572 ( .A1(G2105), .A2(G2104), .ZN(n909) );
  XNOR2_X1 U573 ( .A(n527), .B(KEYINPUT64), .ZN(n714) );
  NOR2_X1 U574 ( .A1(G651), .A2(n577), .ZN(n801) );
  XNOR2_X1 U575 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U576 ( .A(KEYINPUT17), .B(n520), .Z(n531) );
  NAND2_X1 U577 ( .A1(G137), .A2(n531), .ZN(n522) );
  NAND2_X1 U578 ( .A1(G113), .A2(n909), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U580 ( .A(n523), .B(KEYINPUT65), .ZN(n525) );
  INV_X1 U581 ( .A(G2105), .ZN(n526) );
  NAND2_X1 U582 ( .A1(G125), .A2(n908), .ZN(n524) );
  NAND2_X1 U583 ( .A1(n525), .A2(n524), .ZN(n530) );
  NAND2_X1 U584 ( .A1(G101), .A2(n714), .ZN(n528) );
  XNOR2_X1 U585 ( .A(KEYINPUT23), .B(n528), .ZN(n529) );
  INV_X1 U586 ( .A(n531), .ZN(n532) );
  INV_X1 U587 ( .A(n532), .ZN(n904) );
  NAND2_X1 U588 ( .A1(n904), .A2(G138), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n714), .A2(G102), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G126), .A2(n908), .ZN(n538) );
  NAND2_X1 U592 ( .A1(G114), .A2(n909), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n539) );
  NOR2_X1 U594 ( .A1(n540), .A2(n539), .ZN(G164) );
  NAND2_X1 U595 ( .A1(n805), .A2(G90), .ZN(n542) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n577) );
  XOR2_X1 U597 ( .A(G651), .B(KEYINPUT66), .Z(n546) );
  NOR2_X1 U598 ( .A1(n577), .A2(n546), .ZN(n806) );
  NAND2_X1 U599 ( .A1(G77), .A2(n806), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n545) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(KEYINPUT69), .Z(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT70), .B(n543), .ZN(n544) );
  XNOR2_X1 U603 ( .A(n545), .B(n544), .ZN(n551) );
  NOR2_X1 U604 ( .A1(G543), .A2(n546), .ZN(n547) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n547), .Z(n802) );
  NAND2_X1 U606 ( .A1(n802), .A2(G64), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n801), .A2(G52), .ZN(n548) );
  AND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(G301) );
  INV_X1 U610 ( .A(G301), .ZN(G171) );
  NAND2_X1 U611 ( .A1(n801), .A2(G53), .ZN(n553) );
  NAND2_X1 U612 ( .A1(G65), .A2(n802), .ZN(n552) );
  NAND2_X1 U613 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U614 ( .A(KEYINPUT72), .B(n554), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G78), .A2(n806), .ZN(n555) );
  XNOR2_X1 U616 ( .A(KEYINPUT71), .B(n555), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n805), .A2(G91), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(G299) );
  NAND2_X1 U620 ( .A1(n805), .A2(G89), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT4), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G76), .A2(n806), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n563), .B(KEYINPUT5), .ZN(n569) );
  NAND2_X1 U625 ( .A1(n801), .A2(G51), .ZN(n564) );
  XNOR2_X1 U626 ( .A(n564), .B(KEYINPUT76), .ZN(n566) );
  NAND2_X1 U627 ( .A1(G63), .A2(n802), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n567), .Z(n568) );
  NAND2_X1 U630 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U631 ( .A(n570), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U632 ( .A1(n805), .A2(G88), .ZN(n572) );
  NAND2_X1 U633 ( .A1(G75), .A2(n806), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n572), .A2(n571), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n801), .A2(G50), .ZN(n574) );
  NAND2_X1 U636 ( .A1(G62), .A2(n802), .ZN(n573) );
  NAND2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U638 ( .A1(n576), .A2(n575), .ZN(G166) );
  XOR2_X1 U639 ( .A(KEYINPUT86), .B(G166), .Z(G303) );
  XOR2_X1 U640 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U641 ( .A1(G87), .A2(n577), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n802), .A2(n580), .ZN(n582) );
  NAND2_X1 U645 ( .A1(n801), .A2(G49), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(G288) );
  NAND2_X1 U647 ( .A1(G48), .A2(n801), .ZN(n584) );
  NAND2_X1 U648 ( .A1(G86), .A2(n805), .ZN(n583) );
  NAND2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n806), .A2(G73), .ZN(n585) );
  XOR2_X1 U651 ( .A(KEYINPUT2), .B(n585), .Z(n586) );
  NOR2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G61), .A2(n802), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(G305) );
  NAND2_X1 U655 ( .A1(n801), .A2(G47), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G60), .A2(n802), .ZN(n590) );
  NAND2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U658 ( .A(KEYINPUT68), .B(n592), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G72), .A2(n806), .ZN(n593) );
  XNOR2_X1 U660 ( .A(KEYINPUT67), .B(n593), .ZN(n594) );
  NOR2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n805), .A2(G85), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n597), .A2(n596), .ZN(G290) );
  NAND2_X1 U664 ( .A1(G160), .A2(G40), .ZN(n710) );
  INV_X1 U665 ( .A(n710), .ZN(n598) );
  NOR2_X1 U666 ( .A1(G164), .A2(G1384), .ZN(n711) );
  NAND2_X1 U667 ( .A1(n598), .A2(n711), .ZN(n600) );
  NOR2_X1 U668 ( .A1(G1966), .A2(n705), .ZN(n664) );
  XNOR2_X1 U669 ( .A(n600), .B(KEYINPUT96), .ZN(n605) );
  INV_X1 U670 ( .A(n605), .ZN(n636) );
  XNOR2_X1 U671 ( .A(G2078), .B(KEYINPUT25), .ZN(n964) );
  NAND2_X1 U672 ( .A1(n636), .A2(n964), .ZN(n602) );
  INV_X1 U673 ( .A(G1961), .ZN(n1007) );
  NAND2_X1 U674 ( .A1(n1007), .A2(n670), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(n651) );
  NAND2_X1 U676 ( .A1(n651), .A2(G171), .ZN(n650) );
  NAND2_X1 U677 ( .A1(G2072), .A2(n636), .ZN(n603) );
  XNOR2_X1 U678 ( .A(KEYINPUT27), .B(n603), .ZN(n604) );
  INV_X1 U679 ( .A(n604), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n605), .A2(G1956), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U682 ( .A1(G299), .A2(n610), .ZN(n609) );
  XOR2_X1 U683 ( .A(KEYINPUT97), .B(KEYINPUT28), .Z(n608) );
  XNOR2_X1 U684 ( .A(n609), .B(n608), .ZN(n646) );
  NOR2_X1 U685 ( .A1(G299), .A2(n610), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT98), .B(n611), .Z(n644) );
  NAND2_X1 U687 ( .A1(n805), .A2(G92), .ZN(n613) );
  NAND2_X1 U688 ( .A1(G79), .A2(n806), .ZN(n612) );
  NAND2_X1 U689 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n801), .A2(G54), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G66), .A2(n802), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U694 ( .A(KEYINPUT15), .B(n618), .Z(n987) );
  NAND2_X1 U695 ( .A1(G81), .A2(n805), .ZN(n619) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT12), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n620), .B(KEYINPUT74), .ZN(n622) );
  NAND2_X1 U698 ( .A1(G68), .A2(n806), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U700 ( .A(KEYINPUT13), .B(n623), .ZN(n629) );
  NAND2_X1 U701 ( .A1(n802), .A2(G56), .ZN(n624) );
  XOR2_X1 U702 ( .A(KEYINPUT14), .B(n624), .Z(n627) );
  NAND2_X1 U703 ( .A1(G43), .A2(n801), .ZN(n625) );
  XNOR2_X1 U704 ( .A(KEYINPUT75), .B(n625), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n982) );
  INV_X1 U707 ( .A(G1996), .ZN(n630) );
  NOR2_X1 U708 ( .A1(n600), .A2(n630), .ZN(n631) );
  XOR2_X1 U709 ( .A(n631), .B(KEYINPUT26), .Z(n633) );
  NAND2_X1 U710 ( .A1(n670), .A2(G1341), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U712 ( .A1(n982), .A2(n634), .ZN(n635) );
  OR2_X1 U713 ( .A1(n987), .A2(n635), .ZN(n642) );
  NAND2_X1 U714 ( .A1(n987), .A2(n635), .ZN(n640) );
  NAND2_X1 U715 ( .A1(G2067), .A2(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(G1348), .A2(n670), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n646), .A2(n645), .ZN(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT29), .B(n647), .ZN(n648) );
  INV_X1 U723 ( .A(n648), .ZN(n649) );
  NAND2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n662) );
  NOR2_X1 U725 ( .A1(G171), .A2(n651), .ZN(n657) );
  NOR2_X1 U726 ( .A1(G2084), .A2(n670), .ZN(n667) );
  NAND2_X1 U727 ( .A1(G8), .A2(n652), .ZN(n654) );
  NOR2_X1 U728 ( .A1(n657), .A2(n519), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n675) );
  INV_X1 U731 ( .A(n675), .ZN(n663) );
  NOR2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n669) );
  NAND2_X1 U734 ( .A1(G8), .A2(n667), .ZN(n668) );
  NAND2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n681) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n705), .ZN(n672) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n670), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U739 ( .A1(G303), .A2(n673), .ZN(n674) );
  XNOR2_X1 U740 ( .A(n674), .B(KEYINPUT102), .ZN(n677) );
  NAND2_X1 U741 ( .A1(G286), .A2(n675), .ZN(n676) );
  NAND2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U743 ( .A1(G8), .A2(n678), .ZN(n679) );
  XNOR2_X1 U744 ( .A(KEYINPUT32), .B(n679), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n681), .A2(n680), .ZN(n701) );
  NOR2_X1 U746 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U747 ( .A1(G303), .A2(G1971), .ZN(n682) );
  NOR2_X1 U748 ( .A1(n685), .A2(n682), .ZN(n995) );
  NAND2_X1 U749 ( .A1(n701), .A2(n995), .ZN(n683) );
  NOR2_X1 U750 ( .A1(n684), .A2(n705), .ZN(n692) );
  NAND2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n994) );
  INV_X1 U752 ( .A(KEYINPUT33), .ZN(n694) );
  INV_X1 U753 ( .A(n705), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n694), .A2(n687), .ZN(n688) );
  XOR2_X1 U756 ( .A(n688), .B(KEYINPUT104), .Z(n693) );
  AND2_X1 U757 ( .A1(n994), .A2(n693), .ZN(n690) );
  XNOR2_X1 U758 ( .A(G1981), .B(G305), .ZN(n992) );
  INV_X1 U759 ( .A(n992), .ZN(n689) );
  AND2_X1 U760 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n709) );
  INV_X1 U762 ( .A(n693), .ZN(n695) );
  OR2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n992), .A2(n696), .ZN(n700) );
  NOR2_X1 U765 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U766 ( .A(n697), .B(KEYINPUT24), .Z(n698) );
  NOR2_X1 U767 ( .A1(n705), .A2(n698), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n707) );
  NOR2_X1 U769 ( .A1(G2090), .A2(G303), .ZN(n702) );
  NAND2_X1 U770 ( .A1(G8), .A2(n702), .ZN(n703) );
  NAND2_X1 U771 ( .A1(n701), .A2(n703), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  AND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n764) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n768) );
  XNOR2_X1 U776 ( .A(KEYINPUT94), .B(n768), .ZN(n731) );
  NAND2_X1 U777 ( .A1(n904), .A2(G141), .ZN(n720) );
  NAND2_X1 U778 ( .A1(G129), .A2(n908), .ZN(n713) );
  NAND2_X1 U779 ( .A1(G117), .A2(n909), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n718) );
  INV_X1 U781 ( .A(n714), .ZN(n715) );
  INV_X1 U782 ( .A(n715), .ZN(n905) );
  NAND2_X1 U783 ( .A1(n905), .A2(G105), .ZN(n716) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n716), .Z(n717) );
  NOR2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U787 ( .A(KEYINPUT93), .B(n721), .Z(n900) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n900), .ZN(n730) );
  NAND2_X1 U789 ( .A1(G119), .A2(n908), .ZN(n723) );
  NAND2_X1 U790 ( .A1(G107), .A2(n909), .ZN(n722) );
  NAND2_X1 U791 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U792 ( .A1(n904), .A2(G131), .ZN(n724) );
  XOR2_X1 U793 ( .A(KEYINPUT92), .B(n724), .Z(n725) );
  NOR2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U795 ( .A1(G95), .A2(n905), .ZN(n727) );
  NAND2_X1 U796 ( .A1(n728), .A2(n727), .ZN(n915) );
  NAND2_X1 U797 ( .A1(G1991), .A2(n915), .ZN(n729) );
  NAND2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n942) );
  NAND2_X1 U799 ( .A1(n731), .A2(n942), .ZN(n758) );
  NAND2_X1 U800 ( .A1(n764), .A2(n758), .ZN(n732) );
  XOR2_X1 U801 ( .A(KEYINPUT87), .B(G1986), .Z(n733) );
  XNOR2_X1 U802 ( .A(G290), .B(n733), .ZN(n1002) );
  XNOR2_X1 U803 ( .A(G2067), .B(KEYINPUT37), .ZN(n748) );
  NAND2_X1 U804 ( .A1(n908), .A2(G128), .ZN(n734) );
  XOR2_X1 U805 ( .A(KEYINPUT91), .B(n734), .Z(n736) );
  NAND2_X1 U806 ( .A1(n909), .A2(G116), .ZN(n735) );
  NAND2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n737) );
  XOR2_X1 U808 ( .A(KEYINPUT35), .B(n737), .Z(n744) );
  NAND2_X1 U809 ( .A1(n905), .A2(G104), .ZN(n740) );
  NAND2_X1 U810 ( .A1(n904), .A2(G140), .ZN(n738) );
  XOR2_X1 U811 ( .A(KEYINPUT89), .B(n738), .Z(n739) );
  NAND2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U813 ( .A(n741), .B(KEYINPUT90), .ZN(n742) );
  XNOR2_X1 U814 ( .A(n742), .B(KEYINPUT34), .ZN(n743) );
  NOR2_X1 U815 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U816 ( .A(KEYINPUT36), .B(n745), .ZN(n919) );
  NOR2_X1 U817 ( .A1(n748), .A2(n919), .ZN(n954) );
  NAND2_X1 U818 ( .A1(n954), .A2(n768), .ZN(n749) );
  AND2_X1 U819 ( .A1(n1002), .A2(n749), .ZN(n746) );
  NAND2_X1 U820 ( .A1(n747), .A2(n746), .ZN(n767) );
  NAND2_X1 U821 ( .A1(n748), .A2(n919), .ZN(n951) );
  INV_X1 U822 ( .A(n749), .ZN(n759) );
  NOR2_X1 U823 ( .A1(G1996), .A2(n900), .ZN(n947) );
  INV_X1 U824 ( .A(n758), .ZN(n753) );
  NOR2_X1 U825 ( .A1(G1991), .A2(n915), .ZN(n943) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n750) );
  XOR2_X1 U827 ( .A(n750), .B(KEYINPUT105), .Z(n751) );
  NOR2_X1 U828 ( .A1(n943), .A2(n751), .ZN(n752) );
  NOR2_X1 U829 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U830 ( .A1(n947), .A2(n754), .ZN(n755) );
  XOR2_X1 U831 ( .A(KEYINPUT39), .B(n755), .Z(n756) );
  OR2_X1 U832 ( .A1(n759), .A2(n756), .ZN(n757) );
  AND2_X1 U833 ( .A1(n951), .A2(n757), .ZN(n765) );
  NAND2_X1 U834 ( .A1(n1002), .A2(n768), .ZN(n762) );
  NAND2_X1 U835 ( .A1(KEYINPUT88), .A2(n758), .ZN(n760) );
  NOR2_X1 U836 ( .A1(n760), .A2(n759), .ZN(n761) );
  AND2_X1 U837 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U838 ( .A1(n764), .A2(n763), .ZN(n770) );
  AND2_X1 U839 ( .A1(n765), .A2(n770), .ZN(n766) );
  NAND2_X1 U840 ( .A1(n767), .A2(n766), .ZN(n772) );
  INV_X1 U841 ( .A(n768), .ZN(n769) );
  NAND2_X1 U842 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U843 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U844 ( .A(n773), .B(n518), .ZN(G329) );
  AND2_X1 U845 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U846 ( .A(G57), .ZN(G237) );
  INV_X1 U847 ( .A(G132), .ZN(G219) );
  NAND2_X1 U848 ( .A1(G7), .A2(G661), .ZN(n774) );
  XNOR2_X1 U849 ( .A(n774), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U850 ( .A(G223), .ZN(n846) );
  NAND2_X1 U851 ( .A1(n846), .A2(G567), .ZN(n775) );
  XOR2_X1 U852 ( .A(KEYINPUT11), .B(n775), .Z(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n780) );
  OR2_X1 U854 ( .A1(n982), .A2(n780), .ZN(G153) );
  NAND2_X1 U855 ( .A1(G868), .A2(G301), .ZN(n777) );
  OR2_X1 U856 ( .A1(n987), .A2(G868), .ZN(n776) );
  NAND2_X1 U857 ( .A1(n777), .A2(n776), .ZN(G284) );
  INV_X1 U858 ( .A(G868), .ZN(n817) );
  NOR2_X1 U859 ( .A1(G286), .A2(n817), .ZN(n779) );
  NOR2_X1 U860 ( .A1(G868), .A2(G299), .ZN(n778) );
  NOR2_X1 U861 ( .A1(n779), .A2(n778), .ZN(G297) );
  NAND2_X1 U862 ( .A1(n780), .A2(G559), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n781), .A2(n987), .ZN(n782) );
  XNOR2_X1 U864 ( .A(n782), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n982), .ZN(n785) );
  NAND2_X1 U866 ( .A1(G868), .A2(n987), .ZN(n783) );
  NOR2_X1 U867 ( .A1(G559), .A2(n783), .ZN(n784) );
  NOR2_X1 U868 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U869 ( .A(KEYINPUT77), .B(n786), .Z(G282) );
  NAND2_X1 U870 ( .A1(G123), .A2(n908), .ZN(n787) );
  XNOR2_X1 U871 ( .A(n787), .B(KEYINPUT78), .ZN(n788) );
  XNOR2_X1 U872 ( .A(n788), .B(KEYINPUT18), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G111), .A2(n909), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U875 ( .A1(G135), .A2(n904), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G99), .A2(n905), .ZN(n791) );
  NAND2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U878 ( .A1(n794), .A2(n793), .ZN(n941) );
  XNOR2_X1 U879 ( .A(n941), .B(G2096), .ZN(n796) );
  INV_X1 U880 ( .A(G2100), .ZN(n795) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G559), .A2(n987), .ZN(n797) );
  XNOR2_X1 U883 ( .A(n797), .B(n982), .ZN(n854) );
  XNOR2_X1 U884 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n799) );
  XNOR2_X1 U885 ( .A(G288), .B(KEYINPUT80), .ZN(n798) );
  XNOR2_X1 U886 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U887 ( .A(G166), .B(n800), .ZN(n814) );
  NAND2_X1 U888 ( .A1(n801), .A2(G55), .ZN(n804) );
  NAND2_X1 U889 ( .A1(G67), .A2(n802), .ZN(n803) );
  NAND2_X1 U890 ( .A1(n804), .A2(n803), .ZN(n810) );
  NAND2_X1 U891 ( .A1(n805), .A2(G93), .ZN(n808) );
  NAND2_X1 U892 ( .A1(G80), .A2(n806), .ZN(n807) );
  NAND2_X1 U893 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U894 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U895 ( .A(n811), .B(KEYINPUT79), .ZN(n855) );
  XOR2_X1 U896 ( .A(n855), .B(G299), .Z(n812) );
  XNOR2_X1 U897 ( .A(n812), .B(G305), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U899 ( .A(n815), .B(G290), .ZN(n925) );
  XNOR2_X1 U900 ( .A(n854), .B(n925), .ZN(n816) );
  NAND2_X1 U901 ( .A1(n816), .A2(G868), .ZN(n819) );
  NAND2_X1 U902 ( .A1(n817), .A2(n855), .ZN(n818) );
  NAND2_X1 U903 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U904 ( .A1(G2084), .A2(G2078), .ZN(n820) );
  XOR2_X1 U905 ( .A(KEYINPUT20), .B(n820), .Z(n821) );
  NAND2_X1 U906 ( .A1(G2090), .A2(n821), .ZN(n823) );
  XNOR2_X1 U907 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n822) );
  XNOR2_X1 U908 ( .A(n823), .B(n822), .ZN(n824) );
  NAND2_X1 U909 ( .A1(G2072), .A2(n824), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U911 ( .A(KEYINPUT73), .B(G82), .ZN(G220) );
  NOR2_X1 U912 ( .A1(G219), .A2(G220), .ZN(n825) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n825), .Z(n826) );
  NOR2_X1 U914 ( .A1(G218), .A2(n826), .ZN(n827) );
  NAND2_X1 U915 ( .A1(G96), .A2(n827), .ZN(n852) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n852), .ZN(n831) );
  NAND2_X1 U917 ( .A1(G69), .A2(G120), .ZN(n828) );
  NOR2_X1 U918 ( .A1(G237), .A2(n828), .ZN(n829) );
  NAND2_X1 U919 ( .A1(G108), .A2(n829), .ZN(n853) );
  NAND2_X1 U920 ( .A1(G567), .A2(n853), .ZN(n830) );
  NAND2_X1 U921 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U922 ( .A(KEYINPUT83), .B(n832), .ZN(G319) );
  INV_X1 U923 ( .A(G319), .ZN(n834) );
  NAND2_X1 U924 ( .A1(G661), .A2(G483), .ZN(n833) );
  NOR2_X1 U925 ( .A1(n834), .A2(n833), .ZN(n849) );
  NAND2_X1 U926 ( .A1(n849), .A2(G36), .ZN(n835) );
  XNOR2_X1 U927 ( .A(KEYINPUT84), .B(n835), .ZN(G176) );
  XOR2_X1 U928 ( .A(G2454), .B(G2430), .Z(n837) );
  XNOR2_X1 U929 ( .A(G2451), .B(G2446), .ZN(n836) );
  XNOR2_X1 U930 ( .A(n837), .B(n836), .ZN(n844) );
  XOR2_X1 U931 ( .A(G2443), .B(G2427), .Z(n839) );
  XNOR2_X1 U932 ( .A(G2438), .B(KEYINPUT107), .ZN(n838) );
  XNOR2_X1 U933 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U934 ( .A(n840), .B(G2435), .Z(n842) );
  XNOR2_X1 U935 ( .A(G1341), .B(G1348), .ZN(n841) );
  XNOR2_X1 U936 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U937 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U938 ( .A1(n845), .A2(G14), .ZN(n930) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(n930), .Z(G401) );
  NAND2_X1 U940 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U941 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U942 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U943 ( .A1(G3), .A2(G1), .ZN(n848) );
  XOR2_X1 U944 ( .A(KEYINPUT109), .B(n848), .Z(n850) );
  NAND2_X1 U945 ( .A1(n850), .A2(n849), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n851), .B(KEYINPUT110), .ZN(G188) );
  INV_X1 U948 ( .A(G120), .ZN(G236) );
  INV_X1 U949 ( .A(G96), .ZN(G221) );
  INV_X1 U950 ( .A(G69), .ZN(G235) );
  NOR2_X1 U951 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U952 ( .A(G325), .ZN(G261) );
  NOR2_X1 U953 ( .A1(n854), .A2(G860), .ZN(n856) );
  XOR2_X1 U954 ( .A(n856), .B(n855), .Z(G145) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1986), .B(G1961), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U958 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n860) );
  XNOR2_X1 U959 ( .A(G1956), .B(KEYINPUT119), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n872) );
  XOR2_X1 U962 ( .A(KEYINPUT113), .B(KEYINPUT118), .Z(n864) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(n868) );
  XOR2_X1 U965 ( .A(KEYINPUT117), .B(KEYINPUT41), .Z(n866) );
  XNOR2_X1 U966 ( .A(KEYINPUT116), .B(G2474), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U968 ( .A(n868), .B(n867), .Z(n870) );
  XNOR2_X1 U969 ( .A(G1966), .B(G1981), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(G229) );
  XOR2_X1 U972 ( .A(KEYINPUT112), .B(KEYINPUT111), .Z(n874) );
  XNOR2_X1 U973 ( .A(G2678), .B(KEYINPUT43), .ZN(n873) );
  XNOR2_X1 U974 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U975 ( .A(KEYINPUT42), .B(G2090), .Z(n876) );
  XNOR2_X1 U976 ( .A(G2067), .B(G2072), .ZN(n875) );
  XNOR2_X1 U977 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U978 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U979 ( .A(G2096), .B(G2100), .ZN(n879) );
  XNOR2_X1 U980 ( .A(n880), .B(n879), .ZN(n882) );
  XOR2_X1 U981 ( .A(G2084), .B(G2078), .Z(n881) );
  XNOR2_X1 U982 ( .A(n882), .B(n881), .ZN(G227) );
  NAND2_X1 U983 ( .A1(n908), .A2(G124), .ZN(n884) );
  XNOR2_X1 U984 ( .A(KEYINPUT120), .B(KEYINPUT44), .ZN(n883) );
  XNOR2_X1 U985 ( .A(n884), .B(n883), .ZN(n891) );
  NAND2_X1 U986 ( .A1(G136), .A2(n904), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G100), .A2(n905), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G112), .A2(n909), .ZN(n887) );
  XNOR2_X1 U990 ( .A(KEYINPUT121), .B(n887), .ZN(n888) );
  NOR2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(KEYINPUT122), .B(n892), .Z(G162) );
  NAND2_X1 U994 ( .A1(G130), .A2(n908), .ZN(n894) );
  NAND2_X1 U995 ( .A1(G118), .A2(n909), .ZN(n893) );
  NAND2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n899) );
  NAND2_X1 U997 ( .A1(G142), .A2(n904), .ZN(n896) );
  NAND2_X1 U998 ( .A1(G106), .A2(n905), .ZN(n895) );
  NAND2_X1 U999 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U1000 ( .A(n897), .B(KEYINPUT45), .Z(n898) );
  NOR2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U1002 ( .A(n901), .B(n900), .ZN(n923) );
  XOR2_X1 U1003 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n903) );
  XNOR2_X1 U1004 ( .A(G160), .B(n941), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(n903), .B(n902), .ZN(n918) );
  NAND2_X1 U1006 ( .A1(G139), .A2(n904), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(G103), .A2(n905), .ZN(n906) );
  NAND2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n914) );
  NAND2_X1 U1009 ( .A1(G127), .A2(n908), .ZN(n911) );
  NAND2_X1 U1010 ( .A1(G115), .A2(n909), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1012 ( .A(KEYINPUT47), .B(n912), .Z(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n936) );
  XNOR2_X1 U1014 ( .A(n936), .B(n915), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n916), .B(G162), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(n918), .B(n917), .ZN(n921) );
  XNOR2_X1 U1017 ( .A(n919), .B(G164), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1019 ( .A(n923), .B(n922), .Z(n924) );
  NOR2_X1 U1020 ( .A1(G37), .A2(n924), .ZN(G395) );
  XOR2_X1 U1021 ( .A(n925), .B(G286), .Z(n927) );
  XNOR2_X1 U1022 ( .A(G171), .B(n987), .ZN(n926) );
  XNOR2_X1 U1023 ( .A(n927), .B(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n928), .B(n982), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(G37), .A2(n929), .ZN(G397) );
  NAND2_X1 U1026 ( .A1(G319), .A2(n930), .ZN(n933) );
  NOR2_X1 U1027 ( .A1(G229), .A2(G227), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(KEYINPUT49), .B(n931), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1034 ( .A(G2072), .B(n936), .Z(n938) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1037 ( .A(KEYINPUT50), .B(n939), .Z(n957) );
  XOR2_X1 U1038 ( .A(G2084), .B(G160), .Z(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n945) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n950) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(n948), .B(KEYINPUT51), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n952) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT123), .B(n955), .ZN(n956) );
  NOR2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1050 ( .A(KEYINPUT52), .B(n958), .ZN(n959) );
  INV_X1 U1051 ( .A(KEYINPUT55), .ZN(n978) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n978), .ZN(n960) );
  NAND2_X1 U1053 ( .A1(n960), .A2(G29), .ZN(n1037) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G35), .ZN(n973) );
  XOR2_X1 U1055 ( .A(G1991), .B(G25), .Z(n961) );
  NAND2_X1 U1056 ( .A1(n961), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1057 ( .A(G2067), .B(G26), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G33), .B(G2072), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n968) );
  XOR2_X1 U1060 ( .A(n964), .B(G27), .Z(n966) );
  XNOR2_X1 U1061 ( .A(G1996), .B(G32), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1067 ( .A(G2084), .B(G34), .Z(n974) );
  XNOR2_X1 U1068 ( .A(KEYINPUT54), .B(n974), .ZN(n975) );
  NAND2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n978), .B(n977), .ZN(n980) );
  INV_X1 U1071 ( .A(G29), .ZN(n979) );
  NAND2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n981), .ZN(n1035) );
  XNOR2_X1 U1074 ( .A(G16), .B(KEYINPUT56), .ZN(n1006) );
  XNOR2_X1 U1075 ( .A(G171), .B(G1961), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(n982), .B(G1341), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(G299), .B(G1956), .ZN(n983) );
  NOR2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n990) );
  XOR2_X1 U1080 ( .A(G1348), .B(n987), .Z(n988) );
  XNOR2_X1 U1081 ( .A(KEYINPUT124), .B(n988), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n1004) );
  XOR2_X1 U1083 ( .A(G168), .B(G1966), .Z(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1085 ( .A(KEYINPUT57), .B(n993), .Z(n1000) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n997) );
  AND2_X1 U1087 ( .A1(G303), .A2(G1971), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT125), .B(n998), .Z(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(n1005), .ZN(n1033) );
  INV_X1 U1094 ( .A(G16), .ZN(n1031) );
  XNOR2_X1 U1095 ( .A(n1007), .B(G5), .ZN(n1027) );
  XOR2_X1 U1096 ( .A(G1966), .B(G21), .Z(n1018) );
  XNOR2_X1 U1097 ( .A(G1348), .B(KEYINPUT59), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(G4), .ZN(n1012) );
  XNOR2_X1 U1099 ( .A(G1956), .B(G20), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G6), .B(G1981), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT126), .B(G1341), .ZN(n1013) );
  XNOR2_X1 U1104 ( .A(G19), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT60), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1025) );
  XNOR2_X1 U1108 ( .A(G1986), .B(G24), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(G1971), .B(G22), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XOR2_X1 U1111 ( .A(G1976), .B(G23), .Z(n1021) );
  NAND2_X1 U1112 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1113 ( .A(KEYINPUT58), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1114 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1116 ( .A(n1028), .B(KEYINPUT61), .ZN(n1029) );
  XNOR2_X1 U1117 ( .A(KEYINPUT127), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NOR2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  NAND2_X1 U1121 ( .A1(n1037), .A2(n1036), .ZN(n1038) );
  XOR2_X1 U1122 ( .A(KEYINPUT62), .B(n1038), .Z(G311) );
  INV_X1 U1123 ( .A(G311), .ZN(G150) );
endmodule

