

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(n620), .A2(n527), .ZN(n638) );
  NOR2_X4 U549 ( .A1(n543), .A2(n542), .ZN(G160) );
  NOR2_X1 U550 ( .A1(G164), .A2(G1384), .ZN(n669) );
  BUF_X1 U551 ( .A(n549), .Z(n550) );
  AND2_X2 U552 ( .A1(n515), .A2(G2104), .ZN(n992) );
  XNOR2_X1 U553 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n513) );
  INV_X1 U554 ( .A(KEYINPUT101), .ZN(n752) );
  XNOR2_X1 U555 ( .A(n534), .B(KEYINPUT7), .ZN(n535) );
  OR2_X1 U556 ( .A1(n698), .A2(n697), .ZN(n511) );
  INV_X1 U557 ( .A(KEYINPUT27), .ZN(n674) );
  OR2_X1 U558 ( .A1(n702), .A2(n701), .ZN(n703) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n705) );
  INV_X1 U560 ( .A(KEYINPUT31), .ZN(n720) );
  INV_X1 U561 ( .A(n931), .ZN(n743) );
  NOR2_X1 U562 ( .A1(n760), .A2(n743), .ZN(n744) );
  INV_X1 U563 ( .A(n926), .ZN(n748) );
  OR2_X1 U564 ( .A1(n749), .A2(n748), .ZN(n750) );
  INV_X1 U565 ( .A(G2105), .ZN(n515) );
  NOR2_X2 U566 ( .A1(G2104), .A2(n515), .ZN(n988) );
  NOR2_X1 U567 ( .A1(G651), .A2(n620), .ZN(n635) );
  OR2_X1 U568 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U569 ( .A(n537), .B(n536), .ZN(n539) );
  AND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(G164) );
  NOR2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n512) );
  XNOR2_X1 U572 ( .A(n513), .B(n512), .ZN(n549) );
  NAND2_X1 U573 ( .A1(n549), .A2(G138), .ZN(n514) );
  XNOR2_X1 U574 ( .A(n514), .B(KEYINPUT86), .ZN(n521) );
  AND2_X1 U575 ( .A1(n988), .A2(G126), .ZN(n519) );
  NAND2_X1 U576 ( .A1(G102), .A2(n992), .ZN(n517) );
  AND2_X1 U577 ( .A1(G2105), .A2(G2104), .ZN(n989) );
  NAND2_X1 U578 ( .A1(G114), .A2(n989), .ZN(n516) );
  NAND2_X1 U579 ( .A1(n517), .A2(n516), .ZN(n518) );
  NOR2_X1 U580 ( .A1(n519), .A2(n518), .ZN(n520) );
  NOR2_X1 U581 ( .A1(G651), .A2(G543), .ZN(n634) );
  NAND2_X1 U582 ( .A1(n634), .A2(G89), .ZN(n522) );
  XNOR2_X1 U583 ( .A(KEYINPUT4), .B(n522), .ZN(n525) );
  XOR2_X1 U584 ( .A(G543), .B(KEYINPUT0), .Z(n620) );
  XNOR2_X1 U585 ( .A(KEYINPUT69), .B(G651), .ZN(n527) );
  NAND2_X1 U586 ( .A1(G76), .A2(n638), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT77), .B(n523), .Z(n524) );
  NAND2_X1 U588 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U589 ( .A(n526), .B(KEYINPUT5), .Z(n533) );
  NAND2_X1 U590 ( .A1(n635), .A2(G51), .ZN(n530) );
  NOR2_X1 U591 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X2 U592 ( .A(KEYINPUT1), .B(n528), .Z(n642) );
  NAND2_X1 U593 ( .A1(G63), .A2(n642), .ZN(n529) );
  NAND2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U595 ( .A(KEYINPUT6), .B(n531), .ZN(n532) );
  XNOR2_X1 U596 ( .A(KEYINPUT78), .B(n535), .ZN(G168) );
  XOR2_X1 U597 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U598 ( .A1(G101), .A2(n992), .ZN(n537) );
  XOR2_X1 U599 ( .A(KEYINPUT23), .B(KEYINPUT66), .Z(n536) );
  NAND2_X1 U600 ( .A1(n549), .A2(G137), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U602 ( .A1(G125), .A2(n988), .ZN(n541) );
  NAND2_X1 U603 ( .A1(G113), .A2(n989), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G99), .A2(n992), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G111), .A2(n989), .ZN(n544) );
  NAND2_X1 U607 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n988), .A2(G123), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT18), .B(n546), .Z(n547) );
  NOR2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n550), .A2(G135), .ZN(n551) );
  NAND2_X1 U612 ( .A1(n552), .A2(n551), .ZN(n980) );
  XNOR2_X1 U613 ( .A(G2096), .B(n980), .ZN(n553) );
  OR2_X1 U614 ( .A1(G2100), .A2(n553), .ZN(G156) );
  NAND2_X1 U615 ( .A1(n635), .A2(G53), .ZN(n555) );
  NAND2_X1 U616 ( .A1(G65), .A2(n642), .ZN(n554) );
  NAND2_X1 U617 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G91), .A2(n634), .ZN(n557) );
  NAND2_X1 U619 ( .A1(G78), .A2(n638), .ZN(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U621 ( .A1(n559), .A2(n558), .ZN(n933) );
  INV_X1 U622 ( .A(n933), .ZN(G299) );
  INV_X1 U623 ( .A(G132), .ZN(G219) );
  INV_X1 U624 ( .A(G82), .ZN(G220) );
  NAND2_X1 U625 ( .A1(G94), .A2(G452), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT72), .B(n560), .Z(G173) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT74), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT10), .B(n562), .Z(n829) );
  NAND2_X1 U630 ( .A1(n829), .A2(G567), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n563), .Z(G234) );
  NAND2_X1 U632 ( .A1(G81), .A2(n634), .ZN(n564) );
  XOR2_X1 U633 ( .A(KEYINPUT75), .B(n564), .Z(n565) );
  XNOR2_X1 U634 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U635 ( .A1(G68), .A2(n638), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U638 ( .A1(G43), .A2(n635), .ZN(n569) );
  NAND2_X1 U639 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n642), .A2(G56), .ZN(n571) );
  XOR2_X1 U641 ( .A(KEYINPUT14), .B(n571), .Z(n572) );
  NOR2_X2 U642 ( .A1(n573), .A2(n572), .ZN(n1005) );
  NAND2_X1 U643 ( .A1(n1005), .A2(G860), .ZN(G153) );
  NAND2_X1 U644 ( .A1(G77), .A2(n638), .ZN(n574) );
  XNOR2_X1 U645 ( .A(n574), .B(KEYINPUT70), .ZN(n576) );
  NAND2_X1 U646 ( .A1(G90), .A2(n634), .ZN(n575) );
  NAND2_X1 U647 ( .A1(n576), .A2(n575), .ZN(n578) );
  XOR2_X1 U648 ( .A(KEYINPUT71), .B(KEYINPUT9), .Z(n577) );
  XNOR2_X1 U649 ( .A(n578), .B(n577), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n642), .A2(G64), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n635), .A2(G52), .ZN(n579) );
  AND2_X1 U652 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U653 ( .A1(n582), .A2(n581), .ZN(G301) );
  NAND2_X1 U654 ( .A1(n634), .A2(G92), .ZN(n584) );
  NAND2_X1 U655 ( .A1(G66), .A2(n642), .ZN(n583) );
  NAND2_X1 U656 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n635), .A2(G54), .ZN(n586) );
  NAND2_X1 U658 ( .A1(G79), .A2(n638), .ZN(n585) );
  NAND2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n595) );
  XNOR2_X1 U661 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n594) );
  XNOR2_X1 U662 ( .A(n595), .B(n594), .ZN(n698) );
  NOR2_X1 U663 ( .A1(n698), .A2(G868), .ZN(n590) );
  INV_X1 U664 ( .A(G868), .ZN(n654) );
  NOR2_X1 U665 ( .A1(n654), .A2(G301), .ZN(n589) );
  NOR2_X1 U666 ( .A1(n590), .A2(n589), .ZN(G284) );
  XOR2_X1 U667 ( .A(KEYINPUT79), .B(n654), .Z(n591) );
  NOR2_X1 U668 ( .A1(G286), .A2(n591), .ZN(n593) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n592) );
  NOR2_X1 U670 ( .A1(n593), .A2(n592), .ZN(G297) );
  INV_X1 U671 ( .A(G860), .ZN(n610) );
  NAND2_X1 U672 ( .A1(n610), .A2(G559), .ZN(n596) );
  XOR2_X1 U673 ( .A(n595), .B(n594), .Z(n1006) );
  NAND2_X1 U674 ( .A1(n596), .A2(n1006), .ZN(n597) );
  XNOR2_X1 U675 ( .A(n597), .B(KEYINPUT80), .ZN(n598) );
  XNOR2_X1 U676 ( .A(KEYINPUT16), .B(n598), .ZN(G148) );
  NOR2_X1 U677 ( .A1(G559), .A2(n654), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n599), .A2(n1006), .ZN(n600) );
  XNOR2_X1 U679 ( .A(n600), .B(KEYINPUT81), .ZN(n602) );
  AND2_X1 U680 ( .A1(n1005), .A2(n654), .ZN(n601) );
  NOR2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G282) );
  NAND2_X1 U682 ( .A1(n634), .A2(G93), .ZN(n604) );
  NAND2_X1 U683 ( .A1(G67), .A2(n642), .ZN(n603) );
  NAND2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n635), .A2(G55), .ZN(n606) );
  NAND2_X1 U686 ( .A1(G80), .A2(n638), .ZN(n605) );
  NAND2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n607) );
  OR2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n653) );
  XNOR2_X1 U689 ( .A(n653), .B(KEYINPUT82), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n1006), .A2(G559), .ZN(n609) );
  XNOR2_X1 U691 ( .A(n609), .B(n1005), .ZN(n651) );
  NAND2_X1 U692 ( .A1(n651), .A2(n610), .ZN(n611) );
  XNOR2_X1 U693 ( .A(n612), .B(n611), .ZN(G145) );
  NAND2_X1 U694 ( .A1(G88), .A2(n634), .ZN(n614) );
  NAND2_X1 U695 ( .A1(G50), .A2(n635), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n642), .A2(G62), .ZN(n615) );
  XOR2_X1 U698 ( .A(KEYINPUT84), .B(n615), .Z(n616) );
  NOR2_X1 U699 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G75), .A2(n638), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(G303) );
  NAND2_X1 U702 ( .A1(G49), .A2(n635), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G87), .A2(n620), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n642), .A2(n623), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n624) );
  XOR2_X1 U707 ( .A(KEYINPUT83), .B(n624), .Z(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G60), .A2(n642), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G72), .A2(n638), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n634), .A2(G85), .ZN(n629) );
  XOR2_X1 U713 ( .A(KEYINPUT68), .B(n629), .Z(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n635), .A2(G47), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G86), .A2(n634), .ZN(n637) );
  NAND2_X1 U718 ( .A1(G48), .A2(n635), .ZN(n636) );
  NAND2_X1 U719 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n638), .A2(G73), .ZN(n639) );
  XOR2_X1 U721 ( .A(KEYINPUT2), .B(n639), .Z(n640) );
  NOR2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U723 ( .A1(G61), .A2(n642), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(G305) );
  XOR2_X1 U725 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n645) );
  XNOR2_X1 U726 ( .A(G288), .B(n645), .ZN(n646) );
  XOR2_X1 U727 ( .A(n653), .B(n646), .Z(n648) );
  XOR2_X1 U728 ( .A(G290), .B(G299), .Z(n647) );
  XNOR2_X1 U729 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U730 ( .A(n649), .B(G305), .Z(n650) );
  XOR2_X1 U731 ( .A(G303), .B(n650), .Z(n1008) );
  XNOR2_X1 U732 ( .A(n651), .B(n1008), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n652), .A2(G868), .ZN(n656) );
  NAND2_X1 U734 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n656), .A2(n655), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U743 ( .A1(G120), .A2(G108), .ZN(n661) );
  NOR2_X1 U744 ( .A1(G237), .A2(n661), .ZN(n662) );
  NAND2_X1 U745 ( .A1(G69), .A2(n662), .ZN(n956) );
  NAND2_X1 U746 ( .A1(n956), .A2(G567), .ZN(n667) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n663) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n663), .Z(n664) );
  NOR2_X1 U749 ( .A1(G218), .A2(n664), .ZN(n665) );
  NAND2_X1 U750 ( .A1(G96), .A2(n665), .ZN(n955) );
  NAND2_X1 U751 ( .A1(n955), .A2(G2106), .ZN(n666) );
  NAND2_X1 U752 ( .A1(n667), .A2(n666), .ZN(n976) );
  NAND2_X1 U753 ( .A1(G483), .A2(G661), .ZN(n668) );
  NOR2_X1 U754 ( .A1(n976), .A2(n668), .ZN(n831) );
  NAND2_X1 U755 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U756 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U757 ( .A(n669), .B(KEYINPUT64), .ZN(n767) );
  INV_X1 U758 ( .A(KEYINPUT94), .ZN(n670) );
  NAND2_X1 U759 ( .A1(G160), .A2(G40), .ZN(n768) );
  XNOR2_X1 U760 ( .A(n670), .B(n768), .ZN(n671) );
  NAND2_X1 U761 ( .A1(n767), .A2(n671), .ZN(n672) );
  BUF_X1 U762 ( .A(n672), .Z(n714) );
  NAND2_X1 U763 ( .A1(n714), .A2(G1956), .ZN(n677) );
  INV_X1 U764 ( .A(n672), .ZN(n673) );
  NAND2_X1 U765 ( .A1(n673), .A2(G2072), .ZN(n675) );
  XNOR2_X1 U766 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U768 ( .A(n678), .B(KEYINPUT97), .ZN(n699) );
  NOR2_X1 U769 ( .A1(n699), .A2(n933), .ZN(n680) );
  INV_X1 U770 ( .A(KEYINPUT28), .ZN(n679) );
  XNOR2_X1 U771 ( .A(n680), .B(n679), .ZN(n704) );
  INV_X1 U772 ( .A(G1341), .ZN(n942) );
  NAND2_X1 U773 ( .A1(n698), .A2(G1348), .ZN(n681) );
  NAND2_X1 U774 ( .A1(n942), .A2(n681), .ZN(n682) );
  NAND2_X1 U775 ( .A1(n714), .A2(n682), .ZN(n686) );
  INV_X1 U776 ( .A(n714), .ZN(n694) );
  NAND2_X1 U777 ( .A1(n694), .A2(G1996), .ZN(n684) );
  XOR2_X1 U778 ( .A(KEYINPUT65), .B(KEYINPUT26), .Z(n687) );
  INV_X1 U779 ( .A(n687), .ZN(n683) );
  NAND2_X1 U780 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n686), .A2(n685), .ZN(n693) );
  NAND2_X1 U782 ( .A1(n698), .A2(G2067), .ZN(n689) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n687), .ZN(n688) );
  NAND2_X1 U784 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U785 ( .A1(n690), .A2(n694), .ZN(n691) );
  NAND2_X1 U786 ( .A1(n1005), .A2(n691), .ZN(n692) );
  NOR2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n702) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n714), .ZN(n696) );
  NAND2_X1 U789 ( .A1(G2067), .A2(n694), .ZN(n695) );
  NAND2_X1 U790 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n699), .A2(n933), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n511), .A2(n700), .ZN(n701) );
  NAND2_X1 U793 ( .A1(n704), .A2(n703), .ZN(n706) );
  XNOR2_X1 U794 ( .A(n706), .B(n705), .ZN(n711) );
  XNOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .ZN(n851) );
  NOR2_X1 U796 ( .A1(n714), .A2(n851), .ZN(n708) );
  AND2_X1 U797 ( .A1(n714), .A2(G1961), .ZN(n707) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n713) );
  AND2_X1 U799 ( .A1(G171), .A2(n713), .ZN(n709) );
  XOR2_X1 U800 ( .A(KEYINPUT96), .B(n709), .Z(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U802 ( .A(n712), .B(KEYINPUT98), .ZN(n723) );
  NOR2_X1 U803 ( .A1(G171), .A2(n713), .ZN(n719) );
  NAND2_X1 U804 ( .A1(G8), .A2(n714), .ZN(n760) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n760), .ZN(n737) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n714), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n737), .A2(n732), .ZN(n715) );
  NAND2_X1 U808 ( .A1(G8), .A2(n715), .ZN(n716) );
  XNOR2_X1 U809 ( .A(KEYINPUT30), .B(n716), .ZN(n717) );
  NOR2_X1 U810 ( .A1(n717), .A2(G168), .ZN(n718) );
  NOR2_X1 U811 ( .A1(n719), .A2(n718), .ZN(n721) );
  XNOR2_X1 U812 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U813 ( .A1(n723), .A2(n722), .ZN(n734) );
  NAND2_X1 U814 ( .A1(n734), .A2(G286), .ZN(n728) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n760), .ZN(n725) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n714), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n726), .A2(G303), .ZN(n727) );
  NAND2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U820 ( .A(n729), .B(KEYINPUT100), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n730), .A2(G8), .ZN(n731) );
  XNOR2_X1 U822 ( .A(n731), .B(KEYINPUT32), .ZN(n740) );
  NAND2_X1 U823 ( .A1(G8), .A2(n732), .ZN(n733) );
  XOR2_X1 U824 ( .A(KEYINPUT95), .B(n733), .Z(n735) );
  NAND2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n736) );
  NOR2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U827 ( .A(KEYINPUT99), .B(n738), .ZN(n739) );
  NAND2_X1 U828 ( .A1(n740), .A2(n739), .ZN(n756) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n930) );
  NOR2_X1 U830 ( .A1(G1971), .A2(G303), .ZN(n741) );
  NOR2_X1 U831 ( .A1(n930), .A2(n741), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n756), .A2(n742), .ZN(n745) );
  NAND2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n931) );
  AND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U835 ( .A1(KEYINPUT33), .A2(n746), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n930), .A2(KEYINPUT33), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n747), .A2(n760), .ZN(n749) );
  XOR2_X1 U838 ( .A(G1981), .B(G305), .Z(n926) );
  NOR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n753) );
  XNOR2_X1 U840 ( .A(n753), .B(n752), .ZN(n764) );
  NOR2_X1 U841 ( .A1(G1981), .A2(G305), .ZN(n754) );
  XOR2_X1 U842 ( .A(n754), .B(KEYINPUT24), .Z(n755) );
  OR2_X1 U843 ( .A1(n760), .A2(n755), .ZN(n762) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n757) );
  NAND2_X1 U845 ( .A1(G8), .A2(n757), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n756), .A2(n758), .ZN(n759) );
  NAND2_X1 U847 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n762), .A2(n761), .ZN(n763) );
  NOR2_X1 U849 ( .A1(n764), .A2(n763), .ZN(n766) );
  INV_X1 U850 ( .A(KEYINPUT102), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n766), .B(n765), .ZN(n803) );
  NOR2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n814) );
  NAND2_X1 U853 ( .A1(n989), .A2(G116), .ZN(n769) );
  XNOR2_X1 U854 ( .A(KEYINPUT88), .B(n769), .ZN(n772) );
  NAND2_X1 U855 ( .A1(n988), .A2(G128), .ZN(n770) );
  XOR2_X1 U856 ( .A(KEYINPUT87), .B(n770), .Z(n771) );
  NAND2_X1 U857 ( .A1(n772), .A2(n771), .ZN(n773) );
  XNOR2_X1 U858 ( .A(n773), .B(KEYINPUT35), .ZN(n778) );
  NAND2_X1 U859 ( .A1(G104), .A2(n992), .ZN(n775) );
  NAND2_X1 U860 ( .A1(G140), .A2(n550), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U862 ( .A(KEYINPUT34), .B(n776), .Z(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U864 ( .A(n779), .B(KEYINPUT36), .Z(n1001) );
  XNOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .ZN(n812) );
  NOR2_X1 U866 ( .A1(n1001), .A2(n812), .ZN(n890) );
  AND2_X1 U867 ( .A1(n814), .A2(n890), .ZN(n810) );
  NAND2_X1 U868 ( .A1(G119), .A2(n988), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G107), .A2(n989), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT89), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G95), .A2(n992), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n550), .A2(G131), .ZN(n785) );
  XOR2_X1 U875 ( .A(KEYINPUT90), .B(n785), .Z(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U877 ( .A(KEYINPUT91), .B(n788), .ZN(n985) );
  AND2_X1 U878 ( .A1(n985), .A2(G1991), .ZN(n797) );
  NAND2_X1 U879 ( .A1(G129), .A2(n988), .ZN(n790) );
  NAND2_X1 U880 ( .A1(G141), .A2(n550), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U882 ( .A1(n992), .A2(G105), .ZN(n791) );
  XOR2_X1 U883 ( .A(KEYINPUT38), .B(n791), .Z(n792) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U885 ( .A1(n989), .A2(G117), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n981) );
  AND2_X1 U887 ( .A1(n981), .A2(G1996), .ZN(n796) );
  NOR2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n900) );
  XOR2_X1 U889 ( .A(n814), .B(KEYINPUT92), .Z(n798) );
  NOR2_X1 U890 ( .A1(n900), .A2(n798), .ZN(n806) );
  OR2_X1 U891 ( .A1(n810), .A2(n806), .ZN(n799) );
  XOR2_X1 U892 ( .A(KEYINPUT93), .B(n799), .Z(n801) );
  XNOR2_X1 U893 ( .A(G1986), .B(G290), .ZN(n939) );
  AND2_X1 U894 ( .A1(n939), .A2(n814), .ZN(n800) );
  NOR2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n817) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n981), .ZN(n894) );
  NOR2_X1 U898 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U899 ( .A1(G1991), .A2(n985), .ZN(n898) );
  NOR2_X1 U900 ( .A1(n804), .A2(n898), .ZN(n805) );
  NOR2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n894), .A2(n807), .ZN(n808) );
  XOR2_X1 U903 ( .A(KEYINPUT39), .B(n808), .Z(n809) );
  NOR2_X1 U904 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U905 ( .A(n811), .B(KEYINPUT103), .ZN(n813) );
  NAND2_X1 U906 ( .A1(n1001), .A2(n812), .ZN(n892) );
  NAND2_X1 U907 ( .A1(n813), .A2(n892), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(n818), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U911 ( .A(G2443), .B(G1348), .ZN(n827) );
  XNOR2_X1 U912 ( .A(G2430), .B(G2446), .ZN(n825) );
  XOR2_X1 U913 ( .A(G2454), .B(G2451), .Z(n820) );
  XNOR2_X1 U914 ( .A(G2427), .B(G2435), .ZN(n819) );
  XNOR2_X1 U915 ( .A(n820), .B(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(n821), .B(G2438), .Z(n823) );
  XOR2_X1 U917 ( .A(n942), .B(KEYINPUT104), .Z(n822) );
  XNOR2_X1 U918 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n827), .B(n826), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(G14), .ZN(n1014) );
  XNOR2_X1 U922 ( .A(KEYINPUT105), .B(n1014), .ZN(G401) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n829), .ZN(G217) );
  INV_X1 U924 ( .A(n829), .ZN(G223) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U926 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G1), .A2(G3), .ZN(n832) );
  NAND2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT106), .ZN(G188) );
  XNOR2_X1 U930 ( .A(G108), .B(KEYINPUT117), .ZN(G238) );
  NAND2_X1 U932 ( .A1(G100), .A2(n992), .ZN(n835) );
  NAND2_X1 U933 ( .A1(G112), .A2(n989), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n836), .B(KEYINPUT109), .ZN(n838) );
  NAND2_X1 U936 ( .A1(G136), .A2(n550), .ZN(n837) );
  NAND2_X1 U937 ( .A1(n838), .A2(n837), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n988), .A2(G124), .ZN(n839) );
  XOR2_X1 U939 ( .A(KEYINPUT44), .B(n839), .Z(n840) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G162) );
  XOR2_X1 U941 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n920) );
  XNOR2_X1 U942 ( .A(G2090), .B(G35), .ZN(n856) );
  XNOR2_X1 U943 ( .A(KEYINPUT119), .B(G2067), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n842), .B(G26), .ZN(n850) );
  XNOR2_X1 U945 ( .A(G1991), .B(G25), .ZN(n844) );
  XNOR2_X1 U946 ( .A(G33), .B(G2072), .ZN(n843) );
  NOR2_X1 U947 ( .A1(n844), .A2(n843), .ZN(n845) );
  NAND2_X1 U948 ( .A1(G28), .A2(n845), .ZN(n848) );
  XNOR2_X1 U949 ( .A(G32), .B(G1996), .ZN(n846) );
  XNOR2_X1 U950 ( .A(KEYINPUT120), .B(n846), .ZN(n847) );
  NOR2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n849) );
  NAND2_X1 U952 ( .A1(n850), .A2(n849), .ZN(n853) );
  XOR2_X1 U953 ( .A(G27), .B(n851), .Z(n852) );
  NOR2_X1 U954 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U955 ( .A(KEYINPUT53), .B(n854), .ZN(n855) );
  NOR2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n859) );
  XOR2_X1 U957 ( .A(G2084), .B(G34), .Z(n857) );
  XNOR2_X1 U958 ( .A(KEYINPUT54), .B(n857), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n920), .B(n860), .ZN(n862) );
  INV_X1 U961 ( .A(G29), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G11), .A2(n863), .ZN(n889) );
  XNOR2_X1 U964 ( .A(G21), .B(G1966), .ZN(n864) );
  XNOR2_X1 U965 ( .A(n864), .B(KEYINPUT125), .ZN(n877) );
  XOR2_X1 U966 ( .A(G1956), .B(G20), .Z(n869) );
  XOR2_X1 U967 ( .A(n942), .B(G19), .Z(n866) );
  XNOR2_X1 U968 ( .A(G6), .B(G1981), .ZN(n865) );
  NOR2_X1 U969 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(KEYINPUT124), .B(n867), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n872) );
  XOR2_X1 U972 ( .A(KEYINPUT59), .B(G1348), .Z(n870) );
  XNOR2_X1 U973 ( .A(G4), .B(n870), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U975 ( .A(KEYINPUT60), .B(n873), .Z(n875) );
  XNOR2_X1 U976 ( .A(G1961), .B(G5), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  NAND2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n884) );
  XNOR2_X1 U979 ( .A(G1971), .B(G22), .ZN(n879) );
  XNOR2_X1 U980 ( .A(G23), .B(G1976), .ZN(n878) );
  NOR2_X1 U981 ( .A1(n879), .A2(n878), .ZN(n881) );
  XOR2_X1 U982 ( .A(G1986), .B(G24), .Z(n880) );
  NAND2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U984 ( .A(KEYINPUT58), .B(n882), .ZN(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U986 ( .A(KEYINPUT61), .B(n885), .Z(n886) );
  NOR2_X1 U987 ( .A1(G16), .A2(n886), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT126), .ZN(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n924) );
  INV_X1 U990 ( .A(n890), .ZN(n891) );
  NAND2_X1 U991 ( .A1(n892), .A2(n891), .ZN(n918) );
  XOR2_X1 U992 ( .A(G2090), .B(G162), .Z(n893) );
  NOR2_X1 U993 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(KEYINPUT51), .B(n895), .Z(n916) );
  XNOR2_X1 U995 ( .A(G160), .B(G2084), .ZN(n896) );
  NAND2_X1 U996 ( .A1(n896), .A2(n980), .ZN(n897) );
  NOR2_X1 U997 ( .A1(n898), .A2(n897), .ZN(n899) );
  NAND2_X1 U998 ( .A1(n900), .A2(n899), .ZN(n914) );
  NAND2_X1 U999 ( .A1(n989), .A2(G115), .ZN(n901) );
  XOR2_X1 U1000 ( .A(KEYINPUT111), .B(n901), .Z(n903) );
  NAND2_X1 U1001 ( .A1(n988), .A2(G127), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n904), .B(KEYINPUT47), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n992), .ZN(n905) );
  NAND2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n909) );
  NAND2_X1 U1006 ( .A1(n550), .A2(G139), .ZN(n907) );
  XOR2_X1 U1007 ( .A(KEYINPUT110), .B(n907), .Z(n908) );
  NOR2_X1 U1008 ( .A1(n909), .A2(n908), .ZN(n1000) );
  XOR2_X1 U1009 ( .A(G2072), .B(n1000), .Z(n911) );
  XOR2_X1 U1010 ( .A(G164), .B(G2078), .Z(n910) );
  NOR2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1012 ( .A(KEYINPUT50), .B(n912), .Z(n913) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT52), .B(n919), .ZN(n921) );
  NAND2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(n922), .A2(G29), .ZN(n923) );
  NAND2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n953) );
  XOR2_X1 U1020 ( .A(G16), .B(KEYINPUT56), .Z(n951) );
  XOR2_X1 U1021 ( .A(G1966), .B(KEYINPUT121), .Z(n925) );
  XNOR2_X1 U1022 ( .A(G168), .B(n925), .ZN(n927) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(n928), .B(KEYINPUT57), .ZN(n941) );
  XOR2_X1 U1025 ( .A(G1971), .B(G303), .Z(n929) );
  XNOR2_X1 U1026 ( .A(n929), .B(KEYINPUT122), .ZN(n937) );
  INV_X1 U1027 ( .A(n930), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1029 ( .A(G1956), .B(n933), .Z(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n948) );
  XOR2_X1 U1034 ( .A(G301), .B(G1961), .Z(n946) );
  XNOR2_X1 U1035 ( .A(n1005), .B(n942), .ZN(n944) );
  XOR2_X1 U1036 ( .A(n1006), .B(G1348), .Z(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1039 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1040 ( .A(KEYINPUT123), .B(n949), .Z(n950) );
  NOR2_X1 U1041 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1042 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(n954), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1044 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1045 ( .A(G120), .ZN(G236) );
  INV_X1 U1046 ( .A(G96), .ZN(G221) );
  INV_X1 U1047 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1048 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1049 ( .A(n957), .B(KEYINPUT107), .Z(G325) );
  INV_X1 U1050 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1051 ( .A(G2100), .B(G2096), .Z(n959) );
  XNOR2_X1 U1052 ( .A(G2072), .B(G2090), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n959), .B(n958), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2678), .B(KEYINPUT42), .Z(n961) );
  XNOR2_X1 U1055 ( .A(G2067), .B(KEYINPUT43), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n961), .B(n960), .ZN(n962) );
  XOR2_X1 U1057 ( .A(n963), .B(n962), .Z(n965) );
  XNOR2_X1 U1058 ( .A(G2084), .B(G2078), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n965), .B(n964), .ZN(G227) );
  XNOR2_X1 U1060 ( .A(G1976), .B(KEYINPUT41), .ZN(n975) );
  XOR2_X1 U1061 ( .A(G1981), .B(G1971), .Z(n967) );
  XNOR2_X1 U1062 ( .A(G1986), .B(G1956), .ZN(n966) );
  XNOR2_X1 U1063 ( .A(n967), .B(n966), .ZN(n971) );
  XOR2_X1 U1064 ( .A(G2474), .B(KEYINPUT108), .Z(n969) );
  XNOR2_X1 U1065 ( .A(G1996), .B(G1991), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(n969), .B(n968), .ZN(n970) );
  XOR2_X1 U1067 ( .A(n971), .B(n970), .Z(n973) );
  XNOR2_X1 U1068 ( .A(G1966), .B(G1961), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(n973), .B(n972), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n975), .B(n974), .ZN(G229) );
  INV_X1 U1071 ( .A(n976), .ZN(G319) );
  XOR2_X1 U1072 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n978), .B(n977), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(n980), .B(n979), .ZN(n983) );
  XOR2_X1 U1076 ( .A(G160), .B(n981), .Z(n982) );
  XNOR2_X1 U1077 ( .A(n983), .B(n982), .ZN(n984) );
  XOR2_X1 U1078 ( .A(n984), .B(G162), .Z(n987) );
  XOR2_X1 U1079 ( .A(G164), .B(n985), .Z(n986) );
  XNOR2_X1 U1080 ( .A(n987), .B(n986), .ZN(n999) );
  NAND2_X1 U1081 ( .A1(G130), .A2(n988), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(G118), .A2(n989), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n997) );
  NAND2_X1 U1084 ( .A1(G106), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(G142), .A2(n550), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1087 ( .A(KEYINPUT45), .B(n995), .Z(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(n999), .B(n998), .Z(n1003) );
  XOR2_X1 U1090 ( .A(n1001), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(n1003), .B(n1002), .ZN(n1004) );
  NOR2_X1 U1092 ( .A1(G37), .A2(n1004), .ZN(G395) );
  XNOR2_X1 U1093 ( .A(n1006), .B(n1005), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G286), .B(n1007), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G301), .B(n1008), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(n1010), .B(n1009), .ZN(n1011) );
  NOR2_X1 U1097 ( .A1(G37), .A2(n1011), .ZN(G397) );
  XNOR2_X1 U1098 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n1013) );
  NOR2_X1 U1099 ( .A1(G227), .A2(G229), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(n1013), .B(n1012), .ZN(n1016) );
  NAND2_X1 U1101 ( .A1(G319), .A2(n1014), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1103 ( .A(KEYINPUT115), .B(n1017), .Z(n1020) );
  NOR2_X1 U1104 ( .A1(G395), .A2(G397), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(KEYINPUT116), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(G225) );
  INV_X1 U1107 ( .A(G225), .ZN(G308) );
  INV_X1 U1108 ( .A(G303), .ZN(G166) );
endmodule

