

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U550 ( .A1(n555), .A2(G2105), .ZN(n679) );
  AND2_X2 U551 ( .A1(n547), .A2(G2104), .ZN(n893) );
  INV_X1 U552 ( .A(KEYINPUT105), .ZN(n782) );
  INV_X1 U553 ( .A(KEYINPUT17), .ZN(n553) );
  OR2_X1 U554 ( .A1(n733), .A2(G171), .ZN(n516) );
  XNOR2_X1 U555 ( .A(n735), .B(KEYINPUT31), .ZN(n747) );
  AND2_X1 U556 ( .A1(n896), .A2(G114), .ZN(n517) );
  XOR2_X1 U557 ( .A(n715), .B(KEYINPUT28), .Z(n518) );
  NOR2_X1 U558 ( .A1(n939), .A2(n714), .ZN(n715) );
  INV_X1 U559 ( .A(G168), .ZN(n731) );
  BUF_X1 U560 ( .A(n704), .Z(n721) );
  NAND2_X1 U561 ( .A1(n734), .A2(n516), .ZN(n735) );
  AND2_X1 U562 ( .A1(n747), .A2(n741), .ZN(n740) );
  AND2_X1 U563 ( .A1(n766), .A2(n765), .ZN(n767) );
  INV_X1 U564 ( .A(G2104), .ZN(n555) );
  INV_X1 U565 ( .A(G2105), .ZN(n547) );
  NOR2_X2 U566 ( .A1(n523), .A2(n524), .ZN(n636) );
  XNOR2_X1 U567 ( .A(n572), .B(KEYINPUT77), .ZN(n693) );
  INV_X1 U568 ( .A(n693), .ZN(n933) );
  NOR2_X1 U569 ( .A1(G543), .A2(G651), .ZN(n635) );
  NAND2_X1 U570 ( .A1(n635), .A2(G89), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n519), .B(KEYINPUT4), .ZN(n521) );
  XOR2_X1 U572 ( .A(G543), .B(KEYINPUT0), .Z(n523) );
  INV_X1 U573 ( .A(G651), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G76), .A2(n636), .ZN(n520) );
  NAND2_X1 U575 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U576 ( .A(n522), .B(KEYINPUT5), .ZN(n530) );
  NOR2_X2 U577 ( .A1(G651), .A2(n523), .ZN(n643) );
  NAND2_X1 U578 ( .A1(G51), .A2(n643), .ZN(n527) );
  NOR2_X1 U579 ( .A1(G543), .A2(n524), .ZN(n525) );
  XOR2_X2 U580 ( .A(KEYINPUT1), .B(n525), .Z(n639) );
  NAND2_X1 U581 ( .A1(G63), .A2(n639), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT6), .B(n528), .Z(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n531), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U586 ( .A1(G52), .A2(n643), .ZN(n533) );
  NAND2_X1 U587 ( .A1(G64), .A2(n639), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n533), .A2(n532), .ZN(n539) );
  NAND2_X1 U589 ( .A1(G90), .A2(n635), .ZN(n535) );
  NAND2_X1 U590 ( .A1(G77), .A2(n636), .ZN(n534) );
  NAND2_X1 U591 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U592 ( .A(KEYINPUT67), .B(n536), .ZN(n537) );
  XNOR2_X1 U593 ( .A(KEYINPUT9), .B(n537), .ZN(n538) );
  NOR2_X1 U594 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U595 ( .A(KEYINPUT68), .B(n540), .Z(G301) );
  INV_X1 U596 ( .A(G301), .ZN(G171) );
  NAND2_X1 U597 ( .A1(G85), .A2(n635), .ZN(n542) );
  NAND2_X1 U598 ( .A1(G72), .A2(n636), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U600 ( .A1(G47), .A2(n643), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G60), .A2(n639), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U603 ( .A1(n546), .A2(n545), .ZN(G290) );
  NAND2_X1 U604 ( .A1(G101), .A2(n893), .ZN(n548) );
  XNOR2_X1 U605 ( .A(n548), .B(KEYINPUT23), .ZN(n549) );
  XNOR2_X1 U606 ( .A(KEYINPUT65), .B(n549), .ZN(n552) );
  AND2_X1 U607 ( .A1(G2105), .A2(G2104), .ZN(n896) );
  NAND2_X1 U608 ( .A1(G113), .A2(n896), .ZN(n550) );
  XNOR2_X1 U609 ( .A(n550), .B(KEYINPUT66), .ZN(n551) );
  AND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n685) );
  NOR2_X1 U611 ( .A1(G2105), .A2(G2104), .ZN(n554) );
  XNOR2_X1 U612 ( .A(n554), .B(n553), .ZN(n675) );
  BUF_X1 U613 ( .A(n675), .Z(n606) );
  NAND2_X1 U614 ( .A1(G137), .A2(n606), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G125), .A2(n679), .ZN(n556) );
  AND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n684) );
  AND2_X1 U617 ( .A1(n685), .A2(n684), .ZN(G160) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U619 ( .A1(G94), .A2(G452), .ZN(n558) );
  XNOR2_X1 U620 ( .A(n558), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U622 ( .A(n559), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U623 ( .A(G223), .B(KEYINPUT74), .Z(n833) );
  NAND2_X1 U624 ( .A1(n833), .A2(G567), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U626 ( .A1(n636), .A2(G68), .ZN(n561) );
  XNOR2_X1 U627 ( .A(KEYINPUT76), .B(n561), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n635), .A2(G81), .ZN(n562) );
  XNOR2_X1 U629 ( .A(KEYINPUT12), .B(n562), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(KEYINPUT13), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G43), .A2(n643), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U634 ( .A1(G56), .A2(n639), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT14), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n569), .B(KEYINPUT75), .ZN(n570) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n933), .A2(G860), .ZN(G153) );
  NAND2_X1 U639 ( .A1(G92), .A2(n635), .ZN(n574) );
  NAND2_X1 U640 ( .A1(G79), .A2(n636), .ZN(n573) );
  NAND2_X1 U641 ( .A1(n574), .A2(n573), .ZN(n578) );
  NAND2_X1 U642 ( .A1(G54), .A2(n643), .ZN(n576) );
  NAND2_X1 U643 ( .A1(G66), .A2(n639), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(KEYINPUT15), .B(n579), .Z(n580) );
  XOR2_X1 U647 ( .A(KEYINPUT78), .B(n580), .Z(n596) );
  INV_X1 U648 ( .A(n596), .ZN(n927) );
  NOR2_X1 U649 ( .A1(G868), .A2(n927), .ZN(n581) );
  XNOR2_X1 U650 ( .A(n581), .B(KEYINPUT79), .ZN(n583) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U652 ( .A1(n583), .A2(n582), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G91), .A2(n635), .ZN(n585) );
  NAND2_X1 U654 ( .A1(G78), .A2(n636), .ZN(n584) );
  NAND2_X1 U655 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U656 ( .A(KEYINPUT70), .B(n586), .Z(n588) );
  NAND2_X1 U657 ( .A1(n639), .A2(G65), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U659 ( .A1(G53), .A2(n643), .ZN(n589) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n589), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n939) );
  XOR2_X1 U662 ( .A(n939), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U663 ( .A1(G299), .A2(G868), .ZN(n592) );
  XNOR2_X1 U664 ( .A(n592), .B(KEYINPUT80), .ZN(n594) );
  INV_X1 U665 ( .A(G868), .ZN(n600) );
  NOR2_X1 U666 ( .A1(n600), .A2(G286), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G297) );
  INV_X1 U668 ( .A(G559), .ZN(n598) );
  NOR2_X1 U669 ( .A1(G860), .A2(n598), .ZN(n595) );
  NOR2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U671 ( .A(KEYINPUT16), .B(n597), .Z(G148) );
  NAND2_X1 U672 ( .A1(n598), .A2(n927), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n599), .A2(G868), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n693), .A2(n600), .ZN(n601) );
  NAND2_X1 U675 ( .A1(n602), .A2(n601), .ZN(G282) );
  XNOR2_X1 U676 ( .A(G2100), .B(KEYINPUT81), .ZN(n612) );
  NAND2_X1 U677 ( .A1(G123), .A2(n679), .ZN(n603) );
  XNOR2_X1 U678 ( .A(n603), .B(KEYINPUT18), .ZN(n605) );
  NAND2_X1 U679 ( .A1(n893), .A2(G99), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n610) );
  NAND2_X1 U681 ( .A1(G135), .A2(n606), .ZN(n608) );
  NAND2_X1 U682 ( .A1(G111), .A2(n896), .ZN(n607) );
  NAND2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n988) );
  XNOR2_X1 U685 ( .A(n988), .B(G2096), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G559), .A2(n927), .ZN(n656) );
  XOR2_X1 U688 ( .A(n933), .B(n656), .Z(n613) );
  NOR2_X1 U689 ( .A1(G860), .A2(n613), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n643), .A2(G55), .ZN(n616) );
  NAND2_X1 U691 ( .A1(G80), .A2(n636), .ZN(n614) );
  XOR2_X1 U692 ( .A(KEYINPUT83), .B(n614), .Z(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U694 ( .A1(G93), .A2(n635), .ZN(n618) );
  NAND2_X1 U695 ( .A1(G67), .A2(n639), .ZN(n617) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n652) );
  XNOR2_X1 U698 ( .A(n652), .B(KEYINPUT82), .ZN(n621) );
  XNOR2_X1 U699 ( .A(n622), .B(n621), .ZN(G145) );
  NAND2_X1 U700 ( .A1(G49), .A2(n643), .ZN(n624) );
  NAND2_X1 U701 ( .A1(G74), .A2(G651), .ZN(n623) );
  NAND2_X1 U702 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U703 ( .A1(n639), .A2(n625), .ZN(n627) );
  NAND2_X1 U704 ( .A1(n523), .A2(G87), .ZN(n626) );
  NAND2_X1 U705 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G86), .A2(n635), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G48), .A2(n643), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n636), .A2(G73), .ZN(n630) );
  XOR2_X1 U710 ( .A(KEYINPUT2), .B(n630), .Z(n631) );
  NOR2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n639), .A2(G61), .ZN(n633) );
  NAND2_X1 U713 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U714 ( .A1(G88), .A2(n635), .ZN(n638) );
  NAND2_X1 U715 ( .A1(G75), .A2(n636), .ZN(n637) );
  NAND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n639), .A2(G62), .ZN(n640) );
  XOR2_X1 U718 ( .A(KEYINPUT84), .B(n640), .Z(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n643), .A2(G50), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(G303) );
  NOR2_X1 U722 ( .A1(G868), .A2(n652), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n646), .B(KEYINPUT87), .ZN(n659) );
  XOR2_X1 U724 ( .A(G290), .B(G305), .Z(n647) );
  XNOR2_X1 U725 ( .A(G288), .B(n647), .ZN(n648) );
  XOR2_X1 U726 ( .A(n648), .B(KEYINPUT86), .Z(n650) );
  XNOR2_X1 U727 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n649) );
  XNOR2_X1 U728 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U729 ( .A(n652), .B(n651), .Z(n654) );
  XOR2_X1 U730 ( .A(G303), .B(G299), .Z(n653) );
  XNOR2_X1 U731 ( .A(n654), .B(n653), .ZN(n655) );
  XNOR2_X1 U732 ( .A(n655), .B(n933), .ZN(n906) );
  XNOR2_X1 U733 ( .A(n906), .B(n656), .ZN(n657) );
  NAND2_X1 U734 ( .A1(G868), .A2(n657), .ZN(n658) );
  NAND2_X1 U735 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n660) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(KEYINPUT88), .B(KEYINPUT21), .ZN(n662) );
  XNOR2_X1 U740 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U741 ( .A1(n664), .A2(G2072), .ZN(n665) );
  XOR2_X1 U742 ( .A(KEYINPUT89), .B(n665), .Z(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U744 ( .A(KEYINPUT73), .B(G57), .ZN(G237) );
  NAND2_X1 U745 ( .A1(G132), .A2(G82), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n666), .B(KEYINPUT90), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(KEYINPUT22), .ZN(n668) );
  NOR2_X1 U748 ( .A1(G218), .A2(n668), .ZN(n669) );
  NAND2_X1 U749 ( .A1(G96), .A2(n669), .ZN(n841) );
  NAND2_X1 U750 ( .A1(n841), .A2(G2106), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G108), .A2(G120), .ZN(n670) );
  NOR2_X1 U752 ( .A1(G237), .A2(n670), .ZN(n671) );
  NAND2_X1 U753 ( .A1(G69), .A2(n671), .ZN(n840) );
  NAND2_X1 U754 ( .A1(G567), .A2(n840), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n842) );
  NAND2_X1 U756 ( .A1(G483), .A2(G661), .ZN(n674) );
  NOR2_X1 U757 ( .A1(n842), .A2(n674), .ZN(n839) );
  NAND2_X1 U758 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U759 ( .A1(n675), .A2(G138), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G102), .A2(n893), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U762 ( .A(n678), .B(KEYINPUT92), .Z(n683) );
  NAND2_X1 U763 ( .A1(G126), .A2(n679), .ZN(n680) );
  XNOR2_X1 U764 ( .A(KEYINPUT91), .B(n680), .ZN(n681) );
  NOR2_X1 U765 ( .A1(n517), .A2(n681), .ZN(n682) );
  AND2_X1 U766 ( .A1(n683), .A2(n682), .ZN(G164) );
  XNOR2_X1 U767 ( .A(G1996), .B(KEYINPUT100), .ZN(n1009) );
  NOR2_X2 U768 ( .A1(G164), .A2(G1384), .ZN(n785) );
  INV_X1 U769 ( .A(n785), .ZN(n687) );
  AND2_X1 U770 ( .A1(G40), .A2(n684), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n686), .A2(n685), .ZN(n784) );
  NOR2_X1 U772 ( .A1(n687), .A2(n784), .ZN(n696) );
  INV_X1 U773 ( .A(n696), .ZN(n726) );
  INV_X1 U774 ( .A(n726), .ZN(n689) );
  NAND2_X1 U775 ( .A1(n1009), .A2(n689), .ZN(n688) );
  XNOR2_X1 U776 ( .A(n688), .B(KEYINPUT26), .ZN(n691) );
  INV_X1 U777 ( .A(n689), .ZN(n736) );
  NAND2_X1 U778 ( .A1(n736), .A2(G1341), .ZN(n690) );
  NAND2_X1 U779 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U781 ( .A1(n927), .A2(n694), .ZN(n703) );
  NAND2_X1 U782 ( .A1(n694), .A2(n927), .ZN(n701) );
  INV_X1 U783 ( .A(KEYINPUT97), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n695), .A2(n696), .ZN(n706) );
  INV_X1 U785 ( .A(n696), .ZN(n697) );
  NAND2_X1 U786 ( .A1(KEYINPUT97), .A2(n697), .ZN(n708) );
  NAND2_X1 U787 ( .A1(n706), .A2(n708), .ZN(n704) );
  NAND2_X1 U788 ( .A1(n721), .A2(G2067), .ZN(n699) );
  NAND2_X1 U789 ( .A1(G1348), .A2(n736), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n713) );
  NAND2_X1 U793 ( .A1(n704), .A2(G2072), .ZN(n705) );
  XNOR2_X1 U794 ( .A(n705), .B(KEYINPUT27), .ZN(n711) );
  AND2_X1 U795 ( .A1(G1956), .A2(n706), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U797 ( .A(n709), .B(KEYINPUT99), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U799 ( .A1(n939), .A2(n714), .ZN(n712) );
  NAND2_X1 U800 ( .A1(n713), .A2(n712), .ZN(n716) );
  NAND2_X1 U801 ( .A1(n716), .A2(n518), .ZN(n718) );
  XNOR2_X1 U802 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n717) );
  XNOR2_X1 U803 ( .A(n718), .B(n717), .ZN(n725) );
  XNOR2_X1 U804 ( .A(G1961), .B(KEYINPUT95), .ZN(n964) );
  NAND2_X1 U805 ( .A1(n726), .A2(n964), .ZN(n719) );
  XNOR2_X1 U806 ( .A(n719), .B(KEYINPUT96), .ZN(n723) );
  XNOR2_X1 U807 ( .A(G2078), .B(KEYINPUT98), .ZN(n720) );
  XNOR2_X1 U808 ( .A(n720), .B(KEYINPUT25), .ZN(n1010) );
  NAND2_X1 U809 ( .A1(n1010), .A2(n721), .ZN(n722) );
  NAND2_X1 U810 ( .A1(n723), .A2(n722), .ZN(n733) );
  NAND2_X1 U811 ( .A1(n733), .A2(G171), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n748) );
  NAND2_X1 U813 ( .A1(G8), .A2(n726), .ZN(n777) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n777), .ZN(n750) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n726), .ZN(n749) );
  NOR2_X1 U816 ( .A1(n750), .A2(n749), .ZN(n727) );
  NAND2_X1 U817 ( .A1(G8), .A2(n727), .ZN(n729) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n728) );
  XNOR2_X1 U819 ( .A(n729), .B(n728), .ZN(n730) );
  INV_X1 U820 ( .A(n730), .ZN(n732) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n734) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n777), .ZN(n738) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n736), .ZN(n737) );
  NOR2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U825 ( .A1(n739), .A2(G303), .ZN(n741) );
  NAND2_X1 U826 ( .A1(n748), .A2(n740), .ZN(n745) );
  INV_X1 U827 ( .A(n741), .ZN(n742) );
  OR2_X1 U828 ( .A1(n742), .A2(G286), .ZN(n743) );
  AND2_X1 U829 ( .A1(G8), .A2(n743), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U831 ( .A(n746), .B(KEYINPUT32), .ZN(n769) );
  NAND2_X1 U832 ( .A1(n748), .A2(n747), .ZN(n753) );
  AND2_X1 U833 ( .A1(G8), .A2(n749), .ZN(n751) );
  NOR2_X1 U834 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U835 ( .A1(n753), .A2(n752), .ZN(n770) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n937) );
  AND2_X1 U837 ( .A1(n770), .A2(n937), .ZN(n754) );
  NAND2_X1 U838 ( .A1(n769), .A2(n754), .ZN(n758) );
  INV_X1 U839 ( .A(n937), .ZN(n756) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n763) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U842 ( .A1(n763), .A2(n755), .ZN(n938) );
  OR2_X1 U843 ( .A1(n756), .A2(n938), .ZN(n757) );
  AND2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U845 ( .A1(n759), .A2(n777), .ZN(n760) );
  XNOR2_X1 U846 ( .A(n760), .B(KEYINPUT64), .ZN(n761) );
  NOR2_X1 U847 ( .A1(KEYINPUT33), .A2(n761), .ZN(n762) );
  XNOR2_X1 U848 ( .A(KEYINPUT103), .B(n762), .ZN(n766) );
  NAND2_X1 U849 ( .A1(n763), .A2(KEYINPUT33), .ZN(n764) );
  OR2_X1 U850 ( .A1(n777), .A2(n764), .ZN(n765) );
  XNOR2_X1 U851 ( .A(n767), .B(KEYINPUT104), .ZN(n768) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n948) );
  NAND2_X1 U853 ( .A1(n768), .A2(n948), .ZN(n781) );
  NAND2_X1 U854 ( .A1(n770), .A2(n769), .ZN(n773) );
  NOR2_X1 U855 ( .A1(G2090), .A2(G303), .ZN(n771) );
  NAND2_X1 U856 ( .A1(G8), .A2(n771), .ZN(n772) );
  NAND2_X1 U857 ( .A1(n773), .A2(n772), .ZN(n774) );
  NAND2_X1 U858 ( .A1(n774), .A2(n777), .ZN(n779) );
  NOR2_X1 U859 ( .A1(G1981), .A2(G305), .ZN(n775) );
  XOR2_X1 U860 ( .A(n775), .B(KEYINPUT24), .Z(n776) );
  OR2_X1 U861 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U862 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U863 ( .A1(n781), .A2(n780), .ZN(n783) );
  XNOR2_X1 U864 ( .A(n783), .B(n782), .ZN(n816) );
  XNOR2_X1 U865 ( .A(G1986), .B(G290), .ZN(n929) );
  NOR2_X1 U866 ( .A1(n785), .A2(n784), .ZN(n827) );
  NAND2_X1 U867 ( .A1(n929), .A2(n827), .ZN(n814) );
  NAND2_X1 U868 ( .A1(G140), .A2(n606), .ZN(n787) );
  NAND2_X1 U869 ( .A1(G104), .A2(n893), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U871 ( .A(KEYINPUT34), .B(n788), .ZN(n794) );
  NAND2_X1 U872 ( .A1(G128), .A2(n679), .ZN(n790) );
  NAND2_X1 U873 ( .A1(G116), .A2(n896), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U875 ( .A(KEYINPUT93), .B(n791), .ZN(n792) );
  XNOR2_X1 U876 ( .A(KEYINPUT35), .B(n792), .ZN(n793) );
  NOR2_X1 U877 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U878 ( .A(KEYINPUT36), .B(n795), .ZN(n873) );
  XNOR2_X1 U879 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NOR2_X1 U880 ( .A1(n873), .A2(n825), .ZN(n796) );
  XNOR2_X1 U881 ( .A(n796), .B(KEYINPUT94), .ZN(n1002) );
  NAND2_X1 U882 ( .A1(n827), .A2(n1002), .ZN(n823) );
  NAND2_X1 U883 ( .A1(G131), .A2(n606), .ZN(n798) );
  NAND2_X1 U884 ( .A1(G119), .A2(n679), .ZN(n797) );
  NAND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G95), .A2(n893), .ZN(n800) );
  NAND2_X1 U887 ( .A1(G107), .A2(n896), .ZN(n799) );
  NAND2_X1 U888 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n802), .A2(n801), .ZN(n902) );
  INV_X1 U890 ( .A(G1991), .ZN(n843) );
  NOR2_X1 U891 ( .A1(n902), .A2(n843), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G141), .A2(n606), .ZN(n804) );
  NAND2_X1 U893 ( .A1(G129), .A2(n679), .ZN(n803) );
  NAND2_X1 U894 ( .A1(n804), .A2(n803), .ZN(n807) );
  NAND2_X1 U895 ( .A1(n893), .A2(G105), .ZN(n805) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n805), .Z(n806) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n809) );
  NAND2_X1 U898 ( .A1(n896), .A2(G117), .ZN(n808) );
  NAND2_X1 U899 ( .A1(n809), .A2(n808), .ZN(n886) );
  AND2_X1 U900 ( .A1(G1996), .A2(n886), .ZN(n810) );
  NOR2_X1 U901 ( .A1(n811), .A2(n810), .ZN(n996) );
  INV_X1 U902 ( .A(n996), .ZN(n812) );
  NAND2_X1 U903 ( .A1(n812), .A2(n827), .ZN(n817) );
  AND2_X1 U904 ( .A1(n823), .A2(n817), .ZN(n813) );
  AND2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U906 ( .A1(n816), .A2(n815), .ZN(n830) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n886), .ZN(n993) );
  INV_X1 U908 ( .A(n817), .ZN(n820) );
  AND2_X1 U909 ( .A1(n843), .A2(n902), .ZN(n989) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U911 ( .A1(n989), .A2(n818), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U913 ( .A1(n993), .A2(n821), .ZN(n822) );
  XNOR2_X1 U914 ( .A(KEYINPUT39), .B(n822), .ZN(n824) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U916 ( .A1(n825), .A2(n873), .ZN(n1003) );
  NAND2_X1 U917 ( .A1(n826), .A2(n1003), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U919 ( .A1(n830), .A2(n829), .ZN(n832) );
  XNOR2_X1 U920 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n831) );
  XNOR2_X1 U921 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U922 ( .A1(n833), .A2(G2106), .ZN(n834) );
  XNOR2_X1 U923 ( .A(n834), .B(KEYINPUT108), .ZN(G217) );
  NAND2_X1 U924 ( .A1(G15), .A2(G2), .ZN(n836) );
  INV_X1 U925 ( .A(G661), .ZN(n835) );
  NOR2_X1 U926 ( .A1(n836), .A2(n835), .ZN(n837) );
  XNOR2_X1 U927 ( .A(n837), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U929 ( .A1(n839), .A2(n838), .ZN(G188) );
  XOR2_X1 U930 ( .A(G96), .B(KEYINPUT110), .Z(G221) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G82), .ZN(G220) );
  INV_X1 U936 ( .A(G69), .ZN(G235) );
  NOR2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U938 ( .A(G325), .ZN(G261) );
  INV_X1 U939 ( .A(n842), .ZN(G319) );
  XOR2_X1 U940 ( .A(G1981), .B(G1966), .Z(n845) );
  XOR2_X1 U941 ( .A(G1996), .B(n843), .Z(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n855) );
  XOR2_X1 U943 ( .A(KEYINPUT41), .B(G2474), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1956), .B(KEYINPUT113), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1961), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U950 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(G229) );
  XOR2_X1 U953 ( .A(KEYINPUT43), .B(KEYINPUT42), .Z(n857) );
  XNOR2_X1 U954 ( .A(G2678), .B(KEYINPUT112), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(KEYINPUT111), .B(G2090), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2100), .B(G2096), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U962 ( .A(G2078), .B(G2084), .Z(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U964 ( .A1(G124), .A2(n679), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U966 ( .A1(n893), .A2(G100), .ZN(n867) );
  NAND2_X1 U967 ( .A1(n868), .A2(n867), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G136), .A2(n606), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G112), .A2(n896), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U971 ( .A1(n872), .A2(n871), .ZN(G162) );
  XNOR2_X1 U972 ( .A(n873), .B(n988), .ZN(n875) );
  XNOR2_X1 U973 ( .A(G164), .B(G160), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n885) );
  NAND2_X1 U975 ( .A1(G130), .A2(n679), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G118), .A2(n896), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n883) );
  NAND2_X1 U978 ( .A1(G142), .A2(n606), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G106), .A2(n893), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U981 ( .A(KEYINPUT116), .B(n880), .Z(n881) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n881), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n885), .B(n884), .Z(n888) );
  XOR2_X1 U985 ( .A(n886), .B(G162), .Z(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n892) );
  XOR2_X1 U987 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n890) );
  XNOR2_X1 U988 ( .A(KEYINPUT118), .B(KEYINPUT48), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U990 ( .A(n892), .B(n891), .Z(n904) );
  NAND2_X1 U991 ( .A1(G139), .A2(n606), .ZN(n895) );
  NAND2_X1 U992 ( .A1(G103), .A2(n893), .ZN(n894) );
  NAND2_X1 U993 ( .A1(n895), .A2(n894), .ZN(n901) );
  NAND2_X1 U994 ( .A1(G127), .A2(n679), .ZN(n898) );
  NAND2_X1 U995 ( .A1(G115), .A2(n896), .ZN(n897) );
  NAND2_X1 U996 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n899), .Z(n900) );
  NOR2_X1 U998 ( .A1(n901), .A2(n900), .ZN(n984) );
  XNOR2_X1 U999 ( .A(n902), .B(n984), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(n906), .B(KEYINPUT119), .ZN(n908) );
  XOR2_X1 U1003 ( .A(n927), .B(G286), .Z(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n909) );
  XOR2_X1 U1005 ( .A(G171), .B(n909), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G397) );
  XOR2_X1 U1007 ( .A(G2454), .B(G2435), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G2438), .B(G2427), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n919) );
  XOR2_X1 U1010 ( .A(KEYINPUT107), .B(G2446), .Z(n914) );
  XNOR2_X1 U1011 ( .A(G2443), .B(G2430), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1013 ( .A(n915), .B(G2451), .Z(n917) );
  XNOR2_X1 U1014 ( .A(G1341), .B(G1348), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(n917), .B(n916), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(n919), .B(n918), .ZN(n920) );
  NAND2_X1 U1017 ( .A1(n920), .A2(G14), .ZN(n926) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n926), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G229), .A2(G227), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(KEYINPUT49), .B(n921), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n925) );
  NOR2_X1 U1022 ( .A1(G395), .A2(G397), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G303), .ZN(G166) );
  INV_X1 U1026 ( .A(n926), .ZN(G401) );
  INV_X1 U1027 ( .A(G16), .ZN(n952) );
  XOR2_X1 U1028 ( .A(G1348), .B(n927), .Z(n928) );
  NOR2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G1961), .B(KEYINPUT122), .ZN(n930) );
  XOR2_X1 U1031 ( .A(n930), .B(G301), .Z(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n936) );
  XOR2_X1 U1033 ( .A(G1341), .B(n933), .Z(n934) );
  XNOR2_X1 U1034 ( .A(KEYINPUT124), .B(n934), .ZN(n935) );
  NOR2_X1 U1035 ( .A1(n936), .A2(n935), .ZN(n946) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(n939), .B(G1956), .ZN(n941) );
  NAND2_X1 U1038 ( .A1(G1971), .A2(G303), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1041 ( .A(KEYINPUT123), .B(n944), .Z(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n951) );
  XNOR2_X1 U1043 ( .A(G1966), .B(G168), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1045 ( .A(KEYINPUT57), .B(n949), .Z(n950) );
  NOR2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n978) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n978), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(KEYINPUT56), .A2(n953), .ZN(n954) );
  NAND2_X1 U1049 ( .A1(G11), .A2(n954), .ZN(n983) );
  XOR2_X1 U1050 ( .A(G1341), .B(G19), .Z(n958) );
  XNOR2_X1 U1051 ( .A(G1956), .B(G20), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G1981), .B(G6), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT126), .B(n959), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT59), .B(G1348), .Z(n960) );
  XNOR2_X1 U1057 ( .A(G4), .B(n960), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT60), .B(n963), .ZN(n974) );
  XNOR2_X1 U1060 ( .A(KEYINPUT125), .B(G5), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(n965), .B(n964), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(G23), .B(G1976), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n969) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1067 ( .A(KEYINPUT58), .B(n970), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(G21), .B(G1966), .ZN(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n977), .B(KEYINPUT61), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(KEYINPUT56), .A2(n978), .ZN(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1075 ( .A1(G16), .A2(n981), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n1008) );
  XOR2_X1 U1077 ( .A(G2072), .B(n984), .Z(n986) );
  XOR2_X1 U1078 ( .A(G164), .B(G2078), .Z(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT50), .B(n987), .ZN(n1000) );
  XNOR2_X1 U1081 ( .A(G160), .B(G2084), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n998) );
  XOR2_X1 U1084 ( .A(G2090), .B(G162), .Z(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1086 ( .A(KEYINPUT51), .B(n994), .Z(n995) );
  NAND2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1004) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(KEYINPUT52), .B(n1005), .ZN(n1006) );
  NAND2_X1 U1093 ( .A1(n1006), .A2(G29), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1031) );
  XOR2_X1 U1095 ( .A(n1009), .B(G32), .Z(n1012) );
  XNOR2_X1 U1096 ( .A(G27), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1097 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(KEYINPUT120), .B(n1013), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(G25), .B(G1991), .Z(n1014) );
  NAND2_X1 U1100 ( .A1(n1014), .A2(G28), .ZN(n1015) );
  NOR2_X1 U1101 ( .A1(n1016), .A2(n1015), .ZN(n1020) );
  XNOR2_X1 U1102 ( .A(G2067), .B(G26), .ZN(n1018) );
  XNOR2_X1 U1103 ( .A(G33), .B(G2072), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(n1021), .B(KEYINPUT53), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(G2084), .B(G34), .Z(n1022) );
  XNOR2_X1 U1108 ( .A(KEYINPUT54), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  XNOR2_X1 U1110 ( .A(G35), .B(G2090), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(KEYINPUT121), .B(n1027), .Z(n1028) );
  NOR2_X1 U1113 ( .A1(G29), .A2(n1028), .ZN(n1029) );
  XOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT55), .Z(n1030) );
  NOR2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1032), .Z(n1033) );
  XOR2_X1 U1117 ( .A(KEYINPUT127), .B(n1033), .Z(G150) );
  INV_X1 U1118 ( .A(G150), .ZN(G311) );
endmodule

