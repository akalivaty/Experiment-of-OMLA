//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n187));
  OAI21_X1  g001(.A(G214), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT66), .B1(new_n190), .B2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT66), .ZN(new_n192));
  INV_X1    g006(.A(G119), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n192), .A2(new_n193), .A3(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(G119), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G113), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT2), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G113), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n196), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n200), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n203), .A2(new_n195), .A3(new_n194), .A4(new_n191), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT67), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT74), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n211), .A2(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n213));
  OAI22_X1  g027(.A1(new_n211), .A2(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT74), .A4(G104), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT4), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G101), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n213), .A2(new_n214), .A3(new_n222), .A4(new_n217), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT75), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n224), .A2(new_n219), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(KEYINPUT75), .A3(G101), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT4), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n225), .A2(KEYINPUT76), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT76), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n226), .A2(KEYINPUT4), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n219), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n210), .B(new_n221), .C1(new_n228), .C2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT5), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n193), .A3(G116), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n196), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n204), .B1(new_n236), .B2(new_n197), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n212), .A2(KEYINPUT77), .A3(G107), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n216), .A2(G104), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT77), .B1(new_n212), .B2(G107), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n223), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(G110), .B(G122), .Z(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n233), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(G143), .B(G146), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(G128), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n249), .A3(new_n250), .ZN(new_n257));
  INV_X1    g071(.A(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G143), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n255), .ZN(new_n260));
  INV_X1    g074(.A(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n253), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G125), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n260), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n252), .A2(KEYINPUT0), .A3(G128), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n266), .B1(new_n265), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT80), .B1(new_n271), .B2(new_n265), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT7), .ZN(new_n274));
  INV_X1    g088(.A(G224), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G953), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n273), .B1(new_n274), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n272), .B(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(new_n246), .B(KEYINPUT8), .Z(new_n279));
  AND2_X1   g093(.A1(new_n237), .A2(new_n243), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(new_n244), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n248), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G902), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT81), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT76), .B1(new_n225), .B2(new_n227), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n230), .A2(new_n229), .A3(new_n231), .ZN(new_n288));
  AOI211_X1 g102(.A(new_n209), .B(new_n220), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n246), .B1(new_n289), .B2(new_n244), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT6), .A3(new_n248), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n272), .B(new_n276), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n293), .B(new_n246), .C1(new_n289), .C2(new_n244), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(KEYINPUT81), .A3(new_n283), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n286), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(G210), .B1(G237), .B2(G902), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n286), .A2(new_n295), .A3(new_n298), .A4(new_n296), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n189), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G952), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n304), .B1(G234), .B2(G237), .ZN(new_n305));
  INV_X1    g119(.A(G234), .ZN(new_n306));
  INV_X1    g120(.A(G237), .ZN(new_n307));
  OAI211_X1 g121(.A(G902), .B(G953), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT92), .Z(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT21), .B(G898), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n302), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT20), .ZN(new_n314));
  NOR2_X1   g128(.A1(G475), .A2(G902), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT86), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G113), .B(G122), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n318), .A2(KEYINPUT84), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(KEYINPUT84), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n319), .A2(G104), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(G104), .B1(new_n319), .B2(new_n320), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n324));
  AND2_X1   g138(.A1(G125), .A2(G140), .ZN(new_n325));
  NOR2_X1   g139(.A1(G125), .A2(G140), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n265), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(G125), .A2(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(KEYINPUT82), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT19), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n325), .A2(new_n326), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(KEYINPUT19), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n258), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT83), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT16), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n328), .A3(G125), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n341), .B1(new_n334), .B2(new_n340), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n342), .A2(new_n258), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n307), .A2(new_n303), .A3(G214), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n254), .ZN(new_n345));
  NOR2_X1   g159(.A1(G237), .A2(G953), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(G143), .A3(G214), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G131), .ZN(new_n349));
  INV_X1    g163(.A(G131), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n333), .A2(KEYINPUT83), .A3(new_n258), .A4(new_n336), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n339), .A2(new_n343), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(KEYINPUT18), .A2(G131), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n348), .B(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n329), .A2(new_n330), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n258), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT72), .ZN(new_n359));
  XNOR2_X1  g173(.A(new_n358), .B(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n258), .B1(new_n327), .B2(new_n331), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n356), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n323), .B1(new_n354), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT17), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n349), .A2(new_n364), .A3(new_n351), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n342), .A2(new_n258), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n348), .A2(KEYINPUT17), .A3(G131), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n365), .A2(new_n366), .A3(new_n343), .A4(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT85), .B1(new_n321), .B2(new_n322), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n319), .A2(new_n320), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n212), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n319), .A2(G104), .A3(new_n320), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n362), .A2(new_n368), .A3(new_n369), .A4(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n314), .B(new_n317), .C1(new_n363), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT87), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n363), .A2(new_n376), .ZN(new_n380));
  OAI21_X1  g194(.A(KEYINPUT20), .B1(new_n380), .B2(new_n316), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT19), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n327), .B2(new_n331), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n383), .A2(G146), .A3(new_n335), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n343), .B(new_n352), .C1(new_n384), .C2(KEYINPUT83), .ZN(new_n385));
  INV_X1    g199(.A(new_n353), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n362), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n323), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n375), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(KEYINPUT87), .A3(new_n314), .A4(new_n317), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n379), .A2(new_n381), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n323), .B1(new_n362), .B2(new_n368), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n283), .B1(new_n376), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G475), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n392), .B2(new_n396), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(KEYINPUT9), .B(G234), .Z(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(G217), .A3(new_n303), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT89), .ZN(new_n403));
  INV_X1    g217(.A(G122), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(G116), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n190), .A2(KEYINPUT89), .A3(G122), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n407), .B1(new_n190), .B2(G122), .ZN(new_n408));
  OR2_X1    g222(.A1(new_n408), .A2(G107), .ZN(new_n409));
  INV_X1    g223(.A(G134), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT64), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT64), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G134), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n254), .A2(G128), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n261), .A2(G143), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n414), .B1(new_n416), .B2(new_n417), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n407), .A2(KEYINPUT14), .ZN(new_n422));
  AOI211_X1 g236(.A(new_n421), .B(new_n422), .C1(G116), .C2(new_n404), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n409), .B1(new_n419), .B2(new_n420), .C1(new_n423), .C2(new_n216), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n408), .A2(G107), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n409), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT90), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n409), .A2(KEYINPUT90), .A3(new_n425), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n417), .A2(KEYINPUT91), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n254), .A2(KEYINPUT13), .A3(G128), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT13), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n416), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT91), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n432), .B(new_n434), .C1(new_n435), .C2(new_n431), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n419), .B1(new_n436), .B2(G134), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n428), .A2(new_n429), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n402), .B1(new_n424), .B2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n424), .A2(new_n438), .A3(new_n402), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G478), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n443), .A2(KEYINPUT15), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n283), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n444), .B1(new_n442), .B2(new_n283), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G140), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n303), .A2(G227), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n271), .B(new_n221), .C1(new_n228), .C2(new_n232), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n253), .A2(KEYINPUT78), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n256), .A2(KEYINPUT1), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT78), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n251), .A2(new_n252), .A3(new_n456), .A4(G128), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n454), .A2(new_n262), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n243), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(KEYINPUT10), .A3(new_n263), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n453), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G137), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n465), .A2(KEYINPUT11), .A3(G134), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(KEYINPUT11), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n414), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n465), .A2(KEYINPUT11), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n350), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n411), .A2(new_n413), .B1(KEYINPUT11), .B2(new_n465), .ZN(new_n472));
  NOR4_X1   g286(.A1(new_n472), .A2(G131), .A3(new_n466), .A4(new_n469), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n464), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n453), .A2(new_n474), .A3(new_n462), .A4(new_n463), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n452), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n452), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT79), .B1(new_n459), .B2(new_n263), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT79), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n264), .A2(new_n481), .A3(new_n243), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n460), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n475), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT12), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n479), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n449), .B(new_n283), .C1(new_n478), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(G469), .A2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n452), .ZN(new_n489));
  INV_X1    g303(.A(new_n477), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n489), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n477), .A3(new_n452), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(G469), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G221), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n495), .B1(new_n400), .B2(new_n283), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n399), .A2(new_n448), .A3(new_n494), .A4(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n187), .B1(new_n313), .B2(new_n498), .ZN(new_n499));
  AND4_X1   g313(.A1(new_n399), .A2(new_n448), .A3(new_n497), .A4(new_n494), .ZN(new_n500));
  AOI211_X1 g314(.A(new_n311), .B(new_n189), .C1(new_n300), .C2(new_n301), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT93), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n261), .A2(G119), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT23), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n504), .B(new_n505), .C1(G119), .C2(new_n261), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n507), .ZN(new_n509));
  XNOR2_X1  g323(.A(G119), .B(G128), .ZN(new_n510));
  XOR2_X1   g324(.A(KEYINPUT24), .B(G110), .Z(new_n511));
  OAI211_X1 g325(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n360), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n343), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n504), .B1(G119), .B2(new_n261), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n515), .A2(G110), .B1(new_n510), .B2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n343), .A2(new_n366), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n303), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT22), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(G137), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n514), .A2(new_n522), .A3(new_n518), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n283), .A3(new_n525), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n527));
  OAI21_X1  g341(.A(G217), .B1(new_n306), .B2(G902), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT70), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(KEYINPUT25), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n524), .A2(new_n525), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n283), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT73), .Z(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n271), .B1(new_n471), .B2(new_n473), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n468), .A2(new_n350), .A3(new_n470), .ZN(new_n539));
  NAND2_X1  g353(.A1(G134), .A2(G137), .ZN(new_n540));
  OAI211_X1 g354(.A(G131), .B(new_n540), .C1(new_n415), .C2(G137), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n263), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n543), .A2(KEYINPUT30), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(KEYINPUT30), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n210), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n209), .A2(new_n538), .A3(new_n542), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT68), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT68), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n209), .A2(new_n538), .A3(new_n549), .A4(new_n542), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT31), .ZN(new_n552));
  XNOR2_X1  g366(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n553), .B(G101), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n346), .A2(G210), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n546), .A2(new_n551), .A3(new_n552), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT28), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n547), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n209), .B1(new_n538), .B2(new_n542), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n560), .B1(new_n548), .B2(new_n550), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n559), .B1(new_n561), .B2(new_n558), .ZN(new_n562));
  INV_X1    g376(.A(new_n556), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT31), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n546), .A2(new_n551), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n565), .A2(new_n563), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n557), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT69), .ZN(new_n568));
  NOR2_X1   g382(.A1(G472), .A2(G902), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT69), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n570), .B(new_n557), .C1(new_n564), .C2(new_n566), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT32), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n568), .A2(KEYINPUT32), .A3(new_n569), .A4(new_n571), .ZN(new_n575));
  INV_X1    g389(.A(new_n565), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n562), .A2(new_n556), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT29), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n556), .A2(KEYINPUT29), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n283), .B1(new_n562), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(G472), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n499), .A2(new_n502), .A3(new_n537), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  NAND3_X1  g399(.A1(new_n568), .A2(new_n283), .A3(new_n571), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G472), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n587), .A2(new_n537), .A3(new_n572), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n494), .A2(new_n497), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n441), .ZN(new_n592));
  OAI21_X1  g406(.A(KEYINPUT33), .B1(new_n592), .B2(new_n439), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT33), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n440), .A2(new_n594), .A3(new_n441), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n595), .A3(G478), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n442), .A2(new_n443), .A3(new_n283), .ZN(new_n597));
  NAND2_X1  g411(.A1(G478), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n392), .A2(new_n396), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT88), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n392), .A2(new_n396), .A3(new_n393), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n302), .A2(new_n312), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n591), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT34), .B(G104), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  INV_X1    g421(.A(new_n448), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n381), .A2(new_n377), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n608), .A2(new_n396), .A3(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n591), .A2(new_n313), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT35), .B(G107), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G9));
  NAND2_X1  g427(.A1(new_n587), .A2(new_n572), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n519), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n535), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n532), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT94), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT94), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n587), .A2(new_n621), .A3(new_n572), .A4(new_n618), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n620), .A2(new_n499), .A3(new_n502), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT95), .B(KEYINPUT37), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G110), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G12));
  AND2_X1   g440(.A1(new_n302), .A2(new_n618), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT96), .B(G900), .Z(new_n628));
  AND2_X1   g442(.A1(new_n309), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n629), .A2(new_n305), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT97), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n610), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n583), .A2(new_n627), .A3(new_n590), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  XNOR2_X1  g448(.A(new_n631), .B(KEYINPUT39), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n590), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT40), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(new_n618), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n300), .A2(new_n301), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT38), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT98), .B1(new_n561), .B2(new_n556), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n642), .B1(new_n565), .B2(new_n563), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n561), .A2(KEYINPUT98), .A3(new_n556), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n283), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n574), .A2(new_n575), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n448), .B1(new_n601), .B2(new_n602), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n639), .A2(new_n188), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G143), .ZN(G45));
  INV_X1    g465(.A(new_n631), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n603), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n583), .A2(new_n627), .A3(new_n590), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G146), .ZN(G48));
  AND3_X1   g470(.A1(new_n302), .A2(new_n312), .A3(new_n603), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n283), .B1(new_n478), .B2(new_n486), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(G469), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n497), .A3(new_n487), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT99), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n659), .A2(KEYINPUT99), .A3(new_n497), .A4(new_n487), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n657), .A2(new_n583), .A3(new_n537), .A4(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT100), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT41), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G113), .ZN(G15));
  NAND4_X1  g483(.A1(new_n583), .A2(new_n664), .A3(new_n537), .A4(new_n501), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n670), .A2(new_n610), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  AND3_X1   g486(.A1(new_n659), .A2(new_n497), .A3(new_n487), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n302), .A2(new_n673), .A3(KEYINPUT101), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT101), .B1(new_n302), .B2(new_n673), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n312), .B(new_n618), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n583), .A2(new_n399), .A3(new_n448), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n193), .ZN(G21));
  OR3_X1    g493(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT102), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  OAI211_X1 g495(.A(new_n680), .B(new_n569), .C1(new_n681), .C2(new_n567), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n587), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n683), .A2(new_n537), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n501), .A3(new_n649), .A4(new_n664), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G122), .ZN(G24));
  AND3_X1   g500(.A1(new_n587), .A2(new_n618), .A3(new_n682), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n687), .B(new_n654), .C1(new_n674), .C2(new_n675), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G125), .ZN(G27));
  XNOR2_X1  g503(.A(new_n574), .B(KEYINPUT104), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n575), .A3(new_n582), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n691), .A2(new_n537), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n300), .A2(new_n188), .A3(new_n301), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n694));
  NOR4_X1   g508(.A1(new_n653), .A2(new_n693), .A3(new_n589), .A4(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n589), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n583), .A2(new_n537), .A3(new_n654), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT103), .ZN(new_n698));
  AOI22_X1  g512(.A1(new_n692), .A2(new_n695), .B1(new_n698), .B2(new_n694), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT105), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G131), .ZN(G33));
  AND2_X1   g515(.A1(new_n583), .A2(new_n537), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(KEYINPUT106), .A3(new_n632), .A4(new_n696), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n583), .A2(new_n537), .A3(new_n632), .A4(new_n696), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT106), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G134), .ZN(G36));
  INV_X1    g522(.A(new_n599), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n399), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT43), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT109), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n712), .A2(KEYINPUT109), .A3(new_n714), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n614), .A3(new_n618), .A4(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n491), .A2(new_n492), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n492), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(G469), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n488), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT107), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n727), .A2(new_n732), .A3(KEYINPUT46), .A4(new_n488), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n730), .A2(new_n731), .A3(new_n487), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n497), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n722), .B1(new_n735), .B2(new_n635), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n497), .A4(new_n636), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n721), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n693), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n719), .B2(new_n720), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g556(.A(KEYINPUT110), .B(new_n739), .C1(new_n719), .C2(new_n720), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n738), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n465), .ZN(G39));
  AND3_X1   g559(.A1(new_n734), .A2(KEYINPUT47), .A3(new_n497), .ZN(new_n746));
  AOI21_X1  g560(.A(KEYINPUT47), .B1(new_n734), .B2(new_n497), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n654), .B(new_n739), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n537), .A3(new_n583), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n328), .ZN(G42));
  NAND2_X1  g564(.A1(new_n659), .A2(new_n487), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(KEYINPUT111), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT49), .Z(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n537), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n754), .A2(new_n189), .A3(new_n641), .ZN(new_n755));
  INV_X1    g569(.A(new_n647), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n497), .A3(new_n756), .A4(new_n711), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT53), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n302), .A2(new_n649), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n618), .A2(new_n631), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n647), .A2(new_n759), .A3(new_n590), .A4(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n688), .A2(new_n633), .A3(new_n655), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n300), .A2(new_n188), .A3(new_n301), .A4(new_n396), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n631), .ZN(new_n767));
  AND3_X1   g581(.A1(new_n618), .A2(new_n448), .A3(new_n609), .ZN(new_n768));
  AND4_X1   g582(.A1(new_n583), .A2(new_n590), .A3(new_n767), .A4(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT114), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n583), .A2(new_n590), .A3(new_n767), .A4(new_n768), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n706), .A2(new_n703), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n687), .A2(new_n654), .A3(new_n696), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n765), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n770), .A2(new_n773), .ZN(new_n777));
  AND4_X1   g591(.A1(new_n765), .A2(new_n707), .A3(new_n777), .A4(new_n775), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n764), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n692), .A2(new_n695), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n698), .A2(new_n694), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n604), .A2(KEYINPUT112), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n501), .A2(new_n784), .A3(new_n603), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n588), .A3(new_n785), .A4(new_n590), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n584), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n787), .B1(new_n584), .B2(new_n786), .ZN(new_n790));
  INV_X1    g604(.A(new_n399), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n448), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n588), .A2(new_n501), .A3(new_n590), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n623), .A2(new_n793), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n789), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n665), .A2(new_n666), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n665), .A2(new_n666), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n685), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI22_X1  g612(.A1(new_n676), .A2(new_n677), .B1(new_n610), .B2(new_n670), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n782), .A2(new_n795), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n758), .B1(new_n779), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n762), .B(KEYINPUT52), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n707), .A2(new_n777), .A3(new_n775), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT115), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n774), .A2(new_n765), .A3(new_n775), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n799), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n667), .A3(new_n810), .A4(new_n685), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n795), .A2(new_n811), .A3(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n667), .A3(new_n685), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n699), .B1(KEYINPUT118), .B2(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n808), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n802), .A2(new_n803), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT53), .B1(new_n764), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n818), .B1(new_n779), .B2(new_n801), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n584), .A2(new_n786), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT113), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n623), .A2(new_n793), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n822), .A3(new_n788), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n699), .A2(new_n823), .A3(new_n813), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n758), .B1(new_n804), .B2(KEYINPUT116), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n808), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n816), .A2(KEYINPUT117), .B1(new_n827), .B2(KEYINPUT54), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n827), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n752), .B(KEYINPUT119), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n497), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n831), .A2(new_n747), .A3(new_n746), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n684), .A2(new_n305), .A3(new_n715), .ZN(new_n833));
  OR3_X1    g647(.A1(new_n832), .A2(new_n693), .A3(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n641), .A2(new_n188), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n673), .B1(KEYINPUT120), .B2(KEYINPUT50), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n838), .ZN(new_n840));
  NOR4_X1   g654(.A1(new_n833), .A2(new_n840), .A3(new_n835), .A4(new_n836), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n739), .A2(new_n305), .A3(new_n673), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n715), .A2(new_n687), .A3(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n839), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n791), .A2(new_n709), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n756), .A2(new_n842), .A3(new_n537), .A4(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n834), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n304), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n692), .A2(new_n715), .A3(new_n842), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT48), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n756), .A2(new_n842), .A3(new_n537), .A4(new_n603), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n834), .A2(new_n844), .A3(KEYINPUT51), .A4(new_n846), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n851), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n674), .A2(new_n675), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n833), .A2(new_n855), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n828), .A2(new_n829), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(G952), .A2(G953), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n757), .B1(new_n857), .B2(new_n858), .ZN(G75));
  NOR2_X1   g673(.A1(new_n303), .A2(G952), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n291), .A2(new_n294), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(new_n292), .ZN(new_n863));
  XOR2_X1   g677(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n283), .B1(new_n802), .B2(new_n815), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(G210), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n865), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n866), .B2(G210), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n861), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(G51));
  NAND2_X1  g686(.A1(new_n802), .A2(new_n815), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n816), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n488), .B(KEYINPUT57), .Z(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n478), .A2(new_n486), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT123), .Z(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n727), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n866), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n860), .B1(new_n880), .B2(new_n882), .ZN(G54));
  NAND3_X1  g697(.A1(new_n866), .A2(KEYINPUT58), .A3(G475), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(new_n380), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n380), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n885), .A2(new_n886), .A3(new_n860), .ZN(G60));
  NAND2_X1  g701(.A1(new_n593), .A2(new_n595), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n598), .B(KEYINPUT59), .Z(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n890), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n892), .B1(new_n828), .B2(new_n829), .ZN(new_n893));
  AOI221_X4 g707(.A(new_n860), .B1(new_n875), .B2(new_n891), .C1(new_n893), .C2(new_n889), .ZN(G63));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT60), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n895), .B1(new_n873), .B2(new_n898), .ZN(new_n899));
  AOI211_X1 g713(.A(KEYINPUT124), .B(new_n897), .C1(new_n802), .C2(new_n815), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n616), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n795), .A2(new_n811), .A3(KEYINPUT53), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n782), .B1(new_n800), .B2(new_n810), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n779), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT53), .B1(new_n808), .B2(new_n824), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT124), .ZN(new_n907));
  INV_X1    g721(.A(new_n533), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n873), .A2(new_n895), .A3(new_n898), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n901), .A2(new_n910), .A3(new_n861), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n901), .A2(new_n910), .A3(KEYINPUT61), .A4(new_n861), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(G66));
  OAI21_X1  g729(.A(G953), .B1(new_n310), .B2(new_n275), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n823), .A2(new_n813), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n862), .B1(G898), .B2(new_n303), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G69));
  OR2_X1    g734(.A1(new_n544), .A2(new_n545), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n383), .A2(new_n335), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(G900), .B1(new_n923), .B2(G227), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G953), .ZN(new_n925));
  AND4_X1   g739(.A1(new_n692), .A2(new_n736), .A3(new_n737), .A4(new_n759), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n744), .A2(new_n749), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n688), .A2(new_n633), .A3(new_n655), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n929));
  INV_X1    g743(.A(new_n707), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n699), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n782), .A2(KEYINPUT125), .A3(new_n707), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(G953), .B1(new_n927), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n923), .B1(G227), .B2(new_n303), .ZN(new_n935));
  INV_X1    g749(.A(new_n928), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n650), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT62), .Z(new_n938));
  NOR2_X1   g752(.A1(new_n744), .A2(new_n749), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n702), .A2(new_n696), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n636), .B1(new_n792), .B2(new_n603), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n303), .ZN(new_n943));
  OAI221_X1 g757(.A(new_n925), .B1(new_n934), .B2(new_n935), .C1(new_n943), .C2(new_n923), .ZN(G72));
  NAND2_X1  g758(.A1(G472), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT63), .Z(new_n946));
  INV_X1    g760(.A(new_n917), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n576), .A2(new_n563), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n927), .A2(new_n917), .A3(new_n933), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n577), .B1(new_n951), .B2(new_n946), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n952), .A2(new_n860), .ZN(new_n953));
  INV_X1    g767(.A(new_n949), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n827), .A2(new_n577), .A3(new_n946), .A4(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT126), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT126), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n950), .A2(new_n953), .A3(new_n958), .A4(new_n955), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(G57));
endmodule


