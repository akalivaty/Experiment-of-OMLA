//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  AOI21_X1  g002(.A(G1gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT89), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI211_X1 g005(.A(new_n202), .B(KEYINPUT89), .C1(new_n203), .C2(G1gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G8gat), .ZN(new_n209));
  XOR2_X1   g008(.A(new_n209), .B(KEYINPUT91), .Z(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(G8gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT90), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT96), .ZN(new_n214));
  INV_X1    g013(.A(G71gat), .ZN(new_n215));
  INV_X1    g014(.A(G78gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(G71gat), .B2(G78gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n217), .B(KEYINPUT95), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n221), .A2(new_n218), .B1(new_n215), .B2(new_n216), .ZN(new_n223));
  OAI22_X1  g022(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT21), .ZN(new_n225));
  OR2_X1    g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n213), .A2(new_n214), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n225), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n212), .ZN(new_n229));
  INV_X1    g028(.A(new_n226), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT96), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G183gat), .B(G211gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT97), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n235), .B(new_n236), .Z(new_n237));
  AOI21_X1  g036(.A(new_n228), .B1(new_n227), .B2(new_n231), .ZN(new_n238));
  OR3_X1    g037(.A1(new_n233), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G127gat), .B(G155gat), .Z(new_n240));
  NAND2_X1  g039(.A1(G231gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n237), .B1(new_n233), .B2(new_n238), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n239), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n239), .B2(new_n243), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G43gat), .B(G50gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT15), .ZN(new_n248));
  OAI21_X1  g047(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT86), .ZN(new_n250));
  NOR3_X1   g049(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(G29gat), .A2(G36gat), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n247), .A2(KEYINPUT15), .ZN(new_n255));
  AND4_X1   g054(.A1(new_n248), .A2(new_n253), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  OR2_X1    g055(.A1(new_n251), .A2(KEYINPUT87), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(KEYINPUT87), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n248), .B1(new_n259), .B2(new_n254), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT17), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n262), .B(KEYINPUT88), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(KEYINPUT17), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT92), .ZN(new_n265));
  INV_X1    g064(.A(G99gat), .ZN(new_n266));
  INV_X1    g065(.A(G106gat), .ZN(new_n267));
  OAI21_X1  g066(.A(KEYINPUT8), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT98), .B(G85gat), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(new_n269), .B2(G92gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(G85gat), .A2(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT7), .Z(new_n272));
  XNOR2_X1  g071(.A(G99gat), .B(G106gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(KEYINPUT99), .ZN(new_n274));
  NOR3_X1   g073(.A1(new_n270), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(KEYINPUT99), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n276), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n265), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n261), .ZN(new_n282));
  AND2_X1   g081(.A1(G232gat), .A2(G233gat), .ZN(new_n283));
  AOI22_X1  g082(.A1(new_n282), .A2(new_n279), .B1(KEYINPUT41), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(G190gat), .B(G218gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AND3_X1   g085(.A1(new_n281), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n286), .B1(new_n281), .B2(new_n284), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n283), .A2(KEYINPUT41), .ZN(new_n289));
  XNOR2_X1  g088(.A(G134gat), .B(G162gat), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n289), .B(new_n290), .Z(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OR3_X1    g091(.A1(new_n287), .A2(new_n288), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n287), .B2(new_n288), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n246), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G230gat), .ZN(new_n298));
  INV_X1    g097(.A(G233gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n279), .B(new_n224), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OR3_X1    g102(.A1(new_n280), .A2(new_n302), .A3(new_n224), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n301), .A2(new_n298), .A3(new_n299), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G120gat), .B(G148gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(G176gat), .B(G204gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n305), .B2(new_n306), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n297), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(KEYINPUT93), .A2(KEYINPUT18), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n263), .A2(new_n213), .A3(new_n265), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n229), .A2(new_n282), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G229gat), .A2(G233gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n317), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n213), .A2(new_n261), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(KEYINPUT94), .A3(new_n319), .ZN(new_n325));
  OR3_X1    g124(.A1(new_n213), .A2(KEYINPUT94), .A3(new_n261), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n321), .B(KEYINPUT13), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n317), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n318), .A2(new_n321), .A3(new_n319), .A4(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(G113gat), .B(G141gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(G197gat), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT11), .B(G169gat), .Z(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n336), .B(KEYINPUT12), .Z(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n323), .A2(new_n329), .A3(new_n331), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n316), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT82), .ZN(new_n344));
  XOR2_X1   g143(.A(G211gat), .B(G218gat), .Z(new_n345));
  XOR2_X1   g144(.A(G197gat), .B(G204gat), .Z(new_n346));
  INV_X1    g145(.A(G218gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT72), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G218gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(G211gat), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT22), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT73), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n345), .B1(new_n357), .B2(KEYINPUT74), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT29), .ZN(new_n359));
  INV_X1    g158(.A(new_n346), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n351), .A2(KEYINPUT73), .A3(new_n352), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT73), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n364));
  INV_X1    g163(.A(new_n345), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n358), .A2(new_n359), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G148gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G141gat), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G148gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n375), .A2(KEYINPUT2), .ZN(new_n376));
  AND2_X1   g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT78), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380));
  NOR2_X1   g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n377), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G141gat), .B(G148gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n378), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n372), .A2(G148gat), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n370), .A2(G141gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n373), .A3(KEYINPUT77), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n380), .A3(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n377), .A2(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n385), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n369), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n393), .A2(new_n368), .A3(new_n384), .A4(new_n378), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n358), .A2(new_n366), .B1(new_n359), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n359), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n357), .A2(KEYINPUT74), .A3(new_n345), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n365), .B1(new_n363), .B2(new_n364), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n357), .B2(new_n345), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n363), .A2(new_n365), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT3), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n392), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n371), .A2(new_n373), .A3(KEYINPUT77), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT77), .B1(new_n371), .B2(new_n373), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n407), .B1(new_n410), .B2(new_n380), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n378), .A2(new_n384), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n403), .B1(new_n406), .B2(new_n413), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n398), .B(KEYINPUT81), .Z(new_n415));
  AOI22_X1  g214(.A1(new_n395), .A2(new_n399), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G78gat), .B(G106gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT31), .B(G50gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n344), .B1(new_n416), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n416), .B2(new_n420), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n413), .B1(new_n367), .B2(new_n368), .ZN(new_n424));
  INV_X1    g223(.A(new_n398), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n403), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n415), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n360), .B(new_n345), .C1(new_n361), .C2(new_n362), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n359), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n355), .A2(new_n356), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n345), .B1(new_n431), .B2(new_n360), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n368), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(new_n394), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n428), .B1(new_n434), .B2(new_n403), .ZN(new_n435));
  NOR4_X1   g234(.A1(new_n427), .A2(new_n435), .A3(G22gat), .A4(new_n419), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n421), .B1(new_n423), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n405), .A2(new_n359), .A3(new_n429), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n413), .B1(new_n438), .B2(new_n368), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n415), .B1(new_n439), .B2(new_n397), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n440), .B1(new_n424), .B2(new_n426), .ZN(new_n441));
  OAI21_X1  g240(.A(G22gat), .B1(new_n441), .B2(new_n419), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT82), .B1(new_n441), .B2(new_n419), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n416), .A2(new_n422), .A3(new_n420), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(G113gat), .ZN(new_n446));
  INV_X1    g245(.A(G120gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT1), .ZN(new_n449));
  NAND2_X1  g248(.A1(G113gat), .A2(G120gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G127gat), .B(G134gat), .ZN(new_n452));
  INV_X1    g251(.A(G127gat), .ZN(new_n453));
  OAI21_X1  g252(.A(KEYINPUT68), .B1(new_n453), .B2(G134gat), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n452), .B1(new_n451), .B2(new_n454), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT69), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n452), .ZN(new_n459));
  AND2_X1   g258(.A1(G113gat), .A2(G120gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(G113gat), .A2(G120gat), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT1), .ZN(new_n462));
  INV_X1    g261(.A(new_n454), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT69), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(G169gat), .ZN(new_n468));
  INV_X1    g267(.A(G176gat), .ZN(new_n469));
  AND2_X1   g268(.A1(new_n469), .A2(KEYINPUT64), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n469), .A2(KEYINPUT64), .ZN(new_n471));
  OAI211_X1 g270(.A(KEYINPUT23), .B(new_n468), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(G169gat), .A2(G176gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT23), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G169gat), .B2(G176gat), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n472), .A2(KEYINPUT65), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT65), .B1(new_n472), .B2(new_n475), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT25), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(G183gat), .A2(G190gat), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G183gat), .A2(G190gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n478), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n476), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(G169gat), .A2(G176gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT26), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT67), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT67), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n491), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n489), .A2(new_n490), .A3(new_n473), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(G183gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT27), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT27), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(G183gat), .ZN(new_n497));
  INV_X1    g296(.A(G190gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT28), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT27), .B1(new_n494), .B2(KEYINPUT66), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT66), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n496), .A3(G183gat), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT28), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(new_n498), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n493), .A2(new_n500), .A3(new_n482), .A4(new_n505), .ZN(new_n506));
  NOR3_X1   g305(.A1(new_n484), .A2(new_n480), .A3(new_n479), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n487), .A2(KEYINPUT23), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT23), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(G169gat), .B2(G176gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n508), .B1(new_n510), .B2(new_n487), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT25), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n467), .B1(new_n486), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n506), .A2(new_n512), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n457), .B1(new_n455), .B2(new_n456), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n464), .A2(KEYINPUT69), .A3(new_n465), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n472), .A2(new_n475), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT65), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n485), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n472), .A2(KEYINPUT65), .A3(new_n475), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n516), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n514), .A2(new_n515), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT34), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n514), .A2(KEYINPUT34), .A3(new_n515), .A4(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G15gat), .B(G43gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G71gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT70), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n532), .B(new_n215), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT70), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n534), .A2(new_n537), .A3(G99gat), .ZN(new_n538));
  AOI21_X1  g337(.A(G99gat), .B1(new_n534), .B2(new_n537), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n515), .B1(new_n514), .B2(new_n526), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(KEYINPUT33), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT32), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n514), .A2(new_n526), .ZN(new_n546));
  INV_X1    g345(.A(new_n515), .ZN(new_n547));
  AOI221_X4 g346(.A(new_n543), .B1(new_n540), .B2(KEYINPUT33), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n531), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n516), .A2(new_n519), .A3(new_n525), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n519), .B1(new_n516), .B2(new_n525), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT32), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT33), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n555), .A3(new_n540), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n542), .A2(new_n544), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n529), .A2(new_n530), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n437), .A2(new_n445), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT30), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n401), .A2(new_n402), .ZN(new_n564));
  NAND2_X1  g363(.A1(G226gat), .A2(G233gat), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n516), .A2(new_n525), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(new_n359), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n516), .B2(new_n525), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n566), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n358), .A2(new_n366), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT29), .B1(new_n516), .B2(new_n525), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n571), .B(new_n572), .C1(new_n566), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G8gat), .B(G36gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(G64gat), .B(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT76), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT76), .ZN(new_n581));
  AOI211_X1 g380(.A(new_n581), .B(new_n578), .C1(new_n570), .C2(new_n574), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n563), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n575), .A2(new_n579), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n568), .A2(new_n564), .A3(new_n569), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n359), .B1(new_n486), .B2(new_n513), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n565), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n572), .B1(new_n588), .B2(new_n571), .ZN(new_n589));
  OAI211_X1 g388(.A(KEYINPUT30), .B(new_n579), .C1(new_n586), .C2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT75), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n578), .B1(new_n570), .B2(new_n574), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n593), .A2(KEYINPUT75), .A3(KEYINPUT30), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n583), .A2(new_n585), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(KEYINPUT3), .B1(new_n411), .B2(new_n412), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT79), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n455), .B2(new_n456), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n464), .A2(KEYINPUT79), .A3(new_n465), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n596), .A2(new_n396), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n413), .A2(new_n519), .A3(KEYINPUT4), .ZN(new_n602));
  NAND2_X1  g401(.A1(G225gat), .A2(G233gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n464), .A2(new_n465), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n385), .A2(new_n393), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT4), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT80), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n394), .A2(new_n600), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n603), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n393), .A2(new_n385), .B1(new_n598), .B2(new_n599), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n608), .A2(new_n614), .A3(KEYINPUT5), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n606), .B1(new_n467), .B2(new_n394), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n604), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n611), .A2(KEYINPUT5), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n616), .A2(new_n601), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G1gat), .B(G29gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(G85gat), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT0), .B(G57gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT6), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n615), .A2(new_n619), .A3(new_n624), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(KEYINPUT6), .A3(new_n625), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n595), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n562), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT35), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT71), .ZN(new_n635));
  OAI22_X1  g434(.A1(new_n545), .A2(new_n548), .B1(new_n635), .B2(new_n531), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n556), .A2(new_n557), .A3(new_n558), .A4(KEYINPUT71), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AND4_X1   g437(.A1(KEYINPUT35), .A2(new_n437), .A3(new_n445), .A4(new_n638), .ZN(new_n639));
  AOI22_X1  g438(.A1(new_n633), .A2(new_n634), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n545), .A2(new_n548), .A3(new_n531), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n558), .B1(new_n556), .B2(new_n557), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n637), .A3(KEYINPUT36), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n630), .ZN(new_n647));
  AND2_X1   g446(.A1(new_n592), .A2(new_n594), .ZN(new_n648));
  NAND4_X1  g447(.A1(new_n647), .A2(new_n648), .A3(new_n585), .A4(new_n583), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n437), .A2(new_n445), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n646), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n616), .A2(new_n601), .A3(new_n617), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n611), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n610), .B1(new_n612), .B2(new_n613), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n603), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n653), .A2(KEYINPUT39), .A3(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n611), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n624), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT84), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n659), .A2(KEYINPUT84), .A3(new_n624), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT85), .B1(new_n664), .B2(KEYINPUT40), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n624), .B1(new_n615), .B2(new_n619), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n664), .B2(KEYINPUT40), .ZN(new_n667));
  INV_X1    g466(.A(new_n663), .ZN(new_n668));
  AOI21_X1  g467(.A(KEYINPUT84), .B1(new_n659), .B2(new_n624), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n656), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT85), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND4_X1   g472(.A1(new_n595), .A2(new_n665), .A3(new_n667), .A4(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT37), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n570), .A2(new_n675), .A3(new_n574), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n570), .B2(new_n574), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n578), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT38), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n575), .A2(new_n579), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n581), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT38), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n684), .B(new_n578), .C1(new_n676), .C2(new_n677), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n679), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(new_n445), .B(new_n437), .C1(new_n686), .C2(new_n647), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n651), .B1(new_n674), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n640), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n343), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n647), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT100), .B(G1gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1324gat));
  INV_X1    g492(.A(new_n690), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT16), .B(G8gat), .Z(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n595), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT42), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT30), .B1(new_n681), .B2(new_n682), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n592), .A2(new_n594), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n698), .A2(new_n699), .A3(new_n584), .ZN(new_n700));
  OAI21_X1  g499(.A(G8gat), .B1(new_n690), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n697), .A2(new_n701), .ZN(G1325gat));
  AOI21_X1  g501(.A(G15gat), .B1(new_n694), .B2(new_n560), .ZN(new_n703));
  INV_X1    g502(.A(new_n646), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n690), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(G15gat), .B2(new_n705), .ZN(G1326gat));
  AND2_X1   g505(.A1(new_n437), .A2(new_n445), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n690), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT43), .B(G22gat), .Z(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  NAND2_X1  g509(.A1(new_n639), .A2(new_n632), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n634), .B1(new_n649), .B2(new_n561), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n595), .A2(new_n665), .A3(new_n667), .A4(new_n673), .ZN(new_n714));
  OAI211_X1 g513(.A(new_n714), .B(new_n707), .C1(new_n647), .C2(new_n686), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n651), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n295), .ZN(new_n717));
  OR2_X1    g516(.A1(new_n244), .A2(new_n245), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(new_n342), .A3(new_n314), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(G29gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n722), .A3(new_n631), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n718), .B(KEYINPUT102), .ZN(new_n725));
  AND3_X1   g524(.A1(new_n338), .A2(KEYINPUT101), .A3(new_n340), .ZN(new_n726));
  AOI21_X1  g525(.A(KEYINPUT101), .B1(new_n338), .B2(new_n340), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n315), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT103), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n689), .B2(new_n296), .ZN(new_n732));
  AOI211_X1 g531(.A(KEYINPUT44), .B(new_n295), .C1(new_n640), .C2(new_n688), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n631), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n724), .B1(new_n737), .B2(new_n722), .ZN(G1328gat));
  NOR3_X1   g537(.A1(new_n720), .A2(G36gat), .A3(new_n700), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n735), .A2(new_n595), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(G36gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(G1329gat));
  INV_X1    g544(.A(new_n560), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n720), .A2(G43gat), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n735), .A2(new_n646), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g550(.A1(new_n730), .A2(new_n734), .ZN(new_n752));
  OAI21_X1  g551(.A(G50gat), .B1(new_n752), .B2(new_n707), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n721), .A2(KEYINPUT106), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n650), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n753), .B1(G50gat), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT48), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1331gat));
  INV_X1    g558(.A(new_n728), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n297), .A3(new_n314), .ZN(new_n761));
  XOR2_X1   g560(.A(new_n761), .B(KEYINPUT107), .Z(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(new_n689), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n631), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g565(.A(new_n700), .B(new_n763), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n764), .A2(new_n215), .A3(new_n560), .ZN(new_n770));
  OAI21_X1  g569(.A(G71gat), .B1(new_n763), .B2(new_n704), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g572(.A1(new_n763), .A2(new_n707), .ZN(new_n774));
  XNOR2_X1  g573(.A(KEYINPUT108), .B(G78gat), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n774), .B(new_n775), .ZN(G1335gat));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n689), .B2(new_n296), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT110), .B(new_n295), .C1(new_n640), .C2(new_n688), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n728), .A2(new_n718), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT51), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n716), .B2(new_n295), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n689), .A2(new_n777), .A3(new_n296), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n783), .A2(KEYINPUT51), .A3(new_n781), .A4(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n787), .A2(new_n647), .A3(new_n315), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n246), .B(new_n314), .C1(new_n726), .C2(new_n727), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n732), .B2(new_n733), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT109), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(new_n790), .C1(new_n732), .C2(new_n733), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n631), .ZN(new_n796));
  MUX2_X1   g595(.A(new_n788), .B(new_n796), .S(new_n269), .Z(G1336gat));
  INV_X1    g596(.A(new_n787), .ZN(new_n798));
  INV_X1    g597(.A(G92gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n314), .A2(new_n799), .A3(new_n595), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n734), .A2(new_n595), .A3(new_n790), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(new_n803), .B2(G92gat), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n799), .B1(new_n795), .B2(new_n595), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n806), .B1(new_n798), .B2(new_n801), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(G1337gat));
  NAND2_X1  g608(.A1(new_n795), .A2(new_n646), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n266), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n798), .A2(new_n560), .A3(new_n314), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n266), .ZN(G1338gat));
  NOR2_X1   g612(.A1(new_n707), .A2(G106gat), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n314), .B(new_n814), .C1(new_n782), .C2(new_n786), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n734), .A2(new_n650), .A3(new_n790), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n816), .B2(G106gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n267), .B1(new_n795), .B2(new_n650), .ZN(new_n820));
  INV_X1    g619(.A(new_n814), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n783), .A2(new_n781), .A3(new_n784), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI211_X1 g623(.A(new_n315), .B(new_n821), .C1(new_n824), .C2(new_n785), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n819), .B(KEYINPUT53), .C1(new_n820), .C2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n707), .B1(new_n792), .B2(new_n794), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n815), .B1(new_n267), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n819), .B1(new_n829), .B2(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n818), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT113), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n833), .B(new_n818), .C1(new_n827), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT101), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n341), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n338), .A2(KEYINPUT101), .A3(new_n340), .ZN(new_n838));
  INV_X1    g637(.A(new_n305), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n303), .A2(new_n304), .A3(new_n300), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(KEYINPUT54), .A3(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n311), .B1(new_n305), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n843), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n312), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n837), .A2(new_n838), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n325), .A2(new_n326), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n327), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT114), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n320), .A2(new_n322), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n855), .A3(new_n327), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n336), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT115), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n857), .A2(new_n860), .A3(new_n336), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n859), .A2(new_n340), .A3(new_n314), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n296), .B1(new_n850), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n295), .A2(new_n848), .ZN(new_n864));
  AND4_X1   g663(.A1(new_n340), .A2(new_n864), .A3(new_n859), .A4(new_n861), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n725), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n760), .A2(new_n297), .A3(new_n315), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n647), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n650), .B1(new_n637), .B2(new_n636), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n700), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n446), .A3(new_n728), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n868), .A2(new_n700), .A3(new_n562), .ZN(new_n874));
  OAI21_X1  g673(.A(G113gat), .B1(new_n874), .B2(new_n342), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1340gat));
  NAND3_X1  g675(.A1(new_n872), .A2(new_n447), .A3(new_n314), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n874), .A2(new_n315), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n878), .A2(KEYINPUT116), .A3(G120gat), .ZN(new_n879));
  AOI21_X1  g678(.A(KEYINPUT116), .B1(new_n878), .B2(G120gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(G1341gat));
  NAND3_X1  g680(.A1(new_n872), .A2(new_n453), .A3(new_n718), .ZN(new_n882));
  OAI21_X1  g681(.A(G127gat), .B1(new_n874), .B2(new_n725), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(KEYINPUT117), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT117), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n882), .A2(new_n886), .A3(new_n883), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n887), .ZN(G1342gat));
  OR2_X1    g687(.A1(new_n295), .A2(G134gat), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n871), .A2(KEYINPUT56), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(G134gat), .B1(new_n874), .B2(new_n295), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT56), .B1(new_n871), .B2(new_n889), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G1343gat));
  NOR3_X1   g692(.A1(new_n646), .A2(new_n647), .A3(new_n595), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n845), .A2(KEYINPUT118), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n841), .A2(new_n843), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n844), .A2(KEYINPUT118), .A3(new_n845), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n341), .A2(new_n312), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n296), .B1(new_n862), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n246), .B1(new_n900), .B2(new_n865), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n867), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n650), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n895), .B1(new_n903), .B2(KEYINPUT57), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT57), .B(new_n707), .C1(new_n866), .C2(new_n867), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n904), .A2(new_n906), .A3(new_n341), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(G141gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n707), .B1(new_n866), .B2(new_n867), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n894), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n910), .A2(G141gat), .A3(new_n342), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(KEYINPUT120), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT58), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n914), .B1(new_n904), .B2(new_n906), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n707), .B1(new_n901), .B2(new_n867), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n894), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n918), .A2(new_n905), .A3(KEYINPUT119), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n728), .B1(new_n915), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(KEYINPUT58), .A3(G141gat), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT58), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n911), .B1(KEYINPUT120), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n913), .B1(new_n921), .B2(new_n923), .ZN(G1344gat));
  OAI21_X1  g723(.A(new_n901), .B1(new_n341), .B2(new_n316), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n917), .A3(new_n650), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n909), .B2(new_n917), .ZN(new_n927));
  OR2_X1    g726(.A1(new_n927), .A2(new_n315), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT59), .B(G148gat), .C1(new_n928), .C2(new_n895), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT59), .ZN(new_n930));
  OAI211_X1 g729(.A(new_n930), .B(new_n314), .C1(new_n915), .C2(new_n919), .ZN(new_n931));
  INV_X1    g730(.A(new_n910), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n932), .B2(new_n314), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n929), .B(new_n931), .C1(G148gat), .C2(new_n933), .ZN(G1345gat));
  AOI21_X1  g733(.A(G155gat), .B1(new_n932), .B2(new_n718), .ZN(new_n935));
  INV_X1    g734(.A(new_n915), .ZN(new_n936));
  INV_X1    g735(.A(new_n919), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n725), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n935), .B1(new_n938), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g738(.A(G162gat), .B1(new_n932), .B2(new_n296), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n295), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(G162gat), .ZN(G1347gat));
  AOI21_X1  g741(.A(new_n631), .B1(new_n866), .B2(new_n867), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n943), .A2(new_n595), .A3(new_n869), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT121), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n945), .A2(new_n468), .A3(new_n728), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n943), .A2(new_n595), .A3(new_n562), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n595), .A4(new_n562), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n341), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n946), .B1(new_n468), .B2(new_n952), .ZN(G1348gat));
  AOI21_X1  g752(.A(G176gat), .B1(new_n945), .B2(new_n314), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n470), .A2(new_n471), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n949), .A2(new_n955), .A3(new_n314), .A4(new_n950), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT123), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n954), .A2(new_n958), .A3(new_n959), .ZN(G1349gat));
  NAND2_X1  g759(.A1(new_n495), .A2(new_n497), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n961), .A3(new_n246), .ZN(new_n962));
  INV_X1    g761(.A(new_n725), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n949), .A2(new_n963), .A3(new_n950), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n964), .B2(G183gat), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT124), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(KEYINPUT60), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n965), .B(new_n967), .ZN(G1350gat));
  NAND3_X1  g767(.A1(new_n945), .A2(new_n498), .A3(new_n296), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n949), .A2(new_n296), .A3(new_n950), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n971));
  AND3_X1   g770(.A1(new_n970), .A2(new_n971), .A3(G190gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n971), .B1(new_n970), .B2(G190gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n969), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n646), .A2(new_n700), .A3(new_n631), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n926), .B(new_n977), .C1(new_n917), .C2(new_n909), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n342), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n909), .A2(new_n976), .ZN(new_n981));
  INV_X1    g780(.A(G197gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n981), .A2(new_n982), .A3(new_n728), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n983), .B(KEYINPUT125), .Z(new_n984));
  NAND2_X1  g783(.A1(new_n980), .A2(new_n984), .ZN(G1352gat));
  OAI21_X1  g784(.A(G204gat), .B1(new_n979), .B2(new_n315), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n315), .A2(G204gat), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n981), .A2(new_n987), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n986), .A2(new_n992), .ZN(G1353gat));
  INV_X1    g792(.A(G211gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n981), .A2(new_n994), .A3(new_n718), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n718), .A2(new_n976), .ZN(new_n996));
  OAI21_X1  g795(.A(G211gat), .B1(new_n927), .B2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n995), .B1(new_n999), .B2(new_n1000), .ZN(G1354gat));
  AOI21_X1  g800(.A(G218gat), .B1(new_n981), .B2(new_n296), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n348), .A2(new_n350), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n979), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g803(.A(new_n1002), .B1(new_n1004), .B2(new_n296), .ZN(G1355gat));
endmodule


