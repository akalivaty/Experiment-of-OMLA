//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n567, new_n568, new_n569, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n632,
    new_n634, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G234));
  NAND2_X1  g025(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT66), .Z(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n464), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n468), .A2(G136), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(new_n469), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n473), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G162));
  OR2_X1    g054(.A1(new_n462), .A2(new_n463), .ZN(new_n480));
  AND2_X1   g055(.A1(G126), .A2(G2105), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n480), .A2(KEYINPUT67), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n481), .B1(new_n462), .B2(new_n463), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(KEYINPUT68), .A2(G114), .ZN(new_n486));
  NOR2_X1   g061(.A1(KEYINPUT68), .A2(G114), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n482), .A2(new_n485), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n469), .C1(new_n462), .C2(new_n463), .ZN(new_n492));
  XNOR2_X1  g067(.A(new_n492), .B(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(G75), .A2(G543), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n502), .A2(new_n503), .B1(KEYINPUT5), .B2(new_n497), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT71), .B1(new_n505), .B2(new_n497), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n496), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(G50), .A2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OAI21_X1  g089(.A(KEYINPUT69), .B1(new_n514), .B2(G651), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT6), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n515), .A2(new_n518), .B1(new_n514), .B2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n510), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n498), .A2(KEYINPUT70), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n503), .B(G543), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n506), .A2(new_n523), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n528), .B(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n514), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n516), .B1(KEYINPUT6), .B2(new_n517), .ZN(new_n532));
  NOR3_X1   g107(.A1(new_n514), .A2(KEYINPUT69), .A3(G651), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT73), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n536), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n535), .A2(G51), .A3(G543), .A4(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n504), .A2(new_n506), .A3(new_n519), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n538), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n530), .A2(new_n543), .ZN(G168));
  NAND2_X1  g119(.A1(G77), .A2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n507), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n535), .A2(G52), .A3(G543), .A4(new_n537), .ZN(new_n549));
  NAND4_X1  g124(.A1(new_n504), .A2(G90), .A3(new_n506), .A4(new_n519), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n551), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n548), .B1(new_n553), .B2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  XNOR2_X1  g131(.A(KEYINPUT75), .B(G43), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n535), .A2(G543), .A3(new_n537), .A4(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n504), .A2(G81), .A3(new_n506), .A4(new_n519), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n506), .A2(G56), .A3(new_n526), .A4(new_n523), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n517), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g144(.A(new_n569), .B(KEYINPUT76), .Z(G188));
  NAND4_X1  g145(.A1(new_n535), .A2(G53), .A3(G543), .A4(new_n537), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  XOR2_X1   g148(.A(new_n573), .B(KEYINPUT77), .Z(new_n574));
  XOR2_X1   g149(.A(KEYINPUT78), .B(G65), .Z(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n507), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n542), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(G651), .B1(new_n577), .B2(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n572), .A2(new_n578), .ZN(G299));
  XNOR2_X1  g154(.A(new_n528), .B(KEYINPUT72), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(G89), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n580), .A2(new_n581), .A3(new_n538), .A4(new_n540), .ZN(G286));
  XOR2_X1   g157(.A(new_n521), .B(KEYINPUT79), .Z(G303));
  AND2_X1   g158(.A1(new_n504), .A2(new_n506), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n584), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n577), .A2(G87), .ZN(new_n586));
  AND3_X1   g161(.A1(new_n535), .A2(G543), .A3(new_n537), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(G49), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT80), .Z(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n507), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g168(.A1(G48), .A2(G543), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n593), .A2(G651), .B1(new_n519), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n577), .A2(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(KEYINPUT81), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT81), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n577), .A2(new_n598), .A3(G86), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n595), .A2(new_n597), .A3(new_n599), .ZN(G305));
  NAND3_X1  g175(.A1(new_n535), .A2(G543), .A3(new_n537), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n601), .A2(new_n602), .B1(new_n542), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n507), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n577), .A2(G92), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n612), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n542), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n613), .A2(new_n616), .B1(G54), .B2(new_n587), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n504), .A2(G66), .A3(new_n506), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT83), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n618), .A2(KEYINPUT83), .A3(new_n619), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n622), .A2(G651), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n611), .B1(new_n626), .B2(G868), .ZN(G284));
  OAI21_X1  g202(.A(new_n611), .B1(new_n626), .B2(G868), .ZN(G321));
  XOR2_X1   g203(.A(G299), .B(KEYINPUT84), .Z(new_n629));
  MUX2_X1   g204(.A(new_n629), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g205(.A(new_n629), .B(G286), .S(G868), .Z(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n626), .B1(new_n632), .B2(G860), .ZN(G148));
  OAI21_X1  g208(.A(G868), .B1(new_n625), .B2(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n564), .ZN(G323));
  XOR2_X1   g210(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n636));
  XNOR2_X1  g211(.A(G323), .B(new_n636), .ZN(G282));
  NAND2_X1  g212(.A1(new_n480), .A2(new_n470), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT12), .Z(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT13), .Z(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n468), .A2(G135), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n474), .A2(G123), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n469), .A2(G111), .ZN(new_n646));
  OAI21_X1  g221(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n645), .C1(new_n646), .C2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT86), .ZN(G156));
  INV_X1    g226(.A(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2427), .B(G2438), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n652), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n655), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1341), .B(G1348), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2443), .B(G2446), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(G14), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(G401));
  XNOR2_X1  g242(.A(G2072), .B(G2078), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n669), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT87), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n675), .B(new_n672), .C1(new_n668), .C2(new_n670), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n671), .A2(new_n668), .A3(new_n670), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G2096), .B(G2100), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n679), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G227));
  XNOR2_X1  g258(.A(G1971), .B(G1976), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT19), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(G1956), .B(G2474), .Z(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  AND2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(new_n686), .B2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G160), .ZN(new_n702));
  INV_X1    g277(.A(G29), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT24), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n704), .A2(G34), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n703), .B1(new_n704), .B2(G34), .ZN(new_n706));
  OAI22_X1  g281(.A1(new_n702), .A2(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT25), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n468), .A2(G139), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n480), .A2(G127), .ZN(new_n717));
  NAND2_X1  g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n469), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n720), .A2(new_n703), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n703), .B2(G33), .ZN(new_n722));
  INV_X1    g297(.A(G2072), .ZN(new_n723));
  OAI211_X1 g298(.A(new_n709), .B(new_n710), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n703), .A2(G35), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G162), .B2(new_n703), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT29), .Z(new_n727));
  INV_X1    g302(.A(G2090), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G19), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n564), .B2(G16), .ZN(new_n731));
  OAI221_X1 g306(.A(new_n729), .B1(G1341), .B2(new_n731), .C1(new_n728), .C2(new_n727), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n468), .A2(G141), .B1(G105), .B2(new_n470), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n474), .A2(G129), .ZN(new_n734));
  NAND3_X1  g309(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT26), .Z(new_n736));
  NAND3_X1  g311(.A1(new_n733), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G29), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G32), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(KEYINPUT95), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(KEYINPUT95), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT27), .B(G1996), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT30), .B(G28), .ZN(new_n749));
  OR2_X1    g324(.A1(KEYINPUT31), .A2(G11), .ZN(new_n750));
  NAND2_X1  g325(.A1(KEYINPUT31), .A2(G11), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n749), .A2(new_n703), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n648), .B2(new_n703), .ZN(new_n753));
  NOR2_X1   g328(.A1(G27), .A2(G29), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G164), .B2(G29), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G2078), .ZN(new_n756));
  AOI211_X1 g331(.A(new_n753), .B(new_n756), .C1(new_n723), .C2(new_n722), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n703), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NAND2_X1  g334(.A1(new_n468), .A2(G140), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n474), .A2(G128), .ZN(new_n761));
  OR2_X1    g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n762), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(G2078), .B2(new_n755), .ZN(new_n768));
  NAND4_X1  g343(.A1(new_n747), .A2(new_n748), .A3(new_n757), .A4(new_n768), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n732), .B(new_n769), .C1(G1341), .C2(new_n731), .ZN(new_n770));
  INV_X1    g345(.A(G16), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G20), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT23), .Z(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G299), .B2(G16), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G1956), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(G21), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G168), .B2(new_n771), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1966), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n775), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(G4), .A2(G16), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(new_n626), .B2(G16), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT93), .B(G1348), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n770), .A2(new_n779), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G1961), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n771), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n771), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT96), .Z(new_n788));
  AOI21_X1  g363(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n771), .A2(G23), .ZN(new_n790));
  INV_X1    g365(.A(new_n589), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n771), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT33), .B(G1976), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n771), .A2(G22), .ZN(new_n795));
  XOR2_X1   g370(.A(new_n795), .B(KEYINPUT92), .Z(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n771), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G1971), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(G1971), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT32), .B(G1981), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT34), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n703), .A2(G25), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT89), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n468), .A2(G131), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n474), .A2(G119), .ZN(new_n809));
  OR2_X1    g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n810), .B(G2104), .C1(G107), .C2(new_n469), .ZN(new_n811));
  AND3_X1   g386(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n812), .A2(KEYINPUT90), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(KEYINPUT90), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n807), .B1(new_n815), .B2(G29), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n771), .A2(G24), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n604), .B1(new_n608), .B2(G651), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n821), .B2(new_n771), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT91), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1986), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n805), .A2(new_n819), .A3(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT36), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n788), .A2(new_n785), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT97), .ZN(new_n828));
  AND3_X1   g403(.A1(new_n789), .A2(new_n826), .A3(new_n828), .ZN(G311));
  NAND3_X1  g404(.A1(new_n789), .A2(new_n826), .A3(new_n828), .ZN(G150));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(new_n560), .B2(new_n563), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n506), .A2(G67), .A3(new_n526), .A4(new_n523), .ZN(new_n833));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G651), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n535), .A2(G55), .A3(G543), .A4(new_n537), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n504), .A2(G93), .A3(new_n506), .A4(new_n519), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT99), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n564), .B2(KEYINPUT98), .ZN(new_n842));
  NOR4_X1   g417(.A1(new_n560), .A2(new_n563), .A3(new_n831), .A4(KEYINPUT99), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n840), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n561), .A2(new_n562), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G651), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n846), .A2(KEYINPUT98), .A3(new_n559), .A4(new_n558), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT99), .ZN(new_n848));
  INV_X1    g423(.A(new_n560), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n849), .A2(KEYINPUT98), .A3(new_n841), .A4(new_n846), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n848), .A2(new_n839), .A3(new_n832), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT38), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n625), .A2(new_n632), .ZN(new_n854));
  XOR2_X1   g429(.A(new_n853), .B(new_n854), .Z(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT100), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n839), .A2(G860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n861), .B(KEYINPUT37), .Z(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  XOR2_X1   g438(.A(G160), .B(new_n648), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n478), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n813), .A2(new_n814), .A3(KEYINPUT102), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT102), .B1(new_n813), .B2(new_n814), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n639), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n474), .A2(G130), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n468), .A2(G142), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n874));
  OR3_X1    g449(.A1(new_n874), .A2(new_n469), .A3(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n874), .B1(new_n469), .B2(G118), .ZN(new_n876));
  OR2_X1    g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n875), .A2(G2104), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n873), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n815), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n639), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(new_n883), .A3(new_n868), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n871), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n880), .B1(new_n871), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n867), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n871), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n879), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(KEYINPUT103), .A3(new_n885), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n740), .A2(new_n764), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n740), .A2(new_n764), .ZN(new_n895));
  OAI21_X1  g470(.A(G164), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n897), .A2(new_n494), .A3(new_n893), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n720), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n898), .A3(new_n720), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n888), .A2(new_n891), .A3(new_n902), .A4(new_n901), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n866), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n886), .A2(new_n887), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n866), .B1(new_n903), .B2(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n888), .A2(new_n891), .B1(new_n902), .B2(new_n901), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g487(.A(new_n912), .B(KEYINPUT40), .Z(G395));
  NOR2_X1   g488(.A1(new_n625), .A2(G559), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n852), .B(new_n914), .Z(new_n915));
  NAND2_X1  g490(.A1(new_n613), .A2(new_n616), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n587), .A2(G54), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n622), .A2(G651), .A3(new_n623), .ZN(new_n919));
  OAI21_X1  g494(.A(G299), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n617), .A2(new_n624), .A3(new_n572), .A4(new_n578), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT41), .B1(new_n920), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n915), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n921), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n915), .ZN(new_n927));
  XNOR2_X1  g502(.A(G305), .B(new_n521), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n791), .A2(new_n821), .ZN(new_n929));
  NAND2_X1  g504(.A1(G290), .A2(new_n589), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT104), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT104), .B1(new_n929), .B2(new_n930), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n928), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n928), .A2(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(new_n937), .B(KEYINPUT42), .Z(new_n938));
  XNOR2_X1  g513(.A(new_n927), .B(new_n938), .ZN(new_n939));
  MUX2_X1   g514(.A(new_n839), .B(new_n939), .S(G868), .Z(G295));
  MUX2_X1   g515(.A(new_n839), .B(new_n939), .S(G868), .Z(G331));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n942));
  NAND2_X1  g517(.A1(G301), .A2(G286), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n549), .A2(new_n550), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT74), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n552), .ZN(new_n946));
  NAND3_X1  g521(.A1(G168), .A2(new_n946), .A3(new_n548), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n842), .A2(new_n840), .A3(new_n843), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n848), .A2(new_n850), .B1(new_n839), .B2(new_n832), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n844), .A2(new_n851), .A3(new_n943), .A4(new_n947), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n948), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(KEYINPUT105), .A3(new_n851), .A4(new_n844), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n924), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n951), .A2(KEYINPUT106), .ZN(new_n958));
  INV_X1    g533(.A(new_n926), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT106), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n852), .A2(new_n960), .A3(new_n948), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n958), .A2(new_n959), .A3(new_n953), .A4(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n962), .A3(new_n937), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT107), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n957), .A2(new_n962), .A3(new_n937), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n954), .A2(new_n956), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n958), .A2(new_n953), .A3(new_n961), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n959), .A2(new_n968), .B1(new_n969), .B2(new_n924), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT108), .B1(new_n970), .B2(new_n937), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT108), .ZN(new_n972));
  INV_X1    g547(.A(new_n937), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n969), .A2(new_n924), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n926), .B1(new_n954), .B2(new_n956), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n972), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n967), .A2(new_n971), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT43), .B1(new_n977), .B2(G37), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n957), .A2(new_n962), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n979), .B2(new_n973), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n967), .A2(new_n980), .ZN(new_n981));
  OR2_X1    g556(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n942), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n981), .A2(KEYINPUT43), .ZN(new_n984));
  NOR2_X1   g559(.A1(KEYINPUT43), .A2(G37), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n967), .A2(new_n971), .A3(new_n976), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT44), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n983), .A2(new_n988), .ZN(G397));
  AND3_X1   g564(.A1(new_n467), .A2(new_n471), .A3(G40), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n491), .B2(new_n493), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n991), .A2(KEYINPUT45), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1996), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT109), .Z(new_n996));
  XOR2_X1   g571(.A(new_n996), .B(KEYINPUT46), .Z(new_n997));
  XNOR2_X1  g572(.A(new_n764), .B(G2067), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n740), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n998), .B1(new_n740), .B2(G1996), .ZN(new_n1002));
  INV_X1    g577(.A(new_n993), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n996), .B2(new_n741), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n815), .A2(new_n818), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n764), .A2(G2067), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n993), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1001), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n817), .B1(new_n813), .B2(new_n814), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n993), .B1(new_n1006), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1005), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT126), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  INV_X1    g591(.A(G1986), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n993), .A2(new_n821), .A3(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(new_n1018), .B(KEYINPUT48), .Z(new_n1019));
  NOR2_X1   g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1010), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(G305), .A2(G1981), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n595), .A2(new_n596), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(G1981), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT49), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n992), .A2(new_n990), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G8), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1024), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n791), .B2(G1976), .ZN(new_n1032));
  INV_X1    g607(.A(G1976), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G288), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1031), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1032), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1035), .A2(KEYINPUT111), .ZN(new_n1038));
  OAI221_X1 g613(.A(new_n1030), .B1(new_n1031), .B2(new_n1032), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n990), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT116), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n990), .B(KEYINPUT116), .C1(new_n992), .C2(KEYINPUT45), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1966), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n992), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n990), .B1(new_n992), .B2(new_n1048), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n708), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1047), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G8), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G286), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G303), .A2(G8), .ZN(new_n1057));
  XOR2_X1   g632(.A(new_n1057), .B(KEYINPUT55), .Z(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1052), .A2(new_n728), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT110), .B(G1971), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1043), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n1040), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1059), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1056), .B1(new_n1058), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n1065), .ZN(new_n1066));
  AOI211_X1 g641(.A(G1976), .B(G288), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1067));
  XNOR2_X1  g642(.A(new_n1022), .B(KEYINPUT112), .ZN(new_n1068));
  OAI211_X1 g643(.A(G8), .B(new_n1026), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(new_n1064), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1066), .B(new_n1069), .C1(new_n1039), .C2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(G168), .A2(KEYINPUT121), .A3(new_n1059), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT121), .B1(G168), .B2(new_n1059), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT121), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(G286), .B2(G8), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT122), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1059), .B1(new_n1047), .B2(new_n1053), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT51), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1072), .A2(new_n1078), .A3(KEYINPUT51), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1055), .A2(KEYINPUT123), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  OR3_X1    g660(.A1(new_n1072), .A2(new_n1078), .A3(KEYINPUT51), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1085), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(new_n1084), .A3(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1054), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT62), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1092), .A3(new_n1089), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n785), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1094));
  INV_X1    g669(.A(G2078), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1045), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1062), .A2(new_n1040), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT53), .B1(new_n1098), .B2(new_n1095), .ZN(new_n1099));
  OAI21_X1  g674(.A(G171), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1091), .A2(new_n1093), .A3(new_n1101), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1055), .A2(KEYINPUT63), .A3(G286), .ZN(new_n1103));
  XNOR2_X1  g678(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(G299), .B(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1051), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT113), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1049), .A2(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT113), .B1(new_n992), .B2(new_n1048), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT117), .B(G1956), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(KEYINPUT56), .B(G2072), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1098), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1105), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1105), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1052), .A2(G1348), .B1(G2067), .B2(new_n1026), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n626), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1117), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1120), .A2(new_n1116), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1121), .A2(KEYINPUT60), .A3(new_n625), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1121), .B(new_n626), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1127), .B1(new_n1128), .B2(KEYINPUT60), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1120), .A2(new_n1116), .A3(KEYINPUT61), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1126), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(KEYINPUT58), .B(G1341), .Z(new_n1132));
  NAND2_X1  g707(.A1(new_n1026), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT119), .B1(new_n1098), .B2(new_n994), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n1135));
  NOR4_X1   g710(.A1(new_n1062), .A2(new_n1040), .A3(new_n1135), .A4(G1996), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g714(.A(KEYINPUT120), .B(new_n1133), .C1(new_n1134), .C2(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT59), .B1(new_n1141), .B2(new_n564), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1131), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1141), .A2(KEYINPUT59), .A3(new_n564), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1123), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1097), .A2(G171), .A3(new_n1099), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT54), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1098), .A2(KEYINPUT53), .A3(new_n1095), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1094), .ZN(new_n1151));
  OAI21_X1  g726(.A(KEYINPUT124), .B1(new_n1151), .B2(new_n1099), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1099), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n1094), .A4(new_n1150), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1149), .B1(new_n1156), .B2(G171), .ZN(new_n1157));
  AOI211_X1 g732(.A(KEYINPUT125), .B(G301), .C1(new_n1152), .C2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1148), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n1151), .A2(G171), .A3(new_n1099), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1147), .B1(new_n1101), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1159), .A2(new_n1090), .A3(new_n1161), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1102), .B(new_n1103), .C1(new_n1145), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(G2090), .B1(new_n1110), .B2(KEYINPUT114), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1164), .B1(KEYINPUT114), .B2(new_n1110), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1059), .B1(new_n1165), .B2(new_n1063), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1070), .B1(new_n1058), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT115), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1039), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1039), .A2(new_n1168), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1167), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1071), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g747(.A(G290), .B(new_n1017), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1013), .B1(new_n1003), .B2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1021), .B1(new_n1172), .B2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1177));
  OAI211_X1 g751(.A(new_n682), .B(G319), .C1(new_n666), .C2(new_n665), .ZN(new_n1178));
  NOR2_X1   g752(.A1(G229), .A2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n906), .B2(new_n911), .ZN(new_n1180));
  INV_X1    g754(.A(new_n1180), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1177), .B1(new_n987), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g756(.A(KEYINPUT127), .B(new_n1180), .C1(new_n984), .C2(new_n986), .ZN(new_n1183));
  NOR2_X1   g757(.A1(new_n1182), .A2(new_n1183), .ZN(G308));
  NAND2_X1  g758(.A1(new_n987), .A2(new_n1181), .ZN(G225));
endmodule


