//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n629, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NAND4_X1  g030(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT67), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(G325), .B(KEYINPUT68), .Z(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND4_X1  g041(.A1(new_n463), .A2(new_n465), .A3(G137), .A4(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT69), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  XNOR2_X1  g044(.A(KEYINPUT3), .B(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(KEYINPUT69), .A3(G137), .A4(new_n466), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n463), .A2(new_n465), .ZN(new_n474));
  INV_X1    g049(.A(G125), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G101), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n470), .A2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n474), .A2(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G112), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n462), .B1(new_n487), .B2(G2105), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n485), .A2(G136), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n490), .B(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n465), .A3(G126), .A4(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT72), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g075(.A1(new_n463), .A2(new_n465), .A3(G138), .A4(new_n466), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n470), .A2(KEYINPUT4), .A3(G138), .A4(new_n466), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n493), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n500), .A2(new_n503), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AOI21_X1  g082(.A(KEYINPUT5), .B1(KEYINPUT75), .B2(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT74), .A2(G543), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g085(.A1(KEYINPUT74), .A2(KEYINPUT75), .A3(KEYINPUT5), .A4(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n517), .B1(new_n514), .B2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n519), .A2(KEYINPUT6), .A3(G651), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n520), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n515), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND2_X1  g103(.A1(new_n521), .A2(G51), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(KEYINPUT78), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n512), .A2(new_n523), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n512), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT76), .B1(new_n512), .B2(new_n534), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n529), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT77), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT7), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(KEYINPUT79), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n535), .B(new_n536), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT79), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n533), .A2(new_n529), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n542), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G168));
  AOI22_X1  g124(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n514), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n521), .A2(G52), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n524), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  AND2_X1   g131(.A1(new_n510), .A2(new_n511), .ZN(new_n557));
  INV_X1    g132(.A(G56), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n559), .A2(KEYINPUT80), .A3(G651), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n562), .B2(new_n514), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n512), .A2(new_n523), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G81), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n521), .A2(G43), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(G153));
  AND3_X1   g145(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G36), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n571), .A2(new_n574), .ZN(G188));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n523), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n521), .A2(KEYINPUT9), .A3(G53), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT81), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n557), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n565), .B2(G91), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n579), .A2(new_n587), .A3(new_n580), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n582), .A2(new_n586), .A3(new_n588), .ZN(G299));
  INV_X1    g164(.A(G171), .ZN(G301));
  INV_X1    g165(.A(G168), .ZN(G286));
  NAND2_X1  g166(.A1(new_n565), .A2(G87), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT82), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n521), .A2(G49), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  AOI22_X1  g172(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n599), .A2(KEYINPUT83), .A3(G651), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT83), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n598), .B2(new_n514), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n521), .A2(G48), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n565), .A2(G86), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n607), .A2(KEYINPUT84), .A3(new_n514), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT84), .B1(new_n607), .B2(new_n514), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n608), .A2(new_n609), .B1(G47), .B2(new_n521), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n565), .A2(G85), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(G290));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(G92), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n524), .B2(new_n614), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n512), .A2(KEYINPUT10), .A3(G92), .A4(new_n523), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(new_n514), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n521), .A2(G54), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n622), .B2(G171), .ZN(G284));
  OAI21_X1  g199(.A(new_n623), .B1(new_n622), .B2(G171), .ZN(G321));
  NAND2_X1  g200(.A1(G299), .A2(new_n622), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G168), .B2(new_n622), .ZN(G297));
  OAI21_X1  g202(.A(new_n626), .B1(G168), .B2(new_n622), .ZN(G280));
  AND3_X1   g203(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n629));
  INV_X1    g204(.A(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G860), .ZN(G148));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(G868), .B2(new_n569), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n470), .A2(new_n478), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(KEYINPUT12), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n483), .A2(G123), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n485), .A2(G135), .ZN(new_n641));
  NOR2_X1   g216(.A1(G99), .A2(G2105), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2096), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT85), .Z(G156));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XOR2_X1   g224(.A(G2443), .B(G2446), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XOR2_X1   g230(.A(KEYINPUT15), .B(G2435), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n653), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(G14), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  XNOR2_X1  g237(.A(G2072), .B(G2078), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT17), .ZN(new_n664));
  XOR2_X1   g239(.A(G2067), .B(G2678), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n662), .B1(new_n664), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n663), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT87), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n662), .A3(new_n663), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  INV_X1    g246(.A(new_n664), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n672), .A2(new_n662), .A3(new_n665), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(KEYINPUT89), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1971), .B(G1976), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n686), .B(new_n687), .Z(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(new_n685), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT20), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n678), .A2(new_n680), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  OR3_X1    g268(.A1(new_n689), .A2(new_n682), .A3(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT90), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n695), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1986), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n699), .B(new_n702), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G21), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G168), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1966), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT25), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n485), .A2(G139), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n470), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n710), .B(new_n711), .C1(new_n466), .C2(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G33), .B(new_n713), .S(G29), .Z(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT96), .Z(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT97), .A2(G2072), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NOR2_X1   g292(.A1(KEYINPUT97), .A2(G2072), .ZN(new_n718));
  AND2_X1   g293(.A1(KEYINPUT24), .A2(G34), .ZN(new_n719));
  NOR2_X1   g294(.A1(KEYINPUT24), .A2(G34), .ZN(new_n720));
  NOR3_X1   g295(.A1(new_n719), .A2(new_n720), .A3(G29), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(new_n480), .B2(G29), .ZN(new_n722));
  INV_X1    g297(.A(G2084), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n483), .A2(G129), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT98), .B(KEYINPUT26), .Z(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n725), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G29), .B2(G32), .ZN(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  AOI211_X1 g308(.A(new_n718), .B(new_n724), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n717), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT99), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2090), .ZN(new_n738));
  NOR2_X1   g313(.A1(G29), .A2(G35), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G162), .B2(G29), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n737), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n569), .A2(new_n705), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(new_n705), .B2(G19), .ZN(new_n745));
  INV_X1    g320(.A(G1341), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI22_X1  g322(.A1(new_n742), .A2(new_n738), .B1(new_n746), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n732), .A2(new_n733), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n705), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n629), .B2(new_n705), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT93), .B(G1348), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(G2078), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(G171), .A2(G16), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G5), .B2(G16), .ZN(new_n761));
  INV_X1    g336(.A(G1961), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT103), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT100), .B(G28), .ZN(new_n765));
  INV_X1    g340(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(G29), .B1(new_n766), .B2(KEYINPUT30), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT101), .Z(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(KEYINPUT30), .B2(new_n766), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT31), .B(G11), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n769), .B(new_n770), .C1(new_n754), .C2(new_n644), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT102), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n754), .A2(G26), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n483), .A2(G128), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n485), .A2(G140), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n466), .A2(G116), .ZN(new_n778));
  OR3_X1    g353(.A1(KEYINPUT94), .A2(G104), .A3(G2105), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT94), .B1(G104), .B2(G2105), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n779), .A2(G2104), .A3(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n776), .B(new_n777), .C1(new_n778), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2067), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n761), .A2(new_n762), .B1(new_n723), .B2(new_n722), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n764), .A2(new_n772), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n748), .A2(new_n749), .A3(new_n759), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n705), .A2(G20), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n582), .A2(new_n586), .A3(new_n588), .ZN(new_n789));
  OAI211_X1 g364(.A(KEYINPUT23), .B(new_n788), .C1(new_n789), .C2(new_n705), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(KEYINPUT23), .B2(new_n788), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1956), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n743), .A2(new_n747), .A3(new_n787), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n705), .A2(G23), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G288), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT33), .ZN(new_n796));
  INV_X1    g371(.A(G1976), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G305), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n705), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G6), .B2(new_n705), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT32), .B(G1981), .Z(new_n802));
  AND2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NOR2_X1   g379(.A1(G166), .A2(new_n705), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n705), .B2(G22), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR3_X1   g383(.A1(new_n803), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n807), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n798), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  INV_X1    g387(.A(G290), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(new_n705), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n705), .B2(G24), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n483), .A2(G119), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(KEYINPUT92), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(KEYINPUT92), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n820), .A2(new_n821), .B1(G131), .B2(new_n485), .ZN(new_n822));
  OR2_X1    g397(.A1(G95), .A2(G2105), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n823), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(G29), .Z(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT35), .B(G1991), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n815), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(G1986), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n812), .A2(new_n817), .A3(new_n818), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(KEYINPUT36), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n818), .A2(new_n830), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n833), .A2(new_n834), .A3(new_n817), .A4(new_n812), .ZN(new_n835));
  AOI211_X1 g410(.A(new_n708), .B(new_n793), .C1(new_n832), .C2(new_n835), .ZN(G311));
  AOI21_X1  g411(.A(new_n793), .B1(new_n832), .B2(new_n835), .ZN(new_n837));
  INV_X1    g412(.A(new_n708), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  AOI22_X1  g414(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n840), .A2(new_n514), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n521), .A2(G55), .ZN(new_n842));
  INV_X1    g417(.A(G93), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n524), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT104), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n568), .A2(new_n845), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n846), .A2(new_n564), .A3(new_n566), .A4(new_n567), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT39), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n629), .A2(G559), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT38), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n853), .B(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n849), .B1(new_n856), .B2(G860), .ZN(G145));
  XNOR2_X1  g432(.A(new_n782), .B(new_n713), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n503), .A2(new_n504), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT105), .B1(new_n859), .B2(new_n498), .ZN(new_n860));
  INV_X1    g435(.A(new_n498), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n861), .A2(new_n862), .A3(new_n503), .A4(new_n504), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n730), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n858), .A2(new_n864), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n782), .B(new_n713), .Z(new_n870));
  INV_X1    g445(.A(new_n864), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n730), .B1(new_n872), .B2(new_n865), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n483), .A2(G130), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n877));
  AND2_X1   g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n485), .A2(G142), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT106), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n822), .B2(new_n824), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT107), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n822), .A2(new_n824), .A3(new_n881), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n822), .A2(new_n824), .A3(new_n881), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT107), .B1(new_n887), .B2(new_n882), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n886), .A2(new_n637), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n637), .B1(new_n886), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n874), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n886), .A2(new_n888), .ZN(new_n892));
  INV_X1    g467(.A(new_n637), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n886), .A2(new_n888), .A3(new_n637), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n867), .B1(new_n866), .B2(new_n868), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n872), .A2(new_n730), .A3(new_n865), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(new_n899), .A3(KEYINPUT108), .ZN(new_n900));
  XNOR2_X1  g475(.A(G162), .B(new_n644), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n480), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT108), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n894), .A2(new_n898), .A3(new_n904), .A4(new_n895), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(G37), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n891), .A2(new_n899), .A3(new_n902), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g485(.A1(new_n846), .A2(G868), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(G303), .ZN(new_n913));
  NAND2_X1  g488(.A1(G288), .A2(G166), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n913), .A2(G305), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(G305), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  OAI21_X1  g492(.A(G290), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(new_n799), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n920), .A2(new_n813), .A3(new_n915), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g497(.A1(new_n922), .A2(KEYINPUT110), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(KEYINPUT42), .A3(new_n924), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n852), .B(new_n632), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n789), .A2(new_n629), .ZN(new_n931));
  NAND2_X1  g506(.A1(G299), .A2(new_n621), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n932), .ZN(new_n936));
  NOR2_X1   g511(.A1(G299), .A2(new_n621), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT41), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n931), .A2(new_n939), .A3(new_n932), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT109), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n931), .A2(new_n939), .A3(new_n932), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT109), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n935), .B1(new_n945), .B2(new_n930), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n929), .A2(KEYINPUT111), .A3(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n946), .A2(KEYINPUT111), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(KEYINPUT111), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n927), .A2(new_n928), .A3(new_n948), .A4(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n911), .B1(new_n951), .B2(G868), .ZN(G295));
  AOI21_X1  g527(.A(new_n911), .B1(new_n951), .B2(G868), .ZN(G331));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n850), .A2(G168), .A3(new_n851), .ZN(new_n955));
  AOI21_X1  g530(.A(G168), .B1(new_n850), .B2(new_n851), .ZN(new_n956));
  OAI21_X1  g531(.A(G301), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n852), .A2(G286), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n850), .A2(G168), .A3(new_n851), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(G171), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT112), .B1(new_n945), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n936), .A2(KEYINPUT41), .A3(new_n937), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n939), .B1(new_n931), .B2(new_n932), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n943), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n968), .A3(new_n960), .A4(new_n957), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n961), .A2(new_n934), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n962), .A2(new_n969), .A3(new_n922), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n907), .ZN(new_n972));
  INV_X1    g547(.A(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n922), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n961), .B1(new_n940), .B2(new_n938), .ZN(new_n975));
  INV_X1    g550(.A(new_n970), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n954), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n962), .A2(new_n969), .A3(new_n970), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n979), .A2(new_n974), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n980), .A2(new_n972), .A3(KEYINPUT43), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n982));
  OR3_X1    g557(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n980), .B2(new_n972), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n977), .A2(new_n971), .A3(new_n954), .A4(new_n907), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(new_n982), .ZN(new_n988));
  AOI211_X1 g563(.A(KEYINPUT113), .B(KEYINPUT44), .C1(new_n985), .C2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(G397));
  AOI21_X1  g565(.A(G1384), .B1(new_n860), .B2(new_n863), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n472), .A2(new_n477), .A3(G40), .A4(new_n479), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n782), .B(G2067), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n995), .A2(new_n996), .A3(KEYINPUT114), .ZN(new_n1000));
  INV_X1    g575(.A(G1996), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n730), .B(new_n1001), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n999), .A2(new_n1000), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n825), .A2(new_n827), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n825), .A2(new_n827), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n995), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(G290), .A2(G1986), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n995), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT48), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n1012));
  INV_X1    g587(.A(new_n995), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(G1996), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n995), .B1(new_n996), .B2(new_n867), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n995), .A2(KEYINPUT46), .A3(new_n1001), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(KEYINPUT47), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n782), .A2(G2067), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1019), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1011), .B(new_n1018), .C1(new_n1013), .C2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(new_n1021), .B(KEYINPUT127), .Z(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n506), .A2(KEYINPUT45), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n994), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1023), .B1(new_n859), .B2(new_n498), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT45), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1025), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G1966), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT120), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n493), .A2(KEYINPUT72), .A3(new_n497), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT72), .B1(new_n493), .B2(new_n497), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n859), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1384), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1033), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1026), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n994), .B1(new_n1041), .B2(new_n1039), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n506), .A2(new_n1023), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT117), .A3(KEYINPUT50), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .A4(new_n723), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT120), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1029), .A2(new_n1046), .A3(new_n1030), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1032), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  NOR2_X1   g625(.A1(G168), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(KEYINPUT51), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(G8), .C1(new_n1048), .C2(G286), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT123), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1048), .A2(KEYINPUT123), .A3(new_n1051), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1053), .B(new_n1055), .C1(new_n1056), .C2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g633(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1059));
  AOI21_X1  g634(.A(new_n994), .B1(new_n991), .B2(KEYINPUT45), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n1043), .B2(new_n1027), .ZN(new_n1062));
  AOI211_X1 g637(.A(KEYINPUT115), .B(KEYINPUT45), .C1(new_n506), .C2(new_n1023), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1060), .B(new_n757), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1040), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1064), .A2(new_n1065), .B1(new_n762), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n993), .A2(new_n1060), .A3(KEYINPUT53), .A4(new_n757), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1067), .A2(G301), .A3(new_n1068), .ZN(new_n1069));
  OR3_X1    g644(.A1(new_n1029), .A2(new_n1065), .A3(G2078), .ZN(new_n1070));
  AOI21_X1  g645(.A(G301), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1059), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(KEYINPUT55), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n1075));
  NAND3_X1  g650(.A1(G303), .A2(new_n1075), .A3(G8), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1025), .B(new_n1078), .C1(new_n1043), .C2(KEYINPUT50), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(G2090), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1060), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1081), .B2(new_n807), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1077), .B1(new_n1082), .B2(new_n1050), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT49), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G305), .A2(G1981), .ZN(new_n1085));
  INV_X1    g660(.A(G1981), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n600), .A2(new_n602), .B1(G86), .B2(new_n565), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n1087), .B2(new_n604), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1084), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1050), .B1(new_n1025), .B2(new_n1041), .ZN(new_n1090));
  NAND2_X1  g665(.A1(G305), .A2(G1981), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n1086), .A3(new_n604), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(KEYINPUT49), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1090), .B1(G288), .B2(new_n797), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT52), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(G288), .B2(new_n797), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(new_n1090), .C1(new_n797), .C2(G288), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1083), .A2(new_n1094), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1025), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n807), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT116), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1066), .A2(G2090), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1081), .A2(new_n1106), .A3(new_n807), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1077), .B(KEYINPUT118), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(G8), .A3(new_n1109), .ZN(new_n1110));
  AND4_X1   g685(.A1(new_n1058), .A2(new_n1072), .A3(new_n1099), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1025), .A2(new_n1041), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1112), .A2(G2067), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n1066), .B2(new_n752), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n629), .B1(new_n1114), .B2(KEYINPUT60), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  AOI211_X1 g691(.A(new_n1116), .B(new_n1113), .C1(new_n1066), .C2(new_n752), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1114), .A2(KEYINPUT60), .A3(new_n621), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1060), .B(new_n1121), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n581), .A2(KEYINPUT57), .ZN(new_n1123));
  AOI22_X1  g698(.A1(G299), .A2(KEYINPUT57), .B1(new_n586), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(G1956), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1079), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1122), .A2(new_n1124), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT61), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1122), .A2(new_n1133), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1132), .A2(new_n1128), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1127), .A2(KEYINPUT61), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT115), .B1(new_n1038), .B2(KEYINPUT45), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1043), .A2(new_n1061), .A3(new_n1027), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1140), .A2(new_n1001), .A3(new_n1060), .ZN(new_n1141));
  XOR2_X1   g716(.A(KEYINPUT58), .B(G1341), .Z(new_n1142));
  NAND2_X1  g717(.A1(new_n1112), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n568), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1144), .B(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1120), .A2(new_n1129), .A3(new_n1137), .A4(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1132), .A2(KEYINPUT121), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1130), .A2(new_n1131), .A3(new_n1149), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1148), .B(new_n1150), .C1(new_n621), .C2(new_n1114), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n1127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G171), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1155), .A2(KEYINPUT125), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1067), .A2(G301), .A3(new_n1070), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(KEYINPUT125), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1156), .A2(KEYINPUT54), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1111), .A2(new_n1153), .A3(new_n1159), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1094), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1049), .A2(G286), .ZN(new_n1162));
  AOI211_X1 g737(.A(KEYINPUT116), .B(G1971), .C1(new_n1140), .C2(new_n1060), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1106), .B1(new_n1081), .B2(new_n807), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1050), .B1(new_n1165), .B2(new_n1105), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1077), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1161), .B(new_n1162), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT63), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1090), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n594), .A2(new_n797), .A3(new_n595), .A4(new_n596), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT119), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1170), .B1(new_n1174), .B2(new_n1092), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1047), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1046), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1050), .B1(new_n1178), .B2(new_n1045), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1083), .A2(new_n1179), .A3(new_n1180), .A4(G168), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1110), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1175), .B1(new_n1182), .B2(new_n1161), .ZN(new_n1183));
  AND2_X1   g758(.A1(new_n1169), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT126), .ZN(new_n1185));
  AND3_X1   g760(.A1(new_n1160), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1160), .B2(new_n1184), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1071), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1099), .A2(new_n1110), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1058), .A2(KEYINPUT62), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1186), .A2(new_n1187), .A3(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n813), .A2(new_n816), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n995), .B1(new_n1194), .B2(new_n1008), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1007), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1022), .B1(new_n1193), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g772(.A1(new_n660), .A2(G319), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n909), .A2(new_n676), .A3(new_n1199), .ZN(new_n1200));
  AND3_X1   g774(.A1(new_n1200), .A2(new_n703), .A3(new_n987), .ZN(G308));
  NAND3_X1  g775(.A1(new_n1200), .A2(new_n703), .A3(new_n987), .ZN(G225));
endmodule


