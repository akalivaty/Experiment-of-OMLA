

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726;

  INV_X1 U376 ( .A(G953), .ZN(n714) );
  INV_X2 U377 ( .A(G143), .ZN(n360) );
  NOR2_X2 U378 ( .A1(n654), .A2(n496), .ZN(n623) );
  OR2_X2 U379 ( .A1(n393), .A2(n392), .ZN(n395) );
  XNOR2_X2 U380 ( .A(n376), .B(n391), .ZN(n393) );
  XOR2_X2 U381 ( .A(KEYINPUT41), .B(n580), .Z(n676) );
  INV_X1 U382 ( .A(KEYINPUT19), .ZN(n365) );
  AND2_X1 U383 ( .A1(n524), .A2(n523), .ZN(n534) );
  AND2_X1 U384 ( .A1(n527), .A2(n526), .ZN(n529) );
  NOR2_X1 U385 ( .A1(n497), .A2(n589), .ZN(n520) );
  BUF_X1 U386 ( .A(n495), .Z(n657) );
  XNOR2_X1 U387 ( .A(n362), .B(G469), .ZN(n545) );
  XNOR2_X1 U388 ( .A(n367), .B(n699), .ZN(n364) );
  NOR2_X1 U389 ( .A1(n623), .A2(n725), .ZN(n528) );
  XNOR2_X1 U390 ( .A(G131), .B(G134), .ZN(n417) );
  XNOR2_X1 U391 ( .A(n459), .B(G472), .ZN(n495) );
  NOR2_X1 U392 ( .A1(n610), .A2(G902), .ZN(n459) );
  NOR2_X1 U393 ( .A1(n688), .A2(G902), .ZN(n362) );
  XNOR2_X1 U394 ( .A(n363), .B(n357), .ZN(n497) );
  XNOR2_X1 U395 ( .A(n578), .B(n577), .ZN(n594) );
  INV_X1 U396 ( .A(KEYINPUT39), .ZN(n577) );
  NOR2_X1 U397 ( .A1(n369), .A2(n576), .ZN(n578) );
  NAND2_X1 U398 ( .A1(n575), .A2(n370), .ZN(n369) );
  INV_X1 U399 ( .A(n651), .ZN(n589) );
  XNOR2_X1 U400 ( .A(n443), .B(n442), .ZN(n444) );
  NOR2_X1 U401 ( .A1(G902), .A2(n695), .ZN(n445) );
  XNOR2_X1 U402 ( .A(n366), .B(n388), .ZN(n699) );
  XNOR2_X1 U403 ( .A(n446), .B(n389), .ZN(n366) );
  NOR2_X1 U404 ( .A1(G952), .A2(n714), .ZN(n698) );
  XOR2_X1 U405 ( .A(KEYINPUT71), .B(KEYINPUT99), .Z(n448) );
  XNOR2_X1 U406 ( .A(KEYINPUT98), .B(KEYINPUT5), .ZN(n447) );
  XNOR2_X1 U407 ( .A(G113), .B(G116), .ZN(n450) );
  NOR2_X1 U408 ( .A1(n573), .A2(n572), .ZN(n584) );
  XNOR2_X1 U409 ( .A(G143), .B(G131), .ZN(n465) );
  XNOR2_X1 U410 ( .A(n419), .B(n418), .ZN(n458) );
  XNOR2_X1 U411 ( .A(n710), .B(G146), .ZN(n418) );
  XOR2_X1 U412 ( .A(KEYINPUT75), .B(G140), .Z(n421) );
  XNOR2_X1 U413 ( .A(n586), .B(n371), .ZN(n640) );
  INV_X1 U414 ( .A(KEYINPUT38), .ZN(n371) );
  NOR2_X1 U415 ( .A1(n640), .A2(n574), .ZN(n370) );
  XNOR2_X1 U416 ( .A(n545), .B(KEYINPUT1), .ZN(n651) );
  NOR2_X1 U417 ( .A1(n651), .A2(n650), .ZN(n512) );
  XNOR2_X1 U418 ( .A(n473), .B(n472), .ZN(n506) );
  XOR2_X1 U419 ( .A(n460), .B(n495), .Z(n518) );
  XNOR2_X1 U420 ( .A(G113), .B(G104), .ZN(n387) );
  XNOR2_X1 U421 ( .A(G110), .B(KEYINPUT73), .ZN(n386) );
  XOR2_X1 U422 ( .A(G116), .B(G107), .Z(n481) );
  XOR2_X1 U423 ( .A(KEYINPUT3), .B(n390), .Z(n446) );
  XOR2_X1 U424 ( .A(G119), .B(KEYINPUT68), .Z(n390) );
  NAND2_X1 U425 ( .A1(n532), .A2(n531), .ZN(n533) );
  OR2_X1 U426 ( .A1(n640), .A2(n641), .ZN(n644) );
  INV_X1 U427 ( .A(KEYINPUT107), .ZN(n507) );
  XNOR2_X1 U428 ( .A(n372), .B(KEYINPUT30), .ZN(n575) );
  XNOR2_X1 U429 ( .A(n610), .B(KEYINPUT62), .ZN(n612) );
  NAND2_X1 U430 ( .A1(n379), .A2(G475), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U432 ( .A(n368), .B(n402), .ZN(n367) );
  NAND2_X1 U433 ( .A1(n395), .A2(n394), .ZN(n368) );
  NAND2_X1 U434 ( .A1(n379), .A2(G210), .ZN(n378) );
  BUF_X1 U435 ( .A(n639), .Z(n675) );
  XNOR2_X1 U436 ( .A(n375), .B(KEYINPUT42), .ZN(n722) );
  XNOR2_X1 U437 ( .A(n374), .B(KEYINPUT40), .ZN(n726) );
  NAND2_X1 U438 ( .A1(n594), .A2(n630), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n504), .B(n503), .ZN(n725) );
  XNOR2_X1 U440 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n503) );
  NAND2_X1 U441 ( .A1(n502), .A2(n354), .ZN(n504) );
  NOR2_X1 U442 ( .A1(n508), .A2(n509), .ZN(n632) );
  XNOR2_X1 U443 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U444 ( .A(n688), .B(n382), .ZN(n691) );
  OR2_X1 U445 ( .A1(n540), .A2(n411), .ZN(n353) );
  XOR2_X1 U446 ( .A(n501), .B(n500), .Z(n354) );
  NOR2_X1 U447 ( .A1(n638), .A2(n595), .ZN(n355) );
  AND2_X1 U448 ( .A1(n353), .A2(n412), .ZN(n356) );
  XOR2_X1 U449 ( .A(KEYINPUT22), .B(KEYINPUT69), .Z(n357) );
  XNOR2_X1 U450 ( .A(KEYINPUT48), .B(KEYINPUT83), .ZN(n358) );
  XNOR2_X1 U451 ( .A(n359), .B(n462), .ZN(n491) );
  NAND2_X1 U452 ( .A1(n639), .A2(n514), .ZN(n359) );
  XNOR2_X2 U453 ( .A(n360), .B(G128), .ZN(n480) );
  NOR2_X2 U454 ( .A1(n586), .A2(n641), .ZN(n407) );
  NAND2_X1 U455 ( .A1(n355), .A2(n361), .ZN(n713) );
  XNOR2_X1 U456 ( .A(n585), .B(n358), .ZN(n361) );
  NOR2_X2 U457 ( .A1(n579), .A2(n644), .ZN(n580) );
  NAND2_X1 U458 ( .A1(n520), .A2(n657), .ZN(n496) );
  NAND2_X1 U459 ( .A1(n514), .A2(n494), .ZN(n363) );
  AND2_X2 U460 ( .A1(n364), .A2(n596), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n364), .B(n683), .ZN(n685) );
  XNOR2_X2 U462 ( .A(n407), .B(n365), .ZN(n546) );
  NOR2_X1 U463 ( .A1(n657), .A2(n641), .ZN(n372) );
  XNOR2_X1 U464 ( .A(n373), .B(n582), .ZN(n583) );
  NAND2_X1 U465 ( .A1(n722), .A2(n726), .ZN(n373) );
  NAND2_X1 U466 ( .A1(n676), .A2(n581), .ZN(n375) );
  XNOR2_X1 U467 ( .A(n376), .B(n710), .ZN(n712) );
  XNOR2_X2 U468 ( .A(n480), .B(KEYINPUT4), .ZN(n376) );
  NOR2_X2 U469 ( .A1(n597), .A2(n596), .ZN(n380) );
  OR2_X1 U470 ( .A1(n597), .A2(n377), .ZN(n601) );
  OR2_X1 U471 ( .A1(n597), .A2(n378), .ZN(n684) );
  INV_X1 U472 ( .A(n596), .ZN(n379) );
  NAND2_X1 U473 ( .A1(n380), .A2(G472), .ZN(n611) );
  NAND2_X1 U474 ( .A1(n380), .A2(G217), .ZN(n694) );
  NAND2_X1 U475 ( .A1(n380), .A2(G478), .ZN(n606) );
  NAND2_X1 U476 ( .A1(n380), .A2(G469), .ZN(n692) );
  NAND2_X1 U477 ( .A1(n546), .A2(n353), .ZN(n414) );
  NAND2_X1 U478 ( .A1(n546), .A2(n356), .ZN(n416) );
  XNOR2_X1 U479 ( .A(n606), .B(n383), .ZN(n608) );
  NOR2_X2 U480 ( .A1(n613), .A2(n698), .ZN(n615) );
  INV_X1 U481 ( .A(n497), .ZN(n502) );
  XOR2_X1 U482 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n381) );
  XOR2_X1 U483 ( .A(n690), .B(n689), .Z(n382) );
  XOR2_X1 U484 ( .A(n605), .B(KEYINPUT122), .Z(n383) );
  XOR2_X1 U485 ( .A(n381), .B(n429), .Z(n384) );
  AND2_X1 U486 ( .A1(G214), .A2(n463), .ZN(n385) );
  XNOR2_X1 U487 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U488 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U489 ( .A(n464), .B(n385), .ZN(n470) );
  XNOR2_X1 U490 ( .A(n461), .B(KEYINPUT33), .ZN(n639) );
  XNOR2_X1 U491 ( .A(n471), .B(G475), .ZN(n472) );
  XNOR2_X1 U492 ( .A(n470), .B(n469), .ZN(n599) );
  INV_X1 U493 ( .A(KEYINPUT34), .ZN(n462) );
  INV_X1 U494 ( .A(n698), .ZN(n607) );
  XNOR2_X1 U495 ( .A(n632), .B(n507), .ZN(n593) );
  INV_X1 U496 ( .A(KEYINPUT63), .ZN(n614) );
  NAND2_X1 U497 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U498 ( .A(n481), .B(KEYINPUT16), .ZN(n389) );
  XNOR2_X1 U499 ( .A(n386), .B(KEYINPUT88), .ZN(n423) );
  XNOR2_X1 U500 ( .A(n387), .B(G122), .ZN(n468) );
  XNOR2_X1 U501 ( .A(n423), .B(n468), .ZN(n388) );
  INV_X1 U502 ( .A(G101), .ZN(n391) );
  INV_X1 U503 ( .A(n393), .ZN(n419) );
  XNOR2_X1 U504 ( .A(G146), .B(G125), .ZN(n392) );
  INV_X1 U505 ( .A(n392), .ZN(n436) );
  NAND2_X1 U506 ( .A1(n393), .A2(n392), .ZN(n394) );
  XOR2_X1 U507 ( .A(KEYINPUT89), .B(KEYINPUT87), .Z(n397) );
  NAND2_X1 U508 ( .A1(G224), .A2(n714), .ZN(n396) );
  XNOR2_X1 U509 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U510 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n399) );
  XNOR2_X1 U511 ( .A(KEYINPUT76), .B(KEYINPUT90), .ZN(n398) );
  XNOR2_X1 U512 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U513 ( .A(n401), .B(n400), .Z(n402) );
  XNOR2_X1 U514 ( .A(G902), .B(KEYINPUT15), .ZN(n596) );
  OR2_X1 U515 ( .A1(G237), .A2(G902), .ZN(n405) );
  AND2_X1 U516 ( .A1(G210), .A2(n405), .ZN(n403) );
  XNOR2_X2 U517 ( .A(n404), .B(n403), .ZN(n586) );
  NAND2_X1 U518 ( .A1(n405), .A2(G214), .ZN(n406) );
  XOR2_X1 U519 ( .A(n406), .B(KEYINPUT91), .Z(n567) );
  INV_X1 U520 ( .A(n567), .ZN(n641) );
  NAND2_X1 U521 ( .A1(G234), .A2(G237), .ZN(n408) );
  XNOR2_X1 U522 ( .A(KEYINPUT14), .B(n408), .ZN(n409) );
  NAND2_X1 U523 ( .A1(G952), .A2(n409), .ZN(n670) );
  NOR2_X1 U524 ( .A1(G953), .A2(n670), .ZN(n540) );
  NAND2_X1 U525 ( .A1(G902), .A2(n409), .ZN(n538) );
  XOR2_X1 U526 ( .A(G898), .B(KEYINPUT92), .Z(n704) );
  NAND2_X1 U527 ( .A1(G953), .A2(n704), .ZN(n701) );
  NOR2_X1 U528 ( .A1(n538), .A2(n701), .ZN(n410) );
  XOR2_X1 U529 ( .A(KEYINPUT93), .B(n410), .Z(n411) );
  XNOR2_X1 U530 ( .A(KEYINPUT86), .B(KEYINPUT0), .ZN(n412) );
  INV_X1 U531 ( .A(n412), .ZN(n413) );
  NAND2_X1 U532 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U533 ( .A1(n416), .A2(n415), .ZN(n514) );
  XNOR2_X1 U534 ( .A(n417), .B(G137), .ZN(n710) );
  NAND2_X1 U535 ( .A1(G227), .A2(n714), .ZN(n420) );
  XNOR2_X1 U536 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U537 ( .A(n422), .B(G104), .Z(n425) );
  XNOR2_X1 U538 ( .A(n423), .B(G107), .ZN(n424) );
  XNOR2_X1 U539 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U540 ( .A(n458), .B(n426), .ZN(n688) );
  NAND2_X1 U541 ( .A1(G234), .A2(n596), .ZN(n427) );
  XNOR2_X1 U542 ( .A(KEYINPUT20), .B(n427), .ZN(n439) );
  NAND2_X1 U543 ( .A1(G221), .A2(n439), .ZN(n428) );
  XOR2_X1 U544 ( .A(n428), .B(KEYINPUT21), .Z(n655) );
  XNOR2_X1 U545 ( .A(G119), .B(KEYINPUT95), .ZN(n429) );
  XOR2_X1 U546 ( .A(KEYINPUT23), .B(G110), .Z(n431) );
  XNOR2_X1 U547 ( .A(G128), .B(G137), .ZN(n430) );
  XNOR2_X1 U548 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U549 ( .A(n384), .B(n432), .ZN(n435) );
  NAND2_X1 U550 ( .A1(G234), .A2(n714), .ZN(n433) );
  XOR2_X1 U551 ( .A(KEYINPUT8), .B(n433), .Z(n484) );
  NAND2_X1 U552 ( .A1(G221), .A2(n484), .ZN(n434) );
  XNOR2_X1 U553 ( .A(n435), .B(n434), .ZN(n438) );
  XNOR2_X1 U554 ( .A(G140), .B(KEYINPUT10), .ZN(n437) );
  XOR2_X1 U555 ( .A(n437), .B(n436), .Z(n464) );
  INV_X1 U556 ( .A(n464), .ZN(n711) );
  XOR2_X1 U557 ( .A(n438), .B(n711), .Z(n695) );
  NAND2_X1 U558 ( .A1(n439), .A2(G217), .ZN(n443) );
  XOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT25), .Z(n441) );
  XNOR2_X1 U560 ( .A(KEYINPUT74), .B(KEYINPUT96), .ZN(n440) );
  XNOR2_X1 U561 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X2 U562 ( .A(n445), .B(n444), .ZN(n654) );
  NAND2_X1 U563 ( .A1(n655), .A2(n654), .ZN(n650) );
  XNOR2_X1 U564 ( .A(KEYINPUT109), .B(KEYINPUT6), .ZN(n460) );
  INV_X1 U565 ( .A(n446), .ZN(n454) );
  XNOR2_X1 U566 ( .A(n448), .B(n447), .ZN(n452) );
  INV_X1 U567 ( .A(KEYINPUT72), .ZN(n449) );
  XNOR2_X1 U568 ( .A(n454), .B(n453), .ZN(n456) );
  NOR2_X1 U569 ( .A1(G953), .A2(G237), .ZN(n463) );
  NAND2_X1 U570 ( .A1(n463), .A2(G210), .ZN(n455) );
  XNOR2_X1 U571 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U572 ( .A(n458), .B(n457), .ZN(n610) );
  NAND2_X1 U573 ( .A1(n512), .A2(n518), .ZN(n461) );
  XOR2_X1 U574 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n466) );
  XNOR2_X1 U575 ( .A(n466), .B(n465), .ZN(n467) );
  XOR2_X1 U576 ( .A(n468), .B(n467), .Z(n469) );
  NOR2_X1 U577 ( .A1(G902), .A2(n599), .ZN(n473) );
  XNOR2_X1 U578 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n471) );
  XOR2_X1 U579 ( .A(KEYINPUT104), .B(KEYINPUT9), .Z(n475) );
  XNOR2_X1 U580 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n474) );
  XNOR2_X1 U581 ( .A(n475), .B(n474), .ZN(n479) );
  XOR2_X1 U582 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n477) );
  XNOR2_X1 U583 ( .A(G134), .B(G122), .ZN(n476) );
  XNOR2_X1 U584 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U585 ( .A(n479), .B(n478), .Z(n483) );
  XNOR2_X1 U586 ( .A(n480), .B(n481), .ZN(n482) );
  XNOR2_X1 U587 ( .A(n483), .B(n482), .ZN(n486) );
  NAND2_X1 U588 ( .A1(n484), .A2(G217), .ZN(n485) );
  XOR2_X1 U589 ( .A(n486), .B(n485), .Z(n605) );
  NOR2_X1 U590 ( .A1(G902), .A2(n605), .ZN(n488) );
  XNOR2_X1 U591 ( .A(KEYINPUT106), .B(G478), .ZN(n487) );
  XNOR2_X1 U592 ( .A(n488), .B(n487), .ZN(n509) );
  NOR2_X1 U593 ( .A1(n506), .A2(n509), .ZN(n489) );
  XOR2_X1 U594 ( .A(n489), .B(KEYINPUT110), .Z(n555) );
  XNOR2_X1 U595 ( .A(n555), .B(KEYINPUT77), .ZN(n490) );
  NAND2_X1 U596 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X2 U597 ( .A(n492), .B(KEYINPUT35), .ZN(n724) );
  NOR2_X2 U598 ( .A1(n724), .A2(KEYINPUT44), .ZN(n493) );
  XNOR2_X1 U599 ( .A(n493), .B(KEYINPUT66), .ZN(n505) );
  NAND2_X1 U600 ( .A1(n509), .A2(n506), .ZN(n579) );
  INV_X1 U601 ( .A(n579), .ZN(n646) );
  AND2_X1 U602 ( .A1(n646), .A2(n655), .ZN(n494) );
  XNOR2_X1 U603 ( .A(KEYINPUT79), .B(n518), .ZN(n499) );
  NOR2_X1 U604 ( .A1(n654), .A2(n651), .ZN(n498) );
  AND2_X1 U605 ( .A1(n499), .A2(n498), .ZN(n501) );
  INV_X1 U606 ( .A(KEYINPUT78), .ZN(n500) );
  NAND2_X1 U607 ( .A1(n505), .A2(n528), .ZN(n524) );
  INV_X1 U608 ( .A(n506), .ZN(n508) );
  NAND2_X1 U609 ( .A1(n509), .A2(n508), .ZN(n563) );
  INV_X1 U610 ( .A(n563), .ZN(n630) );
  OR2_X1 U611 ( .A1(n593), .A2(n630), .ZN(n510) );
  XNOR2_X1 U612 ( .A(n510), .B(KEYINPUT108), .ZN(n549) );
  INV_X1 U613 ( .A(n549), .ZN(n643) );
  OR2_X1 U614 ( .A1(n545), .A2(n650), .ZN(n576) );
  NAND2_X1 U615 ( .A1(n514), .A2(n657), .ZN(n511) );
  NOR2_X1 U616 ( .A1(n576), .A2(n511), .ZN(n619) );
  INV_X1 U617 ( .A(n512), .ZN(n513) );
  NOR2_X1 U618 ( .A1(n657), .A2(n513), .ZN(n663) );
  NAND2_X1 U619 ( .A1(n663), .A2(n514), .ZN(n515) );
  XNOR2_X1 U620 ( .A(n515), .B(KEYINPUT100), .ZN(n516) );
  XNOR2_X1 U621 ( .A(KEYINPUT31), .B(n516), .ZN(n633) );
  NOR2_X1 U622 ( .A1(n619), .A2(n633), .ZN(n517) );
  NOR2_X1 U623 ( .A1(n643), .A2(n517), .ZN(n522) );
  INV_X1 U624 ( .A(n518), .ZN(n562) );
  AND2_X1 U625 ( .A1(n654), .A2(n562), .ZN(n519) );
  NAND2_X1 U626 ( .A1(n520), .A2(n519), .ZN(n616) );
  INV_X1 U627 ( .A(n616), .ZN(n521) );
  NOR2_X1 U628 ( .A1(n522), .A2(n521), .ZN(n523) );
  INV_X1 U629 ( .A(KEYINPUT84), .ZN(n530) );
  NAND2_X1 U630 ( .A1(n724), .A2(KEYINPUT44), .ZN(n525) );
  NAND2_X1 U631 ( .A1(n530), .A2(n525), .ZN(n527) );
  NAND2_X1 U632 ( .A1(n724), .A2(KEYINPUT84), .ZN(n526) );
  NAND2_X1 U633 ( .A1(n529), .A2(n528), .ZN(n532) );
  OR2_X1 U634 ( .A1(n530), .A2(KEYINPUT44), .ZN(n531) );
  NAND2_X2 U635 ( .A1(n534), .A2(n533), .ZN(n536) );
  INV_X1 U636 ( .A(KEYINPUT45), .ZN(n535) );
  XNOR2_X2 U637 ( .A(n536), .B(n535), .ZN(n705) );
  XOR2_X1 U638 ( .A(KEYINPUT47), .B(KEYINPUT67), .Z(n537) );
  NOR2_X1 U639 ( .A1(n643), .A2(n537), .ZN(n547) );
  OR2_X1 U640 ( .A1(n714), .A2(n538), .ZN(n539) );
  NOR2_X1 U641 ( .A1(G900), .A2(n539), .ZN(n541) );
  NOR2_X1 U642 ( .A1(n541), .A2(n540), .ZN(n574) );
  NOR2_X1 U643 ( .A1(n574), .A2(n654), .ZN(n542) );
  NAND2_X1 U644 ( .A1(n542), .A2(n655), .ZN(n561) );
  NOR2_X1 U645 ( .A1(n657), .A2(n561), .ZN(n543) );
  XOR2_X1 U646 ( .A(KEYINPUT28), .B(n543), .Z(n544) );
  NOR2_X1 U647 ( .A1(n545), .A2(n544), .ZN(n581) );
  NAND2_X1 U648 ( .A1(n581), .A2(n546), .ZN(n558) );
  INV_X1 U649 ( .A(n558), .ZN(n628) );
  NAND2_X1 U650 ( .A1(n547), .A2(n628), .ZN(n548) );
  XNOR2_X1 U651 ( .A(n548), .B(KEYINPUT70), .ZN(n553) );
  NAND2_X1 U652 ( .A1(n558), .A2(KEYINPUT82), .ZN(n550) );
  NAND2_X1 U653 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U654 ( .A1(n551), .A2(KEYINPUT47), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n553), .A2(n552), .ZN(n573) );
  NOR2_X1 U656 ( .A1(n574), .A2(n576), .ZN(n554) );
  NAND2_X1 U657 ( .A1(n554), .A2(n575), .ZN(n556) );
  OR2_X1 U658 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U659 ( .A1(n586), .A2(n557), .ZN(n627) );
  AND2_X1 U660 ( .A1(KEYINPUT47), .A2(n558), .ZN(n559) );
  NOR2_X1 U661 ( .A1(KEYINPUT82), .A2(n559), .ZN(n560) );
  NOR2_X1 U662 ( .A1(n627), .A2(n560), .ZN(n571) );
  INV_X1 U663 ( .A(n561), .ZN(n565) );
  NOR2_X1 U664 ( .A1(n563), .A2(n562), .ZN(n564) );
  NAND2_X1 U665 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U666 ( .A(n566), .B(KEYINPUT111), .ZN(n568) );
  NAND2_X1 U667 ( .A1(n568), .A2(n567), .ZN(n587) );
  NOR2_X1 U668 ( .A1(n586), .A2(n587), .ZN(n569) );
  XNOR2_X1 U669 ( .A(n569), .B(KEYINPUT36), .ZN(n570) );
  NAND2_X1 U670 ( .A1(n570), .A2(n589), .ZN(n636) );
  NAND2_X1 U671 ( .A1(n571), .A2(n636), .ZN(n572) );
  XOR2_X1 U672 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n582) );
  NAND2_X1 U673 ( .A1(n584), .A2(n583), .ZN(n585) );
  INV_X1 U674 ( .A(n586), .ZN(n592) );
  XNOR2_X1 U675 ( .A(KEYINPUT112), .B(n587), .ZN(n588) );
  NOR2_X1 U676 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U677 ( .A(n590), .B(KEYINPUT43), .ZN(n591) );
  NOR2_X1 U678 ( .A1(n592), .A2(n591), .ZN(n638) );
  NAND2_X1 U679 ( .A1(n594), .A2(n593), .ZN(n637) );
  INV_X1 U680 ( .A(n637), .ZN(n595) );
  NOR2_X2 U681 ( .A1(n705), .A2(n713), .ZN(n671) );
  XNOR2_X1 U682 ( .A(n671), .B(KEYINPUT2), .ZN(n597) );
  XOR2_X1 U683 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n598) );
  XNOR2_X1 U684 ( .A(n601), .B(n600), .ZN(n602) );
  NOR2_X1 U685 ( .A1(n602), .A2(n698), .ZN(n604) );
  XOR2_X1 U686 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n603) );
  XNOR2_X1 U687 ( .A(n604), .B(n603), .ZN(G60) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT123), .ZN(G63) );
  XNOR2_X1 U689 ( .A(n612), .B(n611), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n615), .B(n614), .ZN(G57) );
  XNOR2_X1 U691 ( .A(G101), .B(n616), .ZN(G3) );
  XOR2_X1 U692 ( .A(G104), .B(KEYINPUT113), .Z(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n630), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n618), .B(n617), .ZN(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n621) );
  NAND2_X1 U696 ( .A1(n619), .A2(n632), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n621), .B(n620), .ZN(n622) );
  XNOR2_X1 U698 ( .A(G107), .B(n622), .ZN(G9) );
  XOR2_X1 U699 ( .A(G110), .B(n623), .Z(n624) );
  XNOR2_X1 U700 ( .A(KEYINPUT114), .B(n624), .ZN(G12) );
  XOR2_X1 U701 ( .A(G128), .B(KEYINPUT29), .Z(n626) );
  NAND2_X1 U702 ( .A1(n632), .A2(n628), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n626), .B(n625), .ZN(G30) );
  XOR2_X1 U704 ( .A(G143), .B(n627), .Z(G45) );
  NAND2_X1 U705 ( .A1(n628), .A2(n630), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(G146), .ZN(G48) );
  NAND2_X1 U707 ( .A1(n630), .A2(n633), .ZN(n631) );
  XNOR2_X1 U708 ( .A(G113), .B(n631), .ZN(G15) );
  NAND2_X1 U709 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n634), .B(G116), .ZN(G18) );
  XOR2_X1 U711 ( .A(G125), .B(KEYINPUT37), .Z(n635) );
  XNOR2_X1 U712 ( .A(n636), .B(n635), .ZN(G27) );
  XNOR2_X1 U713 ( .A(G134), .B(n637), .ZN(G36) );
  XOR2_X1 U714 ( .A(G140), .B(n638), .Z(G42) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n675), .A2(n642), .ZN(n648) );
  NOR2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U718 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U719 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U720 ( .A(KEYINPUT117), .B(n649), .ZN(n667) );
  XOR2_X1 U721 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n653) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U723 ( .A(n653), .B(n652), .ZN(n661) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U725 ( .A(n656), .B(KEYINPUT49), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT115), .B(n659), .Z(n660) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n664), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n665), .A2(n676), .ZN(n666) );
  NAND2_X1 U732 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U733 ( .A(KEYINPUT52), .B(n668), .Z(n669) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n674) );
  NOR2_X1 U735 ( .A1(n671), .A2(KEYINPUT81), .ZN(n672) );
  XNOR2_X1 U736 ( .A(KEYINPUT2), .B(n672), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n678) );
  NAND2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n679), .A2(G953), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n680), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U742 ( .A(KEYINPUT85), .B(KEYINPUT80), .Z(n682) );
  XNOR2_X1 U743 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n681) );
  XNOR2_X1 U744 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U745 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U746 ( .A1(n686), .A2(n698), .ZN(n687) );
  XNOR2_X1 U747 ( .A(n687), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U748 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n690) );
  XNOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n689) );
  NOR2_X1 U750 ( .A1(n698), .A2(n693), .ZN(G54) );
  XNOR2_X1 U751 ( .A(n694), .B(KEYINPUT124), .ZN(n696) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U753 ( .A1(n698), .A2(n697), .ZN(G66) );
  XOR2_X1 U754 ( .A(G101), .B(n699), .Z(n700) );
  NAND2_X1 U755 ( .A1(n701), .A2(n700), .ZN(n709) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n702) );
  XOR2_X1 U757 ( .A(KEYINPUT61), .B(n702), .Z(n703) );
  NOR2_X1 U758 ( .A1(n704), .A2(n703), .ZN(n707) );
  NOR2_X1 U759 ( .A1(G953), .A2(n705), .ZN(n706) );
  NOR2_X1 U760 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U761 ( .A(n709), .B(n708), .ZN(G69) );
  XOR2_X1 U762 ( .A(n712), .B(n711), .Z(n716) );
  XNOR2_X1 U763 ( .A(n713), .B(n716), .ZN(n715) );
  NAND2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n721) );
  XNOR2_X1 U765 ( .A(G227), .B(n716), .ZN(n717) );
  NAND2_X1 U766 ( .A1(n717), .A2(G900), .ZN(n718) );
  XOR2_X1 U767 ( .A(KEYINPUT125), .B(n718), .Z(n719) );
  NAND2_X1 U768 ( .A1(G953), .A2(n719), .ZN(n720) );
  NAND2_X1 U769 ( .A1(n721), .A2(n720), .ZN(G72) );
  XNOR2_X1 U770 ( .A(n722), .B(G137), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(KEYINPUT126), .ZN(G39) );
  XOR2_X1 U772 ( .A(n724), .B(G122), .Z(G24) );
  XOR2_X1 U773 ( .A(n725), .B(G119), .Z(G21) );
  XNOR2_X1 U774 ( .A(G131), .B(n726), .ZN(G33) );
endmodule

