//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  NAND2_X1  g0012(.A1(G87), .A2(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G116), .B2(G270), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G58), .A2(G232), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G107), .A2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G50), .A2(G226), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G68), .ZN(new_n224));
  INV_X1    g0024(.A(G238), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT1), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT64), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n231), .A2(G1), .A3(G13), .ZN(new_n232));
  AND2_X1   g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n207), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n212), .B(new_n228), .C1(new_n234), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT65), .ZN(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NAND2_X1  g0053(.A1(new_n203), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n207), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G58), .ZN(new_n259));
  XOR2_X1   g0059(.A(new_n259), .B(KEYINPUT8), .Z(new_n260));
  NAND2_X1  g0060(.A1(new_n207), .A2(G33), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n254), .B1(new_n255), .B2(new_n257), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n230), .A2(new_n232), .A3(new_n263), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n202), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n206), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n264), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n269), .B(new_n272), .C1(new_n202), .C2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT66), .B1(new_n233), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n230), .A2(new_n232), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT66), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n256), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(G222), .A2(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n289), .A2(G223), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n283), .B(new_n291), .C1(G77), .C2(new_n287), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n293));
  INV_X1    g0093(.A(G274), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G226), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n293), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n292), .B(new_n296), .C1(new_n297), .C2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n276), .B(new_n301), .C1(new_n302), .C2(new_n300), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT10), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n300), .A2(new_n305), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n306), .B(new_n275), .C1(G179), .C2(new_n300), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G232), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G1698), .ZN(new_n310));
  AND2_X1   g0110(.A1(KEYINPUT3), .A2(G33), .ZN(new_n311));
  NOR2_X1   g0111(.A1(KEYINPUT3), .A2(G33), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n310), .B1(G226), .B2(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G33), .A2(G97), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n316));
  AOI211_X1 g0116(.A(KEYINPUT66), .B(new_n277), .C1(new_n230), .C2(new_n232), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n299), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G238), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n318), .A2(new_n320), .A3(new_n296), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n318), .A2(new_n323), .A3(new_n320), .A4(new_n296), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(G169), .A3(new_n326), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n322), .A2(G179), .A3(new_n324), .ZN(new_n328));
  AND2_X1   g0128(.A1(KEYINPUT70), .A2(KEYINPUT14), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n305), .B(new_n329), .C1(new_n322), .C2(new_n324), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n327), .B(new_n328), .C1(new_n330), .C2(new_n326), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n224), .A2(G20), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n332), .B1(new_n261), .B2(new_n214), .C1(new_n202), .C2(new_n257), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n268), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT11), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n274), .A2(new_n224), .ZN(new_n336));
  INV_X1    g0136(.A(G13), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G1), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n332), .ZN(new_n340));
  XOR2_X1   g0140(.A(new_n340), .B(KEYINPUT12), .Z(new_n341));
  AND2_X1   g0141(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n335), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n331), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n287), .A2(G238), .A3(G1698), .ZN(new_n346));
  AND2_X1   g0146(.A1(KEYINPUT69), .A2(G107), .ZN(new_n347));
  NOR2_X1   g0147(.A1(KEYINPUT69), .A2(G107), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n287), .A2(new_n289), .ZN(new_n351));
  OAI221_X1 g0151(.A(new_n346), .B1(new_n350), .B2(new_n287), .C1(new_n309), .C2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n295), .B1(new_n352), .B2(new_n283), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n215), .B2(new_n299), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n305), .ZN(new_n355));
  XOR2_X1   g0155(.A(KEYINPUT15), .B(G87), .Z(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n261), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT8), .B(G58), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n359), .A2(new_n257), .B1(new_n207), .B2(new_n214), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n268), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n271), .A2(new_n214), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(new_n214), .C2(new_n274), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n355), .B(new_n363), .C1(G179), .C2(new_n354), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n345), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n285), .A2(new_n207), .A3(new_n286), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n286), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n224), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n201), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n207), .A2(new_n256), .A3(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n366), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT72), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n311), .A2(new_n312), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n378), .B2(new_n207), .ZN(new_n379));
  INV_X1    g0179(.A(new_n370), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT71), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n373), .B2(new_n374), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n373), .A2(new_n382), .A3(new_n374), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n381), .A2(KEYINPUT16), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT72), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n387), .B(new_n366), .C1(new_n371), .C2(new_n375), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n377), .A2(new_n268), .A3(new_n386), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G87), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n256), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(G223), .A2(G1698), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n392), .B1(new_n285), .B2(new_n286), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n297), .A2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n395), .B1(new_n278), .B2(new_n282), .ZN(new_n396));
  OAI22_X1  g0196(.A1(new_n299), .A2(new_n309), .B1(new_n294), .B2(new_n293), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI221_X1 g0198(.A(new_n394), .B1(G223), .B2(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n399));
  INV_X1    g0199(.A(new_n391), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n316), .B2(new_n317), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n397), .A2(KEYINPUT73), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT73), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n296), .B(new_n404), .C1(new_n309), .C2(new_n299), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  OAI22_X1  g0206(.A1(new_n398), .A2(G200), .B1(new_n406), .B2(G190), .ZN(new_n407));
  INV_X1    g0207(.A(new_n260), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n274), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n260), .A2(new_n270), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n389), .A2(new_n407), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT17), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n389), .A2(new_n407), .A3(KEYINPUT17), .A4(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  INV_X1    g0216(.A(G179), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n402), .A2(new_n417), .A3(new_n403), .A4(new_n405), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n398), .B2(G169), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n416), .B(new_n419), .C1(new_n389), .C2(new_n411), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n389), .A2(new_n411), .ZN(new_n421));
  INV_X1    g0221(.A(new_n397), .ZN(new_n422));
  AOI21_X1  g0222(.A(G169), .B1(new_n402), .B2(new_n422), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n423), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT18), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n414), .B(new_n415), .C1(new_n420), .C2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n363), .B1(new_n354), .B2(G200), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n302), .B2(new_n354), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n325), .A2(G200), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n322), .A2(G190), .A3(new_n324), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n342), .A3(new_n335), .A4(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n428), .A2(new_n430), .A3(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n308), .A2(new_n365), .A3(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n390), .B(new_n216), .C1(new_n347), .C2(new_n348), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n314), .A2(new_n207), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n436), .A2(KEYINPUT19), .A3(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n287), .A2(new_n207), .A3(G68), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT19), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n261), .B2(new_n216), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n438), .A2(KEYINPUT81), .A3(new_n439), .A4(new_n441), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n268), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n206), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n264), .A2(new_n267), .A3(new_n270), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n356), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n357), .A2(new_n271), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n446), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n225), .A2(new_n289), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n215), .A2(G1698), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n453), .B(new_n454), .C1(new_n311), .C2(new_n312), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n455), .B1(new_n256), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(new_n316), .B2(new_n317), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n206), .A2(G45), .A3(G274), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n298), .B(G250), .C1(G1), .C2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n305), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n452), .A2(new_n463), .ZN(new_n464));
  OR2_X1    g0264(.A1(new_n462), .A2(G179), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n462), .A2(new_n302), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n466), .B1(G200), .B2(new_n462), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n449), .A2(G87), .ZN(new_n468));
  AND3_X1   g0268(.A1(new_n446), .A2(new_n468), .A3(new_n451), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n464), .A2(new_n465), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT79), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n471), .B1(new_n472), .B2(G41), .ZN(new_n473));
  INV_X1    g0273(.A(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n206), .B(G45), .C1(new_n474), .C2(KEYINPUT5), .ZN(new_n477));
  OAI211_X1 g0277(.A(G257), .B(new_n298), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n477), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n475), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(G274), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n482), .B(KEYINPUT80), .ZN(new_n483));
  OAI211_X1 g0283(.A(G250), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT77), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT77), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n287), .A2(new_n486), .A3(G250), .A4(G1698), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n351), .B2(new_n215), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .A4(new_n289), .ZN(new_n491));
  AND3_X1   g0291(.A1(KEYINPUT76), .A2(G33), .A3(G283), .ZN(new_n492));
  AOI21_X1  g0292(.A(KEYINPUT76), .B1(G33), .B2(G283), .ZN(new_n493));
  OR2_X1    g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n488), .A2(new_n490), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n283), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT78), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT78), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n495), .A2(new_n498), .A3(new_n283), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n483), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G200), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n270), .A2(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n448), .A2(new_n216), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT74), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT74), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n505), .B(new_n507), .C1(new_n216), .C2(G107), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n505), .A2(new_n507), .ZN(new_n509));
  XNOR2_X1  g0309(.A(G97), .B(G107), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n511), .A2(new_n207), .B1(new_n214), .B2(new_n257), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n369), .A2(new_n370), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n349), .ZN(new_n516));
  OAI221_X1 g0316(.A(KEYINPUT75), .B1(new_n214), .B2(new_n257), .C1(new_n511), .C2(new_n207), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(new_n502), .B(new_n503), .C1(new_n518), .C2(new_n268), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n482), .B1(new_n495), .B2(new_n283), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(G190), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n501), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n287), .A2(new_n207), .A3(G87), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n256), .A2(new_n456), .A3(G20), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT23), .B(G20), .C1(new_n347), .C2(new_n348), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n207), .B2(G107), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  XOR2_X1   g0330(.A(KEYINPUT85), .B(KEYINPUT22), .Z(new_n531));
  NAND4_X1  g0331(.A1(new_n531), .A2(new_n207), .A3(G87), .A4(new_n287), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n525), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(KEYINPUT86), .A2(KEYINPUT24), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n534), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n525), .A2(new_n530), .A3(new_n532), .A4(new_n536), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n535), .A2(new_n537), .B1(KEYINPUT86), .B2(KEYINPUT24), .ZN(new_n538));
  INV_X1    g0338(.A(new_n268), .ZN(new_n539));
  OR2_X1    g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n289), .C1(new_n311), .C2(new_n312), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n316), .B2(new_n317), .ZN(new_n545));
  OAI211_X1 g0345(.A(G264), .B(new_n298), .C1(new_n476), .C2(new_n477), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n481), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G190), .ZN(new_n549));
  INV_X1    g0349(.A(G107), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n338), .A2(G20), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n551), .B(KEYINPUT25), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n449), .B2(G107), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(G200), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n540), .A2(new_n549), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n502), .B1(new_n518), .B2(new_n268), .ZN(new_n556));
  INV_X1    g0356(.A(new_n503), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n483), .A2(new_n497), .A3(new_n417), .A4(new_n499), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n520), .A2(G169), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AND4_X1   g0361(.A1(new_n470), .A2(new_n522), .A3(new_n555), .A4(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT82), .B1(new_n351), .B2(new_n217), .ZN(new_n563));
  OAI211_X1 g0363(.A(G264), .B(G1698), .C1(new_n311), .C2(new_n312), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT83), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n564), .A2(new_n565), .B1(new_n378), .B2(G303), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n287), .A2(KEYINPUT83), .A3(G264), .A4(G1698), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT82), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n287), .A2(new_n568), .A3(G257), .A4(new_n289), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n563), .A2(new_n566), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n283), .ZN(new_n571));
  OAI211_X1 g0371(.A(G270), .B(new_n298), .C1(new_n476), .C2(new_n477), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n481), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G20), .B1(new_n256), .B2(G97), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n492), .B2(new_n493), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n456), .A2(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n577), .A2(new_n265), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT20), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n577), .A2(new_n265), .A3(KEYINPUT20), .A4(new_n578), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n339), .A2(new_n578), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n583), .B(new_n585), .C1(new_n456), .C2(new_n448), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n575), .A2(new_n586), .A3(G169), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT21), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT84), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n573), .B1(new_n570), .B2(new_n283), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n592), .A2(new_n588), .A3(new_n305), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n572), .A2(G179), .A3(new_n481), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n283), .B2(new_n570), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n586), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n587), .A2(KEYINPUT84), .A3(new_n588), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n591), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n553), .B1(new_n538), .B2(new_n539), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(KEYINPUT87), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT87), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n601), .B(new_n553), .C1(new_n538), .C2(new_n539), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n547), .A2(G169), .ZN(new_n603));
  XNOR2_X1  g0403(.A(new_n603), .B(KEYINPUT88), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n548), .A2(G179), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n600), .A2(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n598), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n586), .B1(new_n575), .B2(G200), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n302), .B2(new_n575), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n435), .A2(new_n562), .A3(new_n607), .A4(new_n609), .ZN(G372));
  AND2_X1   g0410(.A1(new_n414), .A2(new_n415), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n365), .A2(new_n611), .A3(new_n433), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT89), .ZN(new_n613));
  OR3_X1    g0413(.A1(new_n420), .A2(new_n426), .A3(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n420), .B2(new_n426), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n304), .B1(new_n612), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n307), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n604), .A2(new_n605), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n599), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n562), .B1(new_n598), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n464), .A2(new_n465), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n467), .A2(new_n469), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(new_n561), .ZN(new_n627));
  INV_X1    g0427(.A(new_n561), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n470), .A3(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n622), .A2(new_n623), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n435), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n619), .A2(new_n632), .ZN(G369));
  NAND2_X1  g0433(.A1(new_n338), .A2(new_n207), .ZN(new_n634));
  OR3_X1    g0434(.A1(new_n634), .A2(KEYINPUT90), .A3(KEYINPUT27), .ZN(new_n635));
  INV_X1    g0435(.A(G213), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n634), .B2(KEYINPUT27), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT90), .B1(new_n634), .B2(KEYINPUT27), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n635), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(G343), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n586), .A2(new_n641), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n598), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n598), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n609), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g0446(.A(KEYINPUT91), .B(G330), .Z(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n555), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n606), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n600), .A2(new_n602), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n641), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n650), .A2(new_n652), .B1(new_n606), .B2(new_n641), .ZN(new_n653));
  INV_X1    g0453(.A(new_n641), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n598), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n641), .B(KEYINPUT92), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n655), .A2(new_n650), .B1(new_n621), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(G399));
  INV_X1    g0462(.A(new_n210), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G41), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(G1), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n436), .A2(G116), .ZN(new_n667));
  OAI22_X1  g0467(.A1(new_n666), .A2(new_n667), .B1(new_n235), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n631), .A2(new_n660), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(KEYINPUT29), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n630), .A2(new_n623), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT93), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n562), .B1(new_n606), .B2(new_n598), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n630), .A2(KEYINPUT93), .A3(new_n623), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n654), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n671), .B1(new_n678), .B2(KEYINPUT29), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n562), .A2(new_n607), .A3(new_n609), .A4(new_n660), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n545), .A2(new_n546), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n462), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(new_n520), .A3(new_n595), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT30), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n682), .A2(new_n595), .A3(new_n520), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n547), .A2(new_n462), .A3(new_n417), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n592), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n500), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n684), .A2(new_n686), .B1(new_n500), .B2(new_n689), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n654), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n680), .B(new_n692), .C1(KEYINPUT31), .C2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n647), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n679), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n669), .B1(new_n698), .B2(G1), .ZN(G364));
  OR2_X1    g0499(.A1(new_n646), .A2(new_n647), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n337), .A2(G20), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n666), .B1(G45), .B2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n648), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n207), .A2(G190), .ZN(new_n705));
  NOR2_X1   g0505(.A1(G179), .A2(G200), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT95), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n207), .A2(new_n302), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(new_n417), .A3(G200), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n711), .A2(G329), .B1(G303), .B2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(G294), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n207), .B1(new_n706), .B2(G190), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n715), .B(new_n378), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n417), .A2(G200), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n721), .A2(G322), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n705), .A2(new_n417), .A3(G200), .ZN(new_n723));
  INV_X1    g0523(.A(G283), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G190), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OR2_X1    g0528(.A1(KEYINPUT33), .A2(G317), .ZN(new_n729));
  NAND2_X1  g0529(.A1(KEYINPUT33), .A2(G317), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NOR4_X1   g0531(.A1(new_n718), .A2(new_n722), .A3(new_n725), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n705), .A2(new_n719), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G311), .ZN(new_n735));
  INV_X1    g0535(.A(G326), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n726), .A2(new_n302), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n732), .B(new_n735), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT97), .Z(new_n740));
  XNOR2_X1  g0540(.A(new_n717), .B(KEYINPUT96), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI22_X1  g0542(.A1(new_n742), .A2(G97), .B1(G50), .B2(new_n737), .ZN(new_n743));
  INV_X1    g0543(.A(G58), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n743), .B1(new_n744), .B2(new_n720), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n713), .A2(new_n390), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n287), .B1(new_n723), .B2(new_n550), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n748), .B1(new_n224), .B2(new_n728), .C1(new_n214), .C2(new_n733), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n711), .A2(G159), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT32), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n740), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n233), .B1(G20), .B2(new_n305), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n210), .A2(G355), .A3(new_n287), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n252), .A2(G45), .ZN(new_n759));
  XOR2_X1   g0559(.A(new_n759), .B(KEYINPUT94), .Z(new_n760));
  NOR2_X1   g0560(.A1(new_n663), .A2(new_n287), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G45), .B2(new_n235), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n758), .B1(G116), .B2(new_n210), .C1(new_n760), .C2(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n752), .A2(new_n753), .B1(new_n757), .B2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n756), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n646), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n704), .B1(new_n766), .B2(new_n703), .ZN(G396));
  NOR2_X1   g0567(.A1(new_n364), .A2(new_n641), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n363), .A2(new_n641), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n430), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n770), .B2(new_n364), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n670), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n631), .A2(new_n660), .A3(new_n771), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(new_n696), .Z(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n703), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n772), .A2(new_n754), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n711), .A2(G311), .B1(G97), .B2(new_n742), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n727), .A2(G283), .ZN(new_n780));
  INV_X1    g0580(.A(new_n723), .ZN(new_n781));
  AOI22_X1  g0581(.A1(G107), .A2(new_n714), .B1(new_n781), .B2(G87), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n720), .A2(new_n716), .B1(new_n733), .B2(new_n456), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n287), .B(new_n783), .C1(G303), .C2(new_n737), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n723), .A2(new_n224), .ZN(new_n786));
  INV_X1    g0586(.A(G132), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n287), .B1(new_n710), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(KEYINPUT34), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n727), .A2(G150), .B1(new_n737), .B2(G137), .ZN(new_n790));
  INV_X1    g0590(.A(G143), .ZN(new_n791));
  INV_X1    g0591(.A(G159), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(new_n791), .B2(new_n720), .C1(new_n792), .C2(new_n733), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n786), .B(new_n788), .C1(new_n789), .C2(new_n793), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n794), .B1(new_n789), .B2(new_n793), .C1(new_n202), .C2(new_n713), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n717), .A2(new_n744), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n785), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(new_n753), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n753), .A2(new_n754), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n214), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n778), .A2(new_n702), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n777), .A2(new_n801), .ZN(G384));
  INV_X1    g0602(.A(KEYINPUT104), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n691), .A2(new_n803), .A3(new_n641), .ZN(new_n804));
  OAI21_X1  g0604(.A(KEYINPUT104), .B1(new_n693), .B2(new_n654), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT31), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT105), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n694), .A2(KEYINPUT31), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n804), .A2(new_n805), .A3(KEYINPUT105), .A4(new_n806), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n809), .A2(new_n680), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g0612(.A1(new_n331), .A2(new_n343), .A3(new_n654), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n343), .A2(new_n641), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n331), .A2(new_n343), .B1(new_n433), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT99), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT99), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n331), .A2(new_n343), .A3(new_n654), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n433), .A2(new_n814), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n817), .B(new_n818), .C1(new_n344), .C2(new_n819), .ZN(new_n820));
  AND3_X1   g0620(.A1(new_n816), .A2(new_n820), .A3(new_n771), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n812), .A2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n639), .B(KEYINPUT102), .Z(new_n825));
  NAND2_X1  g0625(.A1(new_n421), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(new_n616), .B2(new_n611), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n421), .A2(new_n425), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n828), .A2(new_n826), .A3(new_n412), .ZN(new_n829));
  XOR2_X1   g0629(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n830));
  XNOR2_X1  g0630(.A(new_n829), .B(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n824), .B1(new_n827), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n828), .A2(new_n826), .A3(new_n412), .A4(new_n830), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n386), .A2(new_n268), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n383), .B1(new_n515), .B2(G68), .ZN(new_n835));
  AOI21_X1  g0635(.A(KEYINPUT16), .B1(new_n835), .B2(new_n385), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n411), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n425), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n412), .A2(new_n838), .A3(KEYINPUT101), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT101), .B1(new_n412), .B2(new_n838), .ZN(new_n840));
  INV_X1    g0640(.A(new_n639), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n833), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n427), .A2(KEYINPUT100), .A3(new_n842), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT100), .B1(new_n427), .B2(new_n842), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n845), .B(KEYINPUT38), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n832), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n823), .A2(new_n849), .A3(KEYINPUT40), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n824), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n822), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT106), .B1(new_n853), .B2(KEYINPUT40), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n427), .A2(new_n842), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT100), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n427), .A2(KEYINPUT100), .A3(new_n842), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n859), .B2(new_n845), .ZN(new_n860));
  INV_X1    g0660(.A(new_n848), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n812), .B(new_n821), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT106), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT40), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n850), .B1(new_n854), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT107), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n435), .A2(new_n812), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n867), .B(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n647), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT39), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n849), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n852), .A2(KEYINPUT39), .A3(new_n848), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n813), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n616), .A2(new_n825), .ZN(new_n877));
  INV_X1    g0677(.A(new_n768), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n774), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n816), .A2(new_n820), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n852), .A2(new_n848), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n876), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n435), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n679), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n619), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n884), .B(new_n887), .Z(new_n888));
  XNOR2_X1  g0688(.A(new_n870), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n206), .B2(new_n701), .ZN(new_n890));
  OAI21_X1  g0690(.A(G77), .B1(new_n744), .B2(new_n224), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n891), .A2(new_n235), .B1(G50), .B2(new_n224), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(G1), .A3(new_n337), .ZN(new_n893));
  INV_X1    g0693(.A(new_n511), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n456), .B1(new_n894), .B2(KEYINPUT35), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(new_n234), .C1(KEYINPUT35), .C2(new_n894), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT98), .B(KEYINPUT36), .Z(new_n897));
  XNOR2_X1  g0697(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n890), .A2(new_n893), .A3(new_n898), .ZN(G367));
  XNOR2_X1  g0699(.A(new_n664), .B(KEYINPUT41), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n522), .B(new_n561), .C1(new_n519), .C2(new_n660), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n628), .A2(new_n659), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n661), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT44), .Z(new_n905));
  NAND2_X1  g0705(.A1(new_n661), .A2(new_n903), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT45), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n658), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT110), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n655), .A2(new_n650), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n648), .A2(new_n657), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n658), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n697), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n900), .B1(new_n916), .B2(new_n697), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n206), .B1(new_n701), .B2(G45), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n903), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n920), .A2(new_n911), .A3(KEYINPUT42), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT109), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT42), .B1(new_n920), .B2(new_n911), .ZN(new_n923));
  INV_X1    g0723(.A(new_n606), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n561), .B1(new_n901), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT108), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n922), .B(new_n923), .C1(new_n659), .C2(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT43), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n623), .A2(new_n469), .A3(new_n654), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n470), .B1(new_n469), .B2(new_n654), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n927), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n931), .A2(KEYINPUT43), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n933), .B(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n658), .A2(new_n920), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n919), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n742), .A2(G68), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n939), .B1(new_n744), .B2(new_n713), .C1(new_n791), .C2(new_n738), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n723), .A2(new_n214), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n711), .A2(G137), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n287), .B1(new_n728), .B2(new_n792), .ZN(new_n943));
  NOR4_X1   g0743(.A1(new_n940), .A2(new_n941), .A3(new_n942), .A4(new_n943), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n202), .B2(new_n733), .C1(new_n255), .C2(new_n720), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n711), .A2(G317), .B1(G303), .B2(new_n721), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n724), .B2(new_n733), .C1(new_n350), .C2(new_n717), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT46), .B1(new_n714), .B2(G116), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n714), .A2(KEYINPUT46), .A3(G116), .ZN(new_n949));
  NOR3_X1   g0749(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n781), .A2(G97), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n727), .A2(G294), .B1(new_n737), .B2(G311), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n945), .B1(new_n953), .B2(new_n287), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n753), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n932), .A2(new_n756), .ZN(new_n957));
  INV_X1    g0757(.A(new_n761), .ZN(new_n958));
  OAI221_X1 g0758(.A(new_n757), .B1(new_n210), .B2(new_n357), .C1(new_n958), .C2(new_n244), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n956), .A2(new_n702), .A3(new_n957), .A4(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n938), .A2(new_n960), .ZN(G387));
  AOI21_X1  g0761(.A(new_n665), .B1(new_n697), .B2(new_n913), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n915), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n359), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n202), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT50), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n224), .A2(new_n214), .ZN(new_n967));
  NOR4_X1   g0767(.A1(new_n966), .A2(G45), .A3(new_n967), .A4(new_n667), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n761), .B1(new_n241), .B2(new_n460), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n667), .A2(new_n210), .A3(new_n287), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n210), .A2(G107), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n757), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n734), .A2(G303), .B1(G311), .B2(new_n727), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n721), .A2(G317), .ZN(new_n975));
  XOR2_X1   g0775(.A(KEYINPUT111), .B(G322), .Z(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n975), .C1(new_n738), .C2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT48), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n724), .B2(new_n717), .C1(new_n716), .C2(new_n713), .ZN(new_n979));
  XOR2_X1   g0779(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n287), .B1(new_n781), .B2(G116), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n981), .B(new_n982), .C1(new_n736), .C2(new_n710), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n287), .B1(new_n738), .B2(new_n792), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n951), .B1(new_n710), .B2(new_n255), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n741), .A2(new_n357), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n713), .A2(new_n214), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI211_X1 g0788(.A(new_n984), .B(new_n988), .C1(new_n408), .C2(new_n727), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n202), .B2(new_n720), .C1(new_n224), .C2(new_n733), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n753), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n702), .B(new_n973), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT113), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n994), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n653), .A2(new_n756), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n963), .B1(new_n918), .B2(new_n913), .C1(new_n995), .C2(new_n998), .ZN(G393));
  NOR2_X1   g0799(.A1(new_n908), .A2(new_n658), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n910), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n918), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n757), .B1(new_n216), .B2(new_n210), .C1(new_n249), .C2(new_n958), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(new_n702), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT114), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n378), .B1(new_n724), .B2(new_n713), .C1(new_n710), .C2(new_n976), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n721), .A2(G311), .B1(G317), .B2(new_n737), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n1008), .B(KEYINPUT52), .Z(new_n1009));
  NAND2_X1  g0809(.A1(new_n727), .A2(G303), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n717), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n781), .A2(G107), .B1(new_n1011), .B2(G116), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1007), .B(new_n1013), .C1(G294), .C2(new_n734), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n378), .B1(new_n727), .B2(G50), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G68), .A2(new_n714), .B1(new_n781), .B2(G87), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1015), .B(new_n1016), .C1(new_n710), .C2(new_n791), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n738), .A2(new_n255), .B1(new_n720), .B2(new_n792), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT51), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n214), .B2(new_n741), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1017), .B(new_n1020), .C1(new_n964), .C2(new_n734), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n753), .B1(new_n1014), .B2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1006), .B(new_n1022), .C1(new_n903), .C2(new_n765), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1003), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT115), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n916), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1026), .B(new_n664), .C1(new_n914), .C2(new_n1001), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(G390));
  AND2_X1   g0828(.A1(new_n677), .A2(new_n654), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n770), .A2(new_n364), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n768), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n818), .B(new_n849), .C1(new_n1031), .C2(new_n880), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n874), .B1(new_n881), .B2(new_n813), .ZN(new_n1033));
  NOR3_X1   g0833(.A1(new_n696), .A2(new_n772), .A3(new_n880), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1032), .A2(new_n1033), .B1(G330), .B2(new_n823), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n435), .A2(G330), .A3(new_n812), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n619), .B(new_n1038), .C1(new_n679), .C2(new_n885), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n812), .A2(G330), .A3(new_n771), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1034), .B1(new_n880), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n1031), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n880), .B1(new_n696), .B2(new_n772), .ZN(new_n1043));
  INV_X1    g0843(.A(G330), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1043), .B1(new_n1044), .B2(new_n822), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n879), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1039), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1037), .A2(new_n1049), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n1048), .B(KEYINPUT116), .Z(new_n1051));
  AOI211_X1 g0851(.A(new_n665), .B(new_n1050), .C1(new_n1037), .C2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n875), .A2(new_n755), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n350), .A2(new_n728), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n746), .B(new_n1054), .C1(new_n711), .C2(G294), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n734), .A2(G97), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n786), .B1(new_n742), .B2(G77), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n378), .B1(new_n720), .B2(new_n456), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G283), .B2(new_n737), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(G128), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n741), .A2(new_n792), .B1(new_n738), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G50), .B2(new_n781), .ZN(new_n1063));
  XOR2_X1   g0863(.A(KEYINPUT54), .B(G143), .Z(new_n1064));
  AOI22_X1  g0864(.A1(new_n734), .A2(new_n1064), .B1(G137), .B2(new_n727), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT117), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n287), .B1(new_n720), .B2(new_n787), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n711), .B2(G125), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n713), .A2(new_n255), .ZN(new_n1069));
  XOR2_X1   g0869(.A(KEYINPUT118), .B(KEYINPUT53), .Z(new_n1070));
  XNOR2_X1  g0870(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1063), .A2(new_n1066), .A3(new_n1068), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n992), .B1(new_n1060), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n799), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(new_n408), .ZN(new_n1075));
  OR3_X1    g0875(.A1(new_n1053), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n1037), .A2(new_n918), .B1(new_n703), .B2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1052), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G378));
  INV_X1    g0879(.A(new_n1039), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1037), .B2(new_n1049), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n275), .A2(new_n841), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT120), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n308), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n304), .A2(KEYINPUT120), .A3(new_n307), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  XOR2_X1   g0887(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1088));
  NAND3_X1  g0888(.A1(new_n1084), .A2(new_n1082), .A3(new_n1085), .ZN(new_n1089));
  AND3_X1   g0889(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1088), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT121), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n866), .B2(G330), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n823), .A2(new_n849), .A3(KEYINPUT40), .ZN(new_n1095));
  AOI211_X1 g0895(.A(KEYINPUT106), .B(KEYINPUT40), .C1(new_n823), .C2(new_n882), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n1097));
  OAI211_X1 g0897(.A(G330), .B(new_n1095), .C1(new_n1096), .C2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1098), .A2(KEYINPUT121), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1094), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n854), .A2(new_n865), .ZN(new_n1101));
  NAND4_X1  g0901(.A1(new_n1101), .A2(new_n1093), .A3(G330), .A4(new_n1095), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1092), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1100), .A2(new_n884), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n884), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1098), .A2(KEYINPUT121), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1103), .B1(new_n1107), .B2(new_n1102), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1044), .B(new_n850), .C1(new_n854), .C2(new_n865), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1092), .B1(new_n1109), .B2(new_n1093), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1106), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1081), .A2(new_n1105), .A3(new_n1111), .A4(KEYINPUT57), .ZN(new_n1112));
  AND2_X1   g0912(.A1(new_n1112), .A2(new_n664), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1081), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT122), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n884), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1108), .A2(new_n1110), .A3(new_n1106), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1105), .A2(new_n1111), .A3(KEYINPUT122), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1114), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1113), .B1(new_n1120), .B2(KEYINPUT57), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1103), .A2(new_n754), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n939), .B1(new_n456), .B2(new_n738), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n987), .B1(G58), .B2(new_n781), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n710), .B2(new_n724), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1125), .A2(G41), .A3(new_n287), .ZN(new_n1126));
  XOR2_X1   g0926(.A(new_n1126), .B(KEYINPUT119), .Z(new_n1127));
  AOI211_X1 g0927(.A(new_n1123), .B(new_n1127), .C1(new_n356), .C2(new_n734), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n216), .B2(new_n728), .C1(new_n550), .C2(new_n720), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(new_n1129), .B(KEYINPUT58), .ZN(new_n1130));
  AOI21_X1  g0930(.A(G50), .B1(new_n286), .B2(new_n474), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(G128), .A2(new_n721), .B1(new_n734), .B2(G137), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n714), .A2(new_n1064), .B1(G132), .B2(new_n727), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n737), .A2(G125), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n741), .A2(new_n255), .ZN(new_n1136));
  OR3_X1    g0936(.A1(new_n1135), .A2(KEYINPUT59), .A3(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(G41), .B1(new_n711), .B2(G124), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(new_n256), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G159), .B2(new_n781), .ZN(new_n1140));
  OAI21_X1  g0940(.A(KEYINPUT59), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1131), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1130), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n753), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n799), .A2(new_n202), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1122), .A2(new_n702), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n1002), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1121), .A2(new_n1149), .ZN(G375));
  NAND3_X1  g0950(.A1(new_n1042), .A2(new_n1039), .A3(new_n1047), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1051), .A2(new_n900), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n918), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n755), .B1(new_n816), .B2(new_n820), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n710), .A2(new_n1061), .B1(new_n792), .B2(new_n713), .ZN(new_n1155));
  XOR2_X1   g0955(.A(new_n1155), .B(KEYINPUT123), .Z(new_n1156));
  NAND2_X1  g0956(.A1(new_n1064), .A2(new_n727), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n738), .A2(new_n787), .B1(new_n733), .B2(new_n255), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n742), .B2(G50), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G137), .B2(new_n721), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1161), .B(new_n287), .C1(new_n744), .C2(new_n723), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n720), .A2(new_n724), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1163), .B(new_n986), .C1(G116), .C2(new_n727), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n737), .A2(G294), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n941), .B1(new_n711), .B2(G303), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n350), .A2(new_n733), .B1(new_n713), .B2(new_n216), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n1167), .A2(new_n287), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n992), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1074), .A2(G68), .ZN(new_n1171));
  NOR3_X1   g0971(.A1(new_n1154), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1153), .B1(new_n702), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1152), .A2(new_n1173), .ZN(G381));
  NOR2_X1   g0974(.A1(G390), .A2(G387), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(new_n1176), .A2(G396), .A3(G393), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1121), .A2(new_n1078), .A3(new_n1149), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1178), .A2(G384), .A3(G381), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(G407));
  OAI211_X1 g0980(.A(G407), .B(G213), .C1(G343), .C2(new_n1178), .ZN(G409));
  NAND2_X1  g0981(.A1(new_n1112), .A2(new_n664), .ZN(new_n1182));
  AND3_X1   g0982(.A1(new_n1105), .A2(new_n1111), .A3(KEYINPUT122), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT122), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1081), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT57), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1182), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1002), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1146), .ZN(new_n1189));
  OAI21_X1  g0989(.A(G378), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n636), .A2(G343), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1120), .A2(new_n900), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1105), .A2(new_n1111), .A3(new_n1002), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1193), .A2(new_n1078), .A3(new_n1146), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT60), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1151), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1197), .A2(new_n665), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1151), .A2(new_n1196), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(new_n1049), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n1173), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(G384), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1190), .A2(new_n1192), .A3(new_n1195), .A4(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT63), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1202), .A2(KEYINPUT124), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(KEYINPUT124), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1191), .A2(G2897), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1205), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1191), .B1(G375), .B2(G378), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1209), .B1(new_n1210), .B2(new_n1195), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT61), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g1013(.A(G393), .B(G396), .Z(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT125), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(G390), .A2(G387), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1216), .B1(new_n1218), .B2(new_n1175), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1176), .A2(new_n1217), .A3(new_n1215), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1204), .A2(new_n1213), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1190), .A2(new_n1192), .A3(new_n1195), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(KEYINPUT124), .B2(new_n1202), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1212), .A3(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1203), .A2(KEYINPUT62), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT62), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1210), .A2(new_n1228), .A3(new_n1195), .A4(new_n1202), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT61), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1226), .A2(new_n1227), .A3(new_n1229), .A4(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1221), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1222), .A2(new_n1233), .ZN(G405));
  INV_X1    g1034(.A(KEYINPUT127), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1221), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1219), .A2(new_n1220), .A3(KEYINPUT127), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1190), .A2(new_n1178), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT126), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1238), .A2(new_n1239), .A3(new_n1202), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1202), .B(KEYINPUT126), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n1190), .A3(new_n1178), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1236), .A2(new_n1237), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1242), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n1235), .A3(new_n1221), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(G402));
endmodule


