//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(new_n202), .A2(G50), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  INV_X1    g0020(.A(G257), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n204), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT64), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n222), .A2(new_n223), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n214), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n213), .B(new_n217), .C1(new_n229), .C2(KEYINPUT1), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  INV_X1    g0045(.A(G68), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G50), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G58), .B(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n243), .B(new_n250), .ZN(G351));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G1698), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n252), .A2(G222), .A3(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n252), .A2(G1698), .ZN(new_n256));
  INV_X1    g0056(.A(G223), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n254), .B1(new_n255), .B2(new_n252), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n260), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n261), .A2(new_n265), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(G226), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n262), .A2(KEYINPUT66), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT66), .B1(new_n262), .B2(new_n269), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n210), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G13), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n283));
  NOR3_X1   g0083(.A1(new_n279), .A2(new_n211), .A3(G1), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT68), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G1), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n283), .A2(new_n287), .B1(new_n288), .B2(G20), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G50), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT8), .B(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n211), .A2(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G150), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI22_X1  g0095(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n211), .B1(new_n201), .B2(new_n244), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n277), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT67), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n298), .A2(new_n299), .B1(new_n244), .B2(new_n284), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n290), .B(new_n300), .C1(new_n299), .C2(new_n298), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n275), .B(new_n301), .C1(G179), .C2(new_n273), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT69), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT9), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n301), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n301), .B2(new_n304), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(G190), .B1(new_n271), .B2(new_n272), .ZN(new_n308));
  INV_X1    g0108(.A(new_n272), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G200), .A3(new_n270), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n301), .A2(new_n304), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n308), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n313), .B1(new_n307), .B2(new_n312), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n302), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n252), .A2(G232), .A3(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n322), .A2(new_n324), .A3(G226), .A4(new_n253), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT70), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT70), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n252), .A2(new_n327), .A3(G226), .A4(new_n253), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n260), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n268), .A2(G238), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n266), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT13), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n267), .B1(G238), .B2(new_n268), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n318), .A2(new_n319), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n328), .B2(new_n326), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n334), .B(new_n335), .C1(new_n337), .C2(new_n260), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G169), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n333), .A2(new_n338), .A3(G179), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT14), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n343), .A3(G169), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n288), .A2(G20), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n285), .A2(G68), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT71), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n294), .A2(G50), .B1(G20), .B2(new_n246), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n255), .B2(new_n292), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n350), .A2(new_n277), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n284), .A2(new_n246), .ZN(new_n353));
  XNOR2_X1  g0153(.A(new_n353), .B(KEYINPUT12), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(KEYINPUT11), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n348), .A2(new_n352), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n345), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n356), .ZN(new_n358));
  INV_X1    g0158(.A(G190), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n339), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G200), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n333), .B2(new_n338), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n357), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n252), .A2(G232), .A3(new_n253), .ZN(new_n366));
  INV_X1    g0166(.A(G238), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n366), .B1(new_n205), .B2(new_n252), .C1(new_n256), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n261), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n267), .B1(G244), .B2(new_n268), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n274), .ZN(new_n372));
  INV_X1    g0172(.A(new_n291), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT15), .B(G87), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n374), .B1(new_n292), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(new_n277), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n285), .A2(G77), .A3(new_n346), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n377), .B(new_n378), .C1(G77), .C2(new_n281), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n372), .B(new_n379), .C1(G179), .C2(new_n371), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n371), .A2(G200), .ZN(new_n382));
  INV_X1    g0182(.A(new_n371), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n379), .B1(G190), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n381), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n322), .A2(new_n324), .A3(G226), .A4(G1698), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n322), .A2(new_n324), .A3(G223), .A4(new_n253), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G87), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n261), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n288), .B1(G41), .B2(G45), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n260), .A2(G232), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n266), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n361), .B1(new_n390), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n393), .B1(new_n261), .B2(new_n389), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(G190), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g0197(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n398));
  NAND2_X1  g0198(.A1(new_n294), .A2(G159), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT72), .ZN(new_n400));
  XNOR2_X1  g0200(.A(G58), .B(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(G20), .ZN(new_n402));
  AND2_X1   g0202(.A1(G58), .A2(G68), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n400), .B(G20), .C1(new_n403), .C2(new_n201), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n399), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT7), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n252), .B2(G20), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n323), .A2(G33), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n321), .A2(KEYINPUT3), .ZN(new_n410));
  OAI211_X1 g0210(.A(KEYINPUT7), .B(new_n211), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n246), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n398), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n322), .A2(new_n324), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n414), .B2(new_n211), .ZN(new_n415));
  AOI211_X1 g0215(.A(new_n407), .B(G20), .C1(new_n322), .C2(new_n324), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(G20), .B1(new_n403), .B2(new_n201), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT72), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n404), .B1(G159), .B2(new_n294), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n413), .A2(new_n421), .A3(new_n277), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n373), .A2(new_n281), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n423), .B1(new_n289), .B2(new_n373), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n397), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n425), .B(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n424), .ZN(new_n427));
  INV_X1    g0227(.A(G179), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n390), .A2(new_n428), .A3(new_n394), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G169), .B2(new_n396), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g0232(.A1(KEYINPUT74), .A2(KEYINPUT18), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n422), .B2(new_n424), .ZN(new_n435));
  INV_X1    g0235(.A(new_n433), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(KEYINPUT74), .A2(KEYINPUT18), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n434), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n385), .A2(new_n426), .A3(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n317), .A2(new_n365), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n288), .A2(G33), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n278), .A2(new_n281), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G107), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT25), .B1(new_n284), .B2(new_n205), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n284), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT81), .B(KEYINPUT22), .Z(new_n448));
  NAND4_X1  g0248(.A1(new_n448), .A2(new_n211), .A3(G87), .A4(new_n252), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n322), .A2(new_n324), .A3(new_n211), .A4(G87), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G116), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n211), .B2(G107), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT82), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT24), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n278), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n450), .A2(new_n451), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n450), .A2(new_n451), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n453), .A2(KEYINPUT82), .A3(new_n459), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT24), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n447), .B1(new_n462), .B2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT83), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n264), .A2(G1), .ZN(new_n472));
  AND2_X1   g0272(.A1(KEYINPUT5), .A2(G41), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(G264), .A3(new_n260), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n220), .A2(new_n253), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n221), .A2(G1698), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n322), .A2(new_n477), .A3(new_n324), .A4(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G294), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n471), .B(new_n476), .C1(new_n481), .C2(new_n260), .ZN(new_n482));
  INV_X1    g0282(.A(new_n476), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n260), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT83), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(G274), .ZN(new_n486));
  AND2_X1   g0286(.A1(G1), .A2(G13), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(new_n259), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n472), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n482), .A2(new_n485), .A3(G179), .A4(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n476), .B1(new_n481), .B2(new_n260), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n488), .A2(new_n472), .A3(new_n489), .ZN(new_n493));
  OAI21_X1  g0293(.A(G169), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n470), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n482), .A2(new_n485), .A3(new_n490), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n361), .ZN(new_n498));
  OR3_X1    g0298(.A1(new_n492), .A2(G190), .A3(new_n493), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n496), .B1(new_n470), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n475), .A2(G257), .A3(new_n260), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n490), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n322), .A2(new_n324), .A3(G244), .A4(new_n253), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n253), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n322), .A2(new_n324), .A3(G250), .A4(G1698), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G283), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n506), .A2(new_n507), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n503), .B1(new_n510), .B2(new_n261), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n361), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT6), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n513), .A2(new_n204), .A3(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(G97), .B(G107), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n514), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n516), .A2(new_n211), .B1(new_n255), .B2(new_n295), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n205), .B1(new_n408), .B2(new_n411), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n277), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n281), .A2(G97), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n443), .B2(G97), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n511), .A2(G190), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n508), .B(new_n509), .C1(new_n504), .C2(new_n505), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n504), .A2(new_n505), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n261), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(new_n503), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(G179), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n274), .B2(new_n511), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n523), .A2(new_n524), .B1(new_n522), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n475), .A2(new_n260), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n493), .B1(new_n533), .B2(G270), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n252), .A2(G264), .A3(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n252), .A2(G257), .A3(new_n253), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n414), .A2(G303), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n261), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT20), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n541), .A2(KEYINPUT79), .ZN(new_n542));
  INV_X1    g0342(.A(G116), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n276), .A2(new_n210), .B1(G20), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n509), .B(new_n211), .C1(G33), .C2(new_n204), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT79), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(KEYINPUT20), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n544), .A2(KEYINPUT79), .A3(new_n545), .A4(new_n541), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n285), .A2(G116), .A3(new_n442), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT78), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n281), .B2(G116), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n284), .A2(KEYINPUT78), .A3(new_n543), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n548), .A2(new_n549), .A3(new_n550), .A4(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n540), .A2(new_n555), .A3(KEYINPUT21), .A4(G169), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n555), .A2(G179), .A3(new_n539), .A4(new_n534), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n274), .B1(new_n534), .B2(new_n539), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT21), .B1(new_n559), .B2(new_n555), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT80), .ZN(new_n562));
  INV_X1    g0362(.A(new_n555), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n534), .A2(new_n539), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n564), .C2(new_n361), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n361), .B1(new_n534), .B2(new_n539), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT80), .B1(new_n566), .B2(new_n555), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(G190), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n561), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n211), .B1(new_n319), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(G87), .B2(new_n206), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n322), .A2(new_n324), .A3(new_n211), .A4(G68), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n571), .B1(new_n292), .B2(new_n204), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n277), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n375), .A2(new_n284), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n579), .B1(G87), .B2(new_n443), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n488), .A2(new_n472), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n260), .B(G250), .C1(G1), .C2(new_n264), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(G244), .A2(G1698), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n322), .A2(new_n324), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT75), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n252), .A2(G238), .A3(new_n253), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT75), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n322), .A2(new_n324), .A3(new_n584), .A4(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n454), .A4(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n583), .B1(new_n590), .B2(new_n261), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT77), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n594), .A3(G190), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n591), .B2(G190), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n580), .B(new_n593), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(new_n274), .ZN(new_n599));
  INV_X1    g0399(.A(new_n375), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n443), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n577), .A2(new_n601), .A3(new_n578), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT76), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n591), .A2(new_n428), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT76), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n577), .A2(new_n601), .A3(new_n605), .A4(new_n578), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n599), .A2(new_n603), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n570), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n441), .A2(new_n501), .A3(new_n531), .A4(new_n609), .ZN(new_n610));
  XOR2_X1   g0410(.A(new_n610), .B(KEYINPUT84), .Z(G372));
  AND3_X1   g0411(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n612));
  INV_X1    g0412(.A(new_n583), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  AND3_X1   g0414(.A1(new_n590), .A2(new_n614), .A3(new_n261), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(new_n590), .B2(new_n261), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n274), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n612), .A2(KEYINPUT87), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(KEYINPUT87), .B1(new_n612), .B2(new_n618), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n559), .A2(new_n555), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT21), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n557), .A3(new_n556), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n496), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n470), .A2(new_n500), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n617), .A2(G200), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n590), .A2(new_n261), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n630), .A2(G190), .A3(new_n613), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT77), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n595), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n629), .A2(new_n633), .A3(new_n580), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n612), .A2(new_n618), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n531), .A2(new_n628), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT86), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n627), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n580), .B1(new_n596), .B2(new_n597), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n630), .A2(KEYINPUT85), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n590), .A2(new_n614), .A3(new_n261), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n583), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n361), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(G169), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n639), .A2(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n647), .A2(KEYINPUT86), .A3(new_n628), .A4(new_n531), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n622), .B1(new_n638), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT88), .ZN(new_n651));
  AOI211_X1 g0451(.A(new_n428), .B(new_n503), .C1(new_n510), .C2(new_n261), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n274), .B1(new_n527), .B2(new_n528), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n529), .B(KEYINPUT88), .C1(new_n274), .C2(new_n511), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n522), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n650), .B1(new_n646), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n530), .A2(new_n522), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n598), .A2(new_n660), .A3(new_n607), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(new_n650), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT89), .B(new_n650), .C1(new_n646), .C2(new_n656), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n649), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n441), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n307), .A2(new_n312), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT10), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n314), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT17), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n425), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n364), .A2(new_n381), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n671), .B1(new_n672), .B2(new_n357), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT18), .ZN(new_n674));
  AOI211_X1 g0474(.A(KEYINPUT90), .B(new_n430), .C1(new_n422), .C2(new_n424), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n427), .B2(new_n431), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n674), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n285), .A2(new_n286), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n346), .B(new_n373), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n423), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n417), .A2(new_n420), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n278), .B1(new_n684), .B2(new_n398), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n685), .B2(new_n421), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT90), .B1(new_n686), .B2(new_n430), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n435), .A2(new_n676), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(KEYINPUT18), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n678), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n669), .B1(new_n673), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n692), .A2(new_n302), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n666), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n694), .B(KEYINPUT91), .ZN(G369));
  NAND2_X1  g0495(.A1(new_n280), .A2(new_n211), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(G213), .ZN(new_n699));
  INV_X1    g0499(.A(G343), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n563), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n626), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n570), .B2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n496), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(new_n628), .C1(new_n470), .C2(new_n702), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n708), .B2(new_n702), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n561), .A2(new_n701), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n501), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n496), .A2(new_n702), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n711), .A2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n215), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n208), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n654), .A2(new_n522), .A3(new_n655), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(KEYINPUT26), .A3(new_n635), .A4(new_n634), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n661), .A2(new_n650), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n728), .B(new_n621), .C1(new_n636), .C2(new_n627), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n729), .A2(KEYINPUT95), .A3(KEYINPUT29), .A4(new_n702), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n726), .A2(new_n727), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n621), .B1(new_n636), .B2(new_n627), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT29), .B(new_n702), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n701), .B1(new_n649), .B2(new_n664), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n730), .B(new_n735), .C1(new_n736), .C2(KEYINPUT29), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n609), .A2(new_n501), .A3(new_n531), .A4(new_n702), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n591), .A2(new_n485), .A3(new_n482), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT92), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n534), .A2(new_n539), .A3(G179), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n739), .A2(new_n740), .A3(new_n742), .A4(new_n511), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n511), .A2(new_n591), .A3(new_n485), .A4(new_n482), .ZN(new_n744));
  OAI21_X1  g0544(.A(KEYINPUT92), .B1(new_n744), .B2(new_n741), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT93), .B(KEYINPUT30), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n511), .ZN(new_n748));
  AOI21_X1  g0548(.A(G179), .B1(new_n534), .B2(new_n539), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n617), .A2(new_n497), .A3(new_n748), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n739), .A2(KEYINPUT30), .A3(new_n742), .A4(new_n511), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g0552(.A(KEYINPUT31), .B(new_n701), .C1(new_n747), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT94), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n747), .A2(KEYINPUT94), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n702), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n738), .B(new_n753), .C1(new_n758), .C2(KEYINPUT31), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n737), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n724), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(G13), .A2(G33), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(G20), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n210), .B1(G20), .B2(new_n274), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n250), .A2(new_n264), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n718), .A2(new_n252), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(new_n264), .B2(new_n209), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n770), .B1(KEYINPUT96), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n774), .B1(KEYINPUT96), .B2(new_n773), .ZN(new_n775));
  INV_X1    g0575(.A(G355), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n252), .A2(new_n215), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n775), .B1(G116), .B2(new_n215), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n769), .B1(new_n778), .B2(KEYINPUT97), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(KEYINPUT97), .B2(new_n778), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n279), .A2(G20), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n288), .B1(new_n781), .B2(G45), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n719), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n768), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n211), .A2(new_n428), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n361), .A2(G190), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G322), .A2(new_n790), .B1(new_n793), .B2(G311), .ZN(new_n794));
  INV_X1    g0594(.A(G303), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n359), .A2(new_n361), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n211), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n794), .B(new_n414), .C1(new_n795), .C2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n361), .A2(G190), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n787), .A2(new_n800), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(KEYINPUT33), .B(G317), .Z(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n787), .A2(new_n796), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT102), .Z(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n799), .B(new_n807), .C1(G326), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n797), .A2(new_n791), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT98), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n797), .A2(new_n800), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n816), .A2(G329), .B1(G283), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(KEYINPUT103), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  OAI21_X1  g0621(.A(G20), .B1(new_n789), .B2(G179), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT100), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n822), .A2(new_n823), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n811), .B(new_n820), .C1(new_n821), .C2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n252), .B1(new_n817), .B2(new_n205), .ZN(new_n829));
  INV_X1    g0629(.A(new_n808), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G50), .A2(new_n830), .B1(new_n793), .B2(G77), .ZN(new_n831));
  INV_X1    g0631(.A(G58), .ZN(new_n832));
  INV_X1    g0632(.A(new_n790), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .C1(new_n219), .C2(new_n798), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n829), .B(new_n834), .C1(G68), .C2(new_n804), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n827), .A2(KEYINPUT101), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n827), .A2(KEYINPUT101), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G97), .ZN(new_n840));
  INV_X1    g0640(.A(G159), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n815), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT32), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n835), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n786), .B1(new_n828), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g0645(.A1(new_n780), .A2(new_n785), .A3(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n767), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n705), .B2(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n707), .A2(new_n784), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(G330), .B2(new_n705), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G396));
  NAND2_X1  g0652(.A1(new_n385), .A2(new_n702), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n649), .B2(new_n664), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n380), .A2(new_n701), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n384), .A2(new_n382), .B1(new_n379), .B2(new_n701), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n381), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n736), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n784), .B1(new_n861), .B2(new_n761), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n761), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n768), .A2(new_n765), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n784), .B1(G77), .B2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT104), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n804), .A2(KEYINPUT105), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n804), .A2(KEYINPUT105), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(G283), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(G311), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n815), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n414), .B1(new_n808), .B2(new_n795), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G294), .A2(new_n790), .B1(new_n793), .B2(G116), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n818), .A2(G87), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n876), .B(new_n877), .C1(new_n205), .C2(new_n798), .ZN(new_n878));
  NOR4_X1   g0678(.A1(new_n872), .A2(new_n874), .A3(new_n875), .A4(new_n878), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G137), .A2(new_n830), .B1(new_n793), .B2(G159), .ZN(new_n880));
  INV_X1    g0680(.A(G143), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n880), .B1(new_n881), .B2(new_n833), .C1(new_n805), .C2(new_n293), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT34), .ZN(new_n883));
  INV_X1    g0683(.A(G132), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n252), .B1(new_n815), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n818), .A2(G68), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n244), .B2(new_n798), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT106), .ZN(new_n888));
  INV_X1    g0688(.A(new_n827), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n885), .B(new_n888), .C1(G58), .C2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n879), .A2(new_n840), .B1(new_n883), .B2(new_n890), .ZN(new_n891));
  OAI221_X1 g0691(.A(new_n867), .B1(new_n860), .B2(new_n766), .C1(new_n891), .C2(new_n786), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n863), .A2(new_n892), .ZN(G384));
  NOR2_X1   g0693(.A1(new_n781), .A2(new_n288), .ZN(new_n894));
  INV_X1    g0694(.A(G330), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT108), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n675), .A2(new_n677), .A3(new_n674), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT18), .B1(new_n687), .B2(new_n688), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n426), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT107), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n686), .B2(new_n699), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n699), .B1(new_n422), .B2(new_n424), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(KEYINPUT107), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n425), .B1(new_n675), .B2(new_n677), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n905), .B2(new_n904), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n902), .B(new_n900), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT37), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n432), .A2(new_n908), .A3(new_n425), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n899), .A2(new_n904), .B1(new_n906), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n896), .B1(new_n912), .B2(KEYINPUT38), .ZN(new_n913));
  INV_X1    g0713(.A(new_n437), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n438), .B1(new_n435), .B2(new_n436), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n902), .B1(new_n916), .B2(new_n671), .ZN(new_n917));
  INV_X1    g0717(.A(new_n902), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n425), .A3(new_n432), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT37), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n904), .B2(new_n909), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n917), .A2(new_n921), .A3(KEYINPUT38), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n687), .A2(new_n688), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n907), .A2(new_n924), .A3(new_n425), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n925), .A2(KEYINPUT37), .B1(new_n907), .B2(new_n910), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n907), .B1(new_n690), .B2(new_n426), .ZN(new_n927));
  OAI211_X1 g0727(.A(KEYINPUT108), .B(new_n923), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n913), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n356), .A2(new_n701), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n357), .A2(new_n364), .A3(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n356), .B(new_n701), .C1(new_n345), .C2(new_n363), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n859), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n738), .B1(new_n758), .B2(KEYINPUT31), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT31), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n935), .B(new_n702), .C1(new_n756), .C2(new_n757), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n933), .B(KEYINPUT40), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n929), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(KEYINPUT109), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT109), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n929), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT40), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n933), .B1(new_n934), .B2(new_n936), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n907), .A2(new_n910), .B1(new_n919), .B2(KEYINPUT37), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n918), .B1(new_n439), .B2(new_n426), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n923), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n948), .A2(new_n922), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n944), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n934), .A2(new_n936), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n441), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n895), .B1(new_n951), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n951), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n931), .A2(new_n932), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n854), .B2(new_n856), .ZN(new_n957));
  INV_X1    g0757(.A(new_n699), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n957), .A2(new_n949), .B1(new_n690), .B2(new_n958), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n948), .A2(KEYINPUT39), .A3(new_n922), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT39), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n929), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n345), .A2(new_n356), .A3(new_n702), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n959), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n441), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n693), .B1(new_n737), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n965), .B(new_n967), .Z(new_n968));
  AOI21_X1  g0768(.A(new_n894), .B1(new_n955), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n968), .B2(new_n955), .ZN(new_n970));
  INV_X1    g0770(.A(new_n516), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT35), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(KEYINPUT35), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n972), .A2(G116), .A3(new_n212), .A4(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT36), .ZN(new_n975));
  OAI21_X1  g0775(.A(G77), .B1(new_n832), .B2(new_n246), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n245), .B1(new_n208), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(G1), .A3(new_n279), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n970), .A2(new_n975), .A3(new_n978), .ZN(G367));
  NOR2_X1   g0779(.A1(new_n838), .A2(new_n246), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n809), .A2(new_n881), .B1(new_n293), .B2(new_n833), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n982), .A2(KEYINPUT117), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(KEYINPUT117), .ZN(new_n984));
  INV_X1    g0784(.A(G137), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n815), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n414), .B1(new_n818), .B2(G77), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n244), .B2(new_n792), .C1(new_n832), .C2(new_n798), .ZN(new_n988));
  INV_X1    g0788(.A(new_n870), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n986), .B(new_n988), .C1(new_n989), .C2(G159), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n983), .A2(new_n984), .A3(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT118), .ZN(new_n992));
  INV_X1    g0792(.A(new_n798), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT46), .B1(new_n993), .B2(G116), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n810), .A2(G311), .B1(KEYINPUT116), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(G317), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(KEYINPUT116), .B2(new_n994), .C1(new_n996), .C2(new_n815), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n252), .B1(new_n790), .B2(G303), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n993), .A2(KEYINPUT46), .A3(G116), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n204), .C2(new_n817), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n821), .B2(new_n870), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n827), .A2(new_n205), .B1(new_n871), .B2(new_n792), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT115), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n992), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n768), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n580), .A2(new_n702), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n622), .A2(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1009), .A2(KEYINPUT110), .B1(new_n646), .B2(new_n1008), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(KEYINPUT110), .B2(new_n1009), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n767), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n239), .A2(new_n771), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n769), .C1(new_n215), .C2(new_n375), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1007), .A2(new_n784), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n725), .A2(new_n701), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n522), .A2(new_n701), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n531), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n713), .A2(new_n714), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n716), .C2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1019), .ZN(new_n1025));
  OR2_X1    g0825(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n715), .A2(new_n1024), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1022), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n711), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT112), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT112), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1028), .A2(new_n1032), .A3(new_n1029), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n706), .A2(KEYINPUT113), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n713), .C1(new_n710), .C2(new_n712), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n706), .A2(KEYINPUT113), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1037), .B(new_n1038), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n763), .B1(new_n1035), .B2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n719), .B(KEYINPUT41), .Z(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(KEYINPUT114), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT114), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1040), .A2(new_n1045), .A3(new_n1042), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n783), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1025), .A2(new_n713), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT42), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1025), .A2(new_n708), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n702), .B1(new_n1050), .B2(new_n660), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT43), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n1011), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1011), .A2(new_n1053), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n711), .A2(new_n1025), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1056), .B(new_n1057), .Z(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1015), .B1(new_n1047), .B2(new_n1059), .ZN(G387));
  INV_X1    g0860(.A(new_n1039), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n783), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n833), .A2(new_n996), .B1(new_n792), .B2(new_n795), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n810), .B2(G322), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1064), .B1(new_n870), .B2(new_n873), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(new_n889), .A2(G283), .B1(G294), .B2(new_n993), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT121), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n816), .A2(G326), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n252), .B1(new_n818), .B2(G116), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n798), .A2(new_n255), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G159), .B2(new_n830), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n244), .B2(new_n833), .C1(new_n246), .C2(new_n792), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n414), .B(new_n1079), .C1(G97), .C2(new_n818), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n839), .A2(new_n600), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n373), .A2(new_n804), .B1(new_n816), .B2(G150), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n786), .B1(new_n1076), .B2(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n777), .A2(new_n721), .B1(G107), .B2(new_n215), .ZN(new_n1085));
  XNOR2_X1  g0885(.A(new_n1085), .B(KEYINPUT119), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n236), .A2(G45), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n721), .ZN(new_n1088));
  AOI211_X1 g0888(.A(G45), .B(new_n1088), .C1(G68), .C2(G77), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n291), .A2(G50), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT50), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n772), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1086), .B1(new_n1087), .B2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(KEYINPUT120), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n769), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n784), .B1(new_n1094), .B2(new_n1096), .C1(new_n710), .C2(new_n847), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1061), .A2(new_n763), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n719), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1061), .A2(new_n763), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n1062), .B1(new_n1084), .B2(new_n1097), .C1(new_n1099), .C2(new_n1100), .ZN(G393));
  NAND3_X1  g0901(.A1(new_n1034), .A2(new_n783), .A3(new_n1030), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n769), .B1(new_n204), .B2(new_n215), .C1(new_n243), .C2(new_n772), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n784), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n790), .A2(G311), .B1(new_n830), .B2(G317), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(KEYINPUT52), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n414), .B1(new_n817), .B2(new_n205), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n871), .A2(new_n798), .B1(new_n792), .B2(new_n821), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n816), .A2(G322), .B1(new_n1105), .B2(KEYINPUT52), .ZN(new_n1110));
  AND2_X1   g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n543), .B2(new_n827), .C1(new_n795), .C2(new_n870), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n833), .A2(new_n841), .B1(new_n808), .B2(new_n293), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT122), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT51), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G68), .A2(new_n993), .B1(new_n793), .B2(new_n373), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1116), .A2(new_n252), .A3(new_n877), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G143), .B2(new_n816), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1115), .B(new_n1118), .C1(new_n244), .C2(new_n870), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n838), .A2(new_n255), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1112), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1104), .B1(new_n1121), .B2(new_n768), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(new_n847), .B2(new_n1019), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1102), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1034), .A2(new_n1030), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1098), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT123), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1098), .A2(new_n1126), .A3(KEYINPUT123), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1035), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1098), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n720), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(KEYINPUT124), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT124), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1125), .B1(new_n1136), .B2(new_n1137), .ZN(G390));
  OAI211_X1 g0938(.A(new_n933), .B(G330), .C1(new_n934), .C2(new_n936), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n928), .A2(new_n922), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n899), .A2(new_n904), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n906), .A2(new_n911), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT108), .B1(new_n1144), .B2(new_n923), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n961), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n960), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1146), .A2(new_n1147), .B1(new_n963), .B2(new_n957), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n858), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n380), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n702), .B(new_n1150), .C1(new_n731), .C2(new_n732), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT125), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n1151), .A2(new_n1152), .A3(new_n857), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1152), .B1(new_n1151), .B2(new_n857), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n956), .ZN(new_n1155));
  NOR3_X1   g0955(.A1(new_n1153), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n963), .B1(new_n1141), .B2(new_n1145), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1140), .B1(new_n1148), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1151), .A2(new_n857), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1160), .A2(KEYINPUT125), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1151), .A2(new_n1152), .A3(new_n857), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n956), .A3(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1163), .A2(new_n963), .A3(new_n929), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n760), .A2(new_n860), .A3(new_n956), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n957), .A2(new_n963), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1164), .B(new_n1165), .C1(new_n962), .C2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1159), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n952), .A2(G330), .A3(new_n441), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n693), .B(new_n1169), .C1(new_n737), .C2(new_n966), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n956), .B1(new_n760), .B2(new_n860), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n1171), .A2(new_n1140), .B1(new_n854), .B2(new_n856), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n860), .B(G330), .C1(new_n934), .C2(new_n936), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1155), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1165), .B(new_n1174), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1170), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1159), .A2(new_n1176), .A3(new_n1167), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n719), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1159), .A2(new_n783), .A3(new_n1167), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n784), .B1(new_n373), .B2(new_n865), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n790), .A2(G132), .B1(new_n818), .B2(G50), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n830), .A2(G128), .ZN(new_n1184));
  INV_X1    g0984(.A(G125), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1183), .B(new_n1184), .C1(new_n815), .C2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(KEYINPUT54), .B(G143), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n414), .B1(new_n793), .B2(new_n1188), .ZN(new_n1189));
  OR3_X1    g0989(.A1(new_n798), .A2(KEYINPUT53), .A3(new_n293), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT53), .B1(new_n798), .B2(new_n293), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1186), .A2(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n985), .B2(new_n870), .C1(new_n841), .C2(new_n838), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n886), .B1(new_n815), .B2(new_n821), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n989), .A2(G107), .B1(KEYINPUT126), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n414), .B1(new_n798), .B2(new_n219), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n808), .A2(new_n871), .B1(new_n792), .B2(new_n204), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1197), .B(new_n1198), .C1(G116), .C2(new_n790), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1196), .B(new_n1199), .C1(KEYINPUT126), .C2(new_n1195), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1194), .B1(new_n1200), .B2(new_n1120), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1182), .B1(new_n1201), .B2(new_n768), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n962), .B2(new_n766), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1181), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1180), .A2(new_n1204), .ZN(G378));
  INV_X1    g1005(.A(new_n965), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n317), .A2(new_n301), .A3(new_n958), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n301), .A2(new_n958), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n669), .A2(new_n302), .A3(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n1207), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AND2_X1   g1014(.A1(new_n950), .A2(G330), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1214), .B1(new_n943), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n950), .A2(G330), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1217), .B(new_n1213), .C1(new_n940), .C2(new_n942), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1206), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n929), .A2(new_n941), .A3(new_n938), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n941), .B1(new_n929), .B2(new_n938), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1215), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(new_n1213), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1214), .B(new_n1215), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1223), .A2(new_n965), .A3(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1219), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1213), .A2(new_n765), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n833), .A2(new_n205), .B1(new_n832), .B2(new_n817), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n808), .A2(new_n543), .B1(new_n792), .B2(new_n375), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n414), .A2(new_n263), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1077), .A4(new_n1230), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1231), .B1(new_n204), .B2(new_n805), .C1(new_n871), .C2(new_n815), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1232), .A2(new_n980), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT58), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT58), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n321), .A2(new_n263), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1230), .A2(new_n244), .A3(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n816), .A2(G124), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1236), .B1(new_n818), .B2(G159), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G128), .A2(new_n790), .B1(new_n793), .B2(G137), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G125), .A2(new_n830), .B1(new_n993), .B2(new_n1188), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1241), .B(new_n1242), .C1(new_n805), .C2(new_n884), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n839), .B2(G150), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT59), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1239), .B(new_n1240), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1245), .B2(new_n1244), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n768), .B1(new_n1238), .B2(new_n1247), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT127), .Z(new_n1249));
  AOI211_X1 g1049(.A(new_n785), .B(new_n1249), .C1(new_n244), .C2(new_n864), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1226), .A2(new_n783), .B1(new_n1227), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1170), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1179), .A2(new_n1252), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1223), .A2(new_n965), .A3(new_n1224), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n965), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT57), .B(new_n1253), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n719), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1253), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1251), .B1(new_n1257), .B2(new_n1258), .ZN(G375));
  NAND2_X1  g1059(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1170), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1042), .A3(new_n1177), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1155), .A2(new_n765), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(G294), .A2(new_n830), .B1(new_n993), .B2(G97), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(G283), .A2(new_n790), .B1(new_n793), .B2(G107), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n252), .B1(new_n818), .B2(G77), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G303), .B2(new_n816), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1081), .B(new_n1269), .C1(new_n543), .C2(new_n870), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(G132), .A2(new_n830), .B1(new_n993), .B2(G159), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G137), .A2(new_n790), .B1(new_n793), .B2(G150), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n414), .B1(new_n818), .B2(G58), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1274), .B1(G128), .B2(new_n816), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n838), .B2(new_n244), .C1(new_n870), .C2(new_n1187), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n786), .B1(new_n1270), .B2(new_n1276), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n785), .B(new_n1277), .C1(new_n246), .C2(new_n864), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1260), .A2(new_n783), .B1(new_n1264), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1263), .A2(new_n1279), .ZN(G381));
  NAND2_X1  g1080(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT124), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1124), .B1(new_n1283), .B2(new_n1135), .ZN(new_n1284));
  NOR4_X1   g1084(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OR4_X1    g1086(.A1(G387), .A2(G375), .A3(new_n1286), .A4(G378), .ZN(G407));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n700), .A2(G213), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  OAI211_X1 g1091(.A(G407), .B(G213), .C1(G375), .C2(new_n1291), .ZN(G409));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G378), .B(new_n1251), .C1(new_n1257), .C2(new_n1258), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n783), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1250), .A2(new_n1227), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1253), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1297));
  OAI211_X1 g1097(.A(new_n1295), .B(new_n1296), .C1(new_n1297), .C2(new_n1041), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1288), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1290), .B1(new_n1294), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1262), .B1(new_n1301), .B2(new_n1176), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1260), .A2(new_n1252), .A3(new_n1301), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1303), .A2(new_n720), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1305), .A2(G384), .A3(new_n1279), .ZN(new_n1306));
  AOI21_X1  g1106(.A(G384), .B1(new_n1305), .B2(new_n1279), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G2897), .B(new_n1290), .C1(new_n1306), .C2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1307), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1305), .A2(G384), .A3(new_n1279), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(G2897), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1293), .B1(new_n1300), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1300), .A2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT63), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1046), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1045), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n782), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(new_n1058), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(G390), .A2(new_n1323), .A3(new_n1015), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G387), .A2(new_n1284), .ZN(new_n1325));
  XNOR2_X1  g1125(.A(G393), .B(new_n851), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1326), .B1(new_n1324), .B2(new_n1325), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1316), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1315), .A2(new_n1319), .A3(new_n1329), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  AND3_X1   g1132(.A1(new_n1300), .A2(new_n1332), .A3(new_n1316), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1332), .B1(new_n1300), .B2(new_n1316), .ZN(new_n1334));
  NOR3_X1   g1134(.A1(new_n1333), .A2(new_n1314), .A3(new_n1334), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1331), .B1(new_n1335), .B2(new_n1329), .ZN(G405));
  NAND2_X1  g1136(.A1(G375), .A2(new_n1288), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1316), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1337), .A2(new_n1294), .A3(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1338), .B1(new_n1337), .B2(new_n1294), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(new_n1342), .B(new_n1329), .ZN(G402));
endmodule


