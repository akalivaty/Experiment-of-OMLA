//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n554, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1139, new_n1140;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT66), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT67), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT68), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT69), .ZN(G319));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  AND2_X1   g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n459), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n460), .A2(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT70), .B(G2104), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n465), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT71), .Z(G160));
  XOR2_X1   g050(.A(new_n471), .B(KEYINPUT72), .Z(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n480), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n479), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  NAND3_X1  g062(.A1(new_n480), .A2(G102), .A3(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n490), .B1(new_n471), .B2(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n491), .B2(new_n480), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n480), .A2(KEYINPUT4), .A3(G138), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n459), .B(new_n493), .C1(new_n472), .C2(new_n458), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n459), .A2(new_n461), .A3(G138), .A4(new_n480), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n492), .A2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  AND3_X1   g076(.A1(new_n501), .A2(KEYINPUT74), .A3(G543), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT74), .B1(new_n501), .B2(G543), .ZN(new_n503));
  OAI22_X1  g078(.A1(new_n502), .A2(new_n503), .B1(new_n501), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  XOR2_X1   g081(.A(KEYINPUT73), .B(G651), .Z(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  XOR2_X1   g084(.A(new_n509), .B(KEYINPUT76), .Z(new_n510));
  INV_X1    g085(.A(new_n504), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT6), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n511), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n514), .A2(G543), .A3(new_n513), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n515), .A2(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT75), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n519), .A2(new_n520), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n510), .B1(new_n521), .B2(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  NAND2_X1  g099(.A1(new_n514), .A2(new_n513), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n504), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  INV_X1    g102(.A(new_n518), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n527), .A2(new_n529), .A3(new_n530), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n504), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(new_n508), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n511), .A2(G90), .A3(new_n513), .A4(new_n514), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n514), .A2(G52), .A3(G543), .A4(new_n513), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n526), .A2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n528), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n504), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(new_n508), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n545), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND3_X1  g133(.A1(new_n528), .A2(KEYINPUT9), .A3(G53), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n526), .A2(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n504), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n518), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n559), .A2(new_n560), .A3(new_n564), .A4(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  NAND2_X1  g144(.A1(new_n526), .A2(G87), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n528), .A2(G49), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(G288));
  INV_X1    g148(.A(G86), .ZN(new_n574));
  INV_X1    g149(.A(G48), .ZN(new_n575));
  OAI22_X1  g150(.A1(new_n515), .A2(new_n574), .B1(new_n575), .B2(new_n518), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n507), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(G85), .A2(new_n526), .B1(new_n528), .B2(G47), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n507), .B2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n526), .A2(KEYINPUT10), .A3(G92), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n515), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n591), .A2(G54), .A3(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G651), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n590), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n584), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n584), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  XOR2_X1   g176(.A(new_n601), .B(KEYINPUT79), .Z(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g186(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(KEYINPUT81), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n613), .B(new_n614), .C1(G111), .C2(new_n480), .ZN(new_n615));
  INV_X1    g190(.A(G135), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n481), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(G123), .B2(new_n478), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT82), .Z(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2096), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n462), .A2(new_n472), .A3(new_n480), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT83), .B(KEYINPUT14), .Z(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  NOR2_X1   g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT84), .Z(new_n640));
  INV_X1    g215(.A(G14), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n641), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(G401));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT85), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT86), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT87), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n647), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n653), .B2(new_n649), .ZN(new_n655));
  OR3_X1    g230(.A1(new_n651), .A2(new_n653), .A3(new_n646), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n647), .A2(new_n649), .A3(new_n653), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT88), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2096), .ZN(new_n661));
  INV_X1    g236(.A(G2100), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT89), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT19), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n670), .A2(new_n671), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT91), .Z(new_n678));
  NOR2_X1   g253(.A1(new_n672), .A2(new_n676), .ZN(new_n679));
  AOI211_X1 g254(.A(new_n675), .B(new_n678), .C1(new_n668), .C2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1991), .B(G1996), .ZN(new_n681));
  INV_X1    g256(.A(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n680), .B(new_n685), .Z(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT92), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G229));
  MUX2_X1   g264(.A(G24), .B(G290), .S(G16), .Z(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G1986), .Z(new_n691));
  NOR2_X1   g266(.A1(G25), .A2(G29), .ZN(new_n692));
  OR2_X1    g267(.A1(G95), .A2(G2105), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n693), .B(G2104), .C1(G107), .C2(new_n480), .ZN(new_n694));
  INV_X1    g269(.A(G119), .ZN(new_n695));
  INV_X1    g270(.A(G131), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n694), .B1(new_n477), .B2(new_n695), .C1(new_n696), .C2(new_n481), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n692), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT35), .B(G1991), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G16), .A2(G23), .ZN(new_n707));
  INV_X1    g282(.A(G288), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n702), .A2(G6), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n579), .B2(new_n702), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT32), .B(G1981), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n706), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT34), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n691), .B(new_n701), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  NOR2_X1   g296(.A1(G29), .A2(G35), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G162), .B2(G29), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT29), .ZN(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT28), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n728), .A2(G26), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n731));
  INV_X1    g306(.A(G128), .ZN(new_n732));
  INV_X1    g307(.A(G140), .ZN(new_n733));
  OAI221_X1 g308(.A(new_n731), .B1(new_n477), .B2(new_n732), .C1(new_n733), .C2(new_n481), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n727), .B(new_n729), .C1(new_n734), .C2(G29), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n727), .B2(new_n729), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT95), .B(G2067), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n702), .A2(G4), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n598), .B2(new_n702), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(G16), .A2(G19), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n552), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT94), .B(G1341), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n738), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT96), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n619), .A2(G29), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT24), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G34), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(G160), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n754), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(G2084), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NOR2_X1   g334(.A1(G286), .A2(new_n702), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G21), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n760), .A2(KEYINPUT99), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(KEYINPUT99), .B2(new_n760), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G1966), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n749), .A2(new_n758), .A3(new_n759), .A4(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  NAND2_X1  g342(.A1(G171), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G5), .B2(G16), .ZN(new_n769));
  OAI22_X1  g344(.A1(new_n764), .A2(G1966), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n728), .A2(G33), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n462), .A2(G127), .ZN(new_n772));
  NAND2_X1  g347(.A1(G115), .A2(G2104), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n480), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT25), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n774), .B(new_n776), .C1(new_n482), .C2(G139), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n771), .B1(new_n777), .B2(new_n728), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2072), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n769), .A2(new_n767), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n728), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n728), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(G2078), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n782), .A2(G2078), .B1(new_n728), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT100), .B(G11), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT31), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n780), .A2(new_n783), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  NOR4_X1   g363(.A1(new_n766), .A2(new_n770), .A3(new_n779), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n721), .A2(new_n726), .A3(new_n748), .A4(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n702), .A2(KEYINPUT23), .A3(G20), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT23), .ZN(new_n792));
  INV_X1    g367(.A(G20), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n793), .B2(G16), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n794), .C1(new_n603), .C2(new_n702), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT101), .B(G1956), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(G29), .A2(G32), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n482), .A2(G141), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT97), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n480), .A2(G105), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n478), .A2(G129), .B1(new_n472), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g378(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT98), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT26), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n798), .B1(new_n807), .B2(new_n728), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT27), .B(G1996), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n790), .A2(new_n797), .A3(new_n810), .ZN(G311));
  OR3_X1    g386(.A1(new_n790), .A2(new_n797), .A3(new_n810), .ZN(G150));
  NAND2_X1  g387(.A1(new_n526), .A2(G93), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT102), .B(G55), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n528), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G80), .A2(G543), .ZN(new_n817));
  INV_X1    g392(.A(G67), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n504), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n508), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(G860), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT37), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n598), .A2(G559), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT38), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT39), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT103), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n816), .B2(new_n821), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n813), .A2(new_n815), .A3(KEYINPUT103), .A4(new_n820), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n551), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n822), .A2(new_n552), .A3(KEYINPUT103), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n828), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n825), .B1(new_n835), .B2(G860), .ZN(G145));
  XNOR2_X1  g411(.A(new_n697), .B(new_n623), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n478), .A2(G130), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT106), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(new_n480), .B2(G118), .ZN(new_n841));
  INV_X1    g416(.A(G106), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n480), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n482), .B2(G142), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n837), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT107), .ZN(new_n847));
  OAI211_X1 g422(.A(G126), .B(new_n459), .C1(new_n472), .C2(new_n458), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n489), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G2105), .ZN(new_n850));
  AND3_X1   g425(.A1(new_n494), .A2(new_n497), .A3(KEYINPUT105), .ZN(new_n851));
  AOI21_X1  g426(.A(KEYINPUT105), .B1(new_n494), .B2(new_n497), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n850), .B(new_n488), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n734), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n807), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n777), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n856), .A2(new_n777), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n847), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n857), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n846), .B(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n486), .B(KEYINPUT104), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G160), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n619), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(new_n846), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n859), .A2(new_n870), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g448(.A(new_n834), .B(new_n608), .ZN(new_n874));
  AND4_X1   g449(.A1(G299), .A2(new_n589), .A3(new_n596), .A4(new_n593), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n603), .B1(new_n590), .B2(new_n597), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n593), .A2(new_n596), .ZN(new_n880));
  AOI21_X1  g455(.A(G299), .B1(new_n880), .B2(new_n589), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT108), .B1(new_n881), .B2(new_n875), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n877), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n878), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n879), .B1(new_n888), .B2(new_n874), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(G288), .A2(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g467(.A1(G288), .A2(KEYINPUT109), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n894), .B(G290), .Z(new_n895));
  NAND2_X1  g470(.A1(G303), .A2(new_n579), .ZN(new_n896));
  OAI211_X1 g471(.A(G305), .B(new_n510), .C1(new_n521), .C2(new_n522), .ZN(new_n897));
  AOI21_X1  g472(.A(KEYINPUT110), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n895), .A2(new_n899), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n896), .A2(new_n897), .A3(KEYINPUT110), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n898), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n900), .B1(new_n895), .B2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n891), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(G868), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(G868), .B2(new_n822), .ZN(G295));
  OAI21_X1  g481(.A(new_n905), .B1(G868), .B2(new_n822), .ZN(G331));
  NAND2_X1  g482(.A1(new_n902), .A2(new_n895), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n899), .B2(new_n895), .ZN(new_n909));
  INV_X1    g484(.A(new_n878), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n882), .A2(new_n884), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .ZN(new_n912));
  NAND3_X1  g487(.A1(G168), .A2(G171), .A3(KEYINPUT112), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT112), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n914), .B1(new_n540), .B2(new_n543), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n539), .A2(new_n541), .A3(KEYINPUT112), .A4(new_n542), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n915), .A2(G286), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n834), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n832), .A2(new_n913), .A3(new_n833), .A4(new_n917), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT114), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(KEYINPUT114), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n912), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n919), .A2(new_n920), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n910), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n912), .B(KEYINPUT41), .C1(new_n921), .C2(new_n922), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n909), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n885), .B2(new_n887), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT113), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n921), .A2(new_n922), .A3(new_n910), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT113), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n932), .B(new_n924), .C1(new_n885), .C2(new_n887), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n903), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  INV_X1    g510(.A(G37), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n928), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n937), .A2(KEYINPUT116), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(KEYINPUT116), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n909), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT115), .B1(new_n941), .B2(new_n936), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT115), .ZN(new_n943));
  AOI211_X1 g518(.A(new_n943), .B(G37), .C1(new_n940), .C2(new_n909), .ZN(new_n944));
  INV_X1    g519(.A(new_n934), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI211_X1 g521(.A(new_n938), .B(new_n939), .C1(new_n946), .C2(new_n935), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n946), .A2(KEYINPUT43), .ZN(new_n950));
  AND4_X1   g525(.A1(KEYINPUT43), .A2(new_n928), .A3(new_n936), .A4(new_n934), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT44), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(G397));
  INV_X1    g528(.A(G1384), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n851), .A2(new_n852), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n954), .B1(new_n955), .B2(new_n492), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G40), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n474), .A2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n957), .A2(new_n959), .A3(KEYINPUT45), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n734), .B(G2067), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(new_n807), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n963));
  INV_X1    g538(.A(G1996), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n960), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n966), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n962), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT47), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n807), .A2(G1996), .A3(new_n960), .ZN(new_n970));
  XOR2_X1   g545(.A(new_n970), .B(KEYINPUT117), .Z(new_n971));
  NOR2_X1   g546(.A1(new_n807), .A2(G1996), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n960), .B1(new_n972), .B2(new_n961), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n697), .B(new_n700), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n974), .B1(new_n960), .B2(new_n975), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n977), .B(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT126), .ZN(new_n981));
  INV_X1    g556(.A(new_n698), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n700), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n973), .A3(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n734), .A2(G2067), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n981), .B1(new_n986), .B2(new_n960), .ZN(new_n987));
  AOI211_X1 g562(.A(KEYINPUT126), .B(new_n966), .C1(new_n984), .C2(new_n985), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n969), .B(new_n980), .C1(new_n987), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(G305), .A2(G1981), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n579), .A2(new_n682), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n993), .A2(KEYINPUT49), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(KEYINPUT49), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n956), .A2(KEYINPUT118), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT118), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n853), .A2(new_n997), .A3(new_n954), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n959), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G8), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n994), .A2(new_n995), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1976), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n708), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n992), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(new_n1001), .ZN(new_n1006));
  NAND2_X1  g581(.A1(G303), .A2(G8), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(KEYINPUT55), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1011), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n957), .A2(KEYINPUT45), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n954), .B1(new_n492), .B2(new_n498), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n474), .A2(new_n958), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n705), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1015), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n996), .A2(new_n998), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n1022), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1020), .B1(new_n1026), .B2(G2090), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1013), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1001), .B1(new_n1003), .B2(G288), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  OR2_X1    g605(.A1(new_n1030), .A2(KEYINPUT120), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(G288), .A2(new_n1030), .A3(new_n1003), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(new_n1002), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1028), .A3(new_n1002), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n996), .A2(KEYINPUT50), .A3(new_n998), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n959), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1020), .B1(new_n1041), .B2(G2090), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1013), .B1(G8), .B2(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1037), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT50), .B1(new_n996), .B2(new_n998), .ZN(new_n1045));
  NOR3_X1   g620(.A1(new_n1045), .A2(new_n1023), .A3(G2084), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n996), .A2(new_n1016), .A3(new_n998), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1048), .A2(KEYINPUT121), .A3(new_n1018), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT121), .B1(new_n1048), .B2(new_n1018), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1047), .B1(new_n1052), .B2(G1966), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G286), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT63), .B1(new_n1044), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1027), .A2(G8), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT63), .B1(new_n1057), .B2(new_n1013), .ZN(new_n1058));
  NOR4_X1   g633(.A1(new_n1037), .A2(new_n1058), .A3(G286), .A4(new_n1054), .ZN(new_n1059));
  OAI221_X1 g634(.A(new_n1006), .B1(new_n1028), .B2(new_n1036), .C1(new_n1056), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g636(.A1(G286), .A2(G8), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n1062), .B(KEYINPUT124), .Z(new_n1063));
  NAND3_X1  g638(.A1(new_n1054), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n1063), .B(KEYINPUT125), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1053), .A2(KEYINPUT123), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n853), .A2(new_n997), .A3(new_n954), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n997), .B1(new_n853), .B2(new_n954), .ZN(new_n1069));
  NOR3_X1   g644(.A1(new_n1068), .A2(new_n1069), .A3(KEYINPUT45), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1070), .B2(new_n959), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1051), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1048), .A2(KEYINPUT121), .A3(new_n1018), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n1077), .A3(new_n1047), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1066), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1065), .B1(new_n1079), .B2(G8), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1063), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1077), .B1(new_n1076), .B2(new_n1047), .ZN(new_n1082));
  AOI211_X1 g657(.A(KEYINPUT123), .B(new_n1046), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT51), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1064), .B1(new_n1080), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2078), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1052), .A2(KEYINPUT53), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1019), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT53), .B1(new_n1089), .B2(new_n1087), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1090), .B1(new_n767), .B2(new_n1026), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G301), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1086), .A2(KEYINPUT62), .A3(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n999), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1025), .A2(G1348), .B1(new_n1095), .B2(G2067), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n598), .B(KEYINPUT122), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n598), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1096), .A2(new_n1097), .B1(KEYINPUT122), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1100), .B1(new_n1102), .B2(new_n1098), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G299), .B(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT56), .B(G2072), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1014), .A2(new_n1017), .A3(new_n1018), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(G1956), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1104), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1104), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n1106), .C1(new_n1040), .C2(G1956), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1111), .A3(KEYINPUT61), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  AOI22_X1  g689(.A1(new_n1089), .A2(new_n964), .B1(new_n1095), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1113), .B1(new_n1115), .B2(new_n551), .ZN(new_n1116));
  AND2_X1   g691(.A1(new_n1112), .A2(new_n1116), .ZN(new_n1117));
  OR3_X1    g692(.A1(new_n1115), .A2(new_n1113), .A3(new_n551), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1103), .A2(new_n1117), .A3(new_n1118), .A4(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1111), .A2(new_n1096), .A3(new_n598), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(new_n1123), .A3(new_n1109), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1125), .B1(new_n1016), .B2(new_n956), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(KEYINPUT53), .A3(new_n1087), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1091), .A2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g703(.A(G171), .B(KEYINPUT54), .Z(new_n1129));
  MUX2_X1   g704(.A(new_n1128), .B(new_n1092), .S(new_n1129), .Z(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1124), .A2(new_n1130), .B1(new_n1131), .B2(new_n1093), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1094), .B1(new_n1132), .B2(new_n1086), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1060), .B1(new_n1133), .B2(new_n1044), .ZN(new_n1134));
  XOR2_X1   g709(.A(G290), .B(G1986), .Z(new_n1135));
  OAI21_X1  g710(.A(new_n976), .B1(new_n1135), .B2(new_n966), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n990), .B1(new_n1134), .B2(new_n1136), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g712(.A1(new_n663), .A2(new_n664), .A3(new_n643), .ZN(new_n1139));
  AOI21_X1  g713(.A(new_n1139), .B1(new_n869), .B2(new_n871), .ZN(new_n1140));
  NAND4_X1  g714(.A1(new_n1140), .A2(new_n947), .A3(new_n456), .A4(new_n688), .ZN(G225));
  INV_X1    g715(.A(G225), .ZN(G308));
endmodule


