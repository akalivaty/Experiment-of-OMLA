//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:01 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT65), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  OR4_X1    g028(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT70), .Z(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G101), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(new_n458), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n464), .A2(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n465), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OR3_X1    g050(.A1(new_n475), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(KEYINPUT71), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n475), .A2(new_n465), .ZN(new_n480));
  MUX2_X1   g055(.A(G100), .B(G112), .S(G2105), .Z(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G124), .B1(G2104), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(G126), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n485), .B1(new_n462), .B2(new_n463), .ZN(new_n486));
  AND2_X1   g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  OAI21_X1  g062(.A(G2105), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT4), .A2(G138), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(new_n462), .B2(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n465), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  OAI211_X1 g068(.A(G138), .B(new_n465), .C1(new_n473), .C2(new_n474), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n488), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  NOR2_X1   g073(.A1(KEYINPUT6), .A2(G651), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT72), .B(G651), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT6), .ZN(new_n501));
  XOR2_X1   g076(.A(KEYINPUT5), .B(G543), .Z(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G88), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G50), .ZN(new_n507));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(new_n500), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n504), .A2(new_n507), .A3(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT72), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT72), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI211_X1 g092(.A(G51), .B(G543), .C1(new_n517), .C2(new_n499), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND2_X1  g095(.A1(G63), .A2(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT73), .B1(new_n502), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n523), .A2(new_n524), .A3(G63), .A4(G651), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n518), .A2(new_n520), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n503), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(G168));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n502), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT74), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(KEYINPUT74), .B(new_n531), .C1(new_n502), .C2(new_n532), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(new_n500), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n503), .A2(G90), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT75), .B(G52), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n506), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n502), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n503), .A2(G81), .B1(new_n545), .B2(new_n500), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n506), .A2(G43), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(KEYINPUT76), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n506), .A2(KEYINPUT9), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n503), .A2(KEYINPUT77), .A3(G91), .ZN(new_n558));
  OAI211_X1 g133(.A(G91), .B(new_n523), .C1(new_n517), .C2(new_n499), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n523), .A2(G65), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n564), .A2(KEYINPUT78), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n563), .A2(KEYINPUT79), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT79), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n506), .A2(new_n556), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n568), .A2(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n562), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(new_n528), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT80), .B1(new_n576), .B2(new_n526), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n527), .A2(new_n578), .A3(new_n528), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G286));
  NAND2_X1  g156(.A1(new_n503), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n506), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  OAI211_X1 g160(.A(G86), .B(new_n523), .C1(new_n517), .C2(new_n499), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT83), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n523), .A2(G61), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n523), .A2(KEYINPUT81), .A3(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT82), .Z(new_n593));
  NAND3_X1  g168(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(new_n500), .B1(new_n506), .B2(G48), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n587), .A2(new_n595), .A3(KEYINPUT84), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(KEYINPUT84), .B1(new_n587), .B2(new_n595), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n597), .A2(new_n598), .ZN(G305));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G60), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n502), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n503), .A2(G85), .B1(new_n500), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(new_n506), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n502), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G651), .ZN(new_n610));
  INV_X1    g185(.A(G54), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n503), .A2(G92), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n503), .A2(KEYINPUT10), .A3(G92), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G868), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n618), .B2(G301), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT85), .ZN(G284));
  INV_X1    g196(.A(new_n620), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n618), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n580), .B2(new_n618), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n580), .B2(new_n618), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n617), .B1(new_n626), .B2(G860), .ZN(G148));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n617), .A2(new_n628), .A3(new_n626), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n628), .B1(new_n617), .B2(new_n626), .ZN(new_n631));
  OAI21_X1  g206(.A(G868), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g209(.A1(new_n475), .A2(G2105), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G2104), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  INV_X1    g214(.A(G2100), .ZN(new_n640));
  OR2_X1    g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n480), .A2(G123), .ZN(new_n643));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  OR3_X1    g222(.A1(new_n465), .A2(KEYINPUT87), .A3(G111), .ZN(new_n648));
  OAI21_X1  g223(.A(KEYINPUT87), .B1(new_n465), .B2(G111), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n646), .A2(new_n647), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n476), .A2(new_n477), .ZN(new_n651));
  INV_X1    g226(.A(G135), .ZN(new_n652));
  OAI211_X1 g227(.A(new_n643), .B(new_n650), .C1(new_n651), .C2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(G2096), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n641), .A2(new_n642), .A3(new_n655), .ZN(G156));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT15), .B(G2435), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2427), .ZN(new_n660));
  INV_X1    g235(.A(G2430), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n657), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2443), .B(G2446), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1341), .B(G1348), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n663), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G401));
  XNOR2_X1  g248(.A(G2072), .B(G2078), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT89), .ZN(new_n676));
  XOR2_X1   g251(.A(G2084), .B(G2090), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n674), .B1(new_n679), .B2(KEYINPUT17), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(KEYINPUT17), .A3(new_n674), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n677), .B1(KEYINPUT17), .B2(new_n674), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n676), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n675), .B(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n674), .A3(new_n677), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(new_n654), .A3(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n654), .B1(new_n684), .B2(new_n689), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n640), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n692), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n694), .A2(G2100), .A3(new_n690), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(G227));
  XOR2_X1   g271(.A(G1971), .B(G1976), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT19), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1956), .B(G2474), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1961), .B(G1966), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n698), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n698), .A2(new_n701), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT20), .Z(new_n705));
  AOI211_X1 g280(.A(new_n703), .B(new_n705), .C1(new_n698), .C2(new_n702), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1981), .B(G1986), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT90), .ZN(new_n710));
  XOR2_X1   g285(.A(G1991), .B(G1996), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n708), .B(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(G229));
  NAND3_X1  g289(.A1(new_n478), .A2(KEYINPUT92), .A3(G139), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT92), .ZN(new_n716));
  INV_X1    g291(.A(G139), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n651), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n459), .A2(G103), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  NAND3_X1  g295(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n721), .A2(KEYINPUT93), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT93), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n715), .A2(new_n723), .A3(new_n718), .A4(new_n720), .ZN(new_n724));
  AOI22_X1  g299(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n465), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT94), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(G29), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G33), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(G29), .B2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(G2072), .Z(new_n732));
  INV_X1    g307(.A(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G35), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT101), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n483), .B2(G29), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT29), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  AND3_X1   g315(.A1(new_n739), .A2(G2090), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(G2090), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g318(.A1(KEYINPUT24), .A2(G34), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT24), .A2(G34), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n733), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT95), .Z(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G160), .B2(G29), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G2084), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT99), .Z(new_n750));
  INV_X1    g325(.A(G16), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n751), .A2(G5), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G301), .B2(G16), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(G164), .A2(G29), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G27), .B2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT100), .B(G2078), .Z(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n757), .A2(new_n759), .B1(G2084), .B2(new_n748), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n750), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n733), .A2(G26), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT28), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n478), .A2(G140), .ZN(new_n765));
  MUX2_X1   g340(.A(G104), .B(G116), .S(G2105), .Z(new_n766));
  AOI22_X1  g341(.A1(new_n480), .A2(G128), .B1(G2104), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n764), .B1(new_n768), .B2(G29), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT91), .B(G2067), .Z(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n757), .A2(new_n759), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n733), .A2(G32), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n478), .A2(G141), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n459), .A2(G105), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT26), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n777), .B(new_n779), .C1(G129), .C2(new_n480), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n775), .B1(new_n782), .B2(new_n733), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT27), .B(G1996), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n783), .A2(new_n785), .B1(new_n769), .B2(new_n771), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n548), .A2(G16), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G16), .B2(G19), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n788), .A2(G1341), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(G1341), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n774), .B(new_n786), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n743), .A2(new_n761), .A3(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n775), .B(new_n784), .C1(new_n782), .C2(new_n733), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT96), .Z(new_n794));
  NOR2_X1   g369(.A1(G4), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(new_n617), .B2(G16), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1348), .Z(new_n797));
  XOR2_X1   g372(.A(KEYINPUT31), .B(G11), .Z(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(KEYINPUT30), .A2(G28), .ZN(new_n800));
  NOR2_X1   g375(.A1(KEYINPUT30), .A2(G28), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n799), .A2(KEYINPUT97), .B1(new_n733), .B2(new_n802), .ZN(new_n803));
  OAI221_X1 g378(.A(new_n803), .B1(KEYINPUT97), .B2(new_n799), .C1(new_n653), .C2(new_n733), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n751), .A2(G21), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n529), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n753), .A2(new_n754), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  AND3_X1   g387(.A1(new_n794), .A2(new_n797), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n751), .A2(G20), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT23), .Z(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G299), .B2(G16), .ZN(new_n816));
  INV_X1    g391(.A(G1956), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n808), .A2(new_n809), .A3(new_n810), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(KEYINPUT98), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n732), .A2(new_n792), .A3(new_n813), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(G16), .B1(new_n597), .B2(new_n598), .ZN(new_n822));
  NOR2_X1   g397(.A1(G6), .A2(G16), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT32), .B(G1981), .Z(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT34), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n751), .A2(G23), .ZN(new_n830));
  INV_X1    g405(.A(G288), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n751), .ZN(new_n832));
  XOR2_X1   g407(.A(KEYINPUT33), .B(G1976), .Z(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(G16), .A2(G22), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(G166), .B2(G16), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1971), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n828), .A2(new_n829), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(G16), .A2(G24), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(G290), .B2(new_n751), .ZN(new_n841));
  INV_X1    g416(.A(G1986), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n478), .A2(G131), .ZN(new_n845));
  MUX2_X1   g420(.A(G95), .B(G107), .S(G2105), .Z(new_n846));
  AOI22_X1  g421(.A1(new_n480), .A2(G119), .B1(G2104), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G29), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G25), .B2(G29), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT35), .B(G1991), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n853), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n843), .B(new_n844), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n839), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n829), .B1(new_n828), .B2(new_n838), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT36), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n828), .A2(new_n838), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT34), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT36), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n839), .A4(new_n857), .ZN(new_n864));
  AOI211_X1 g439(.A(KEYINPUT102), .B(new_n821), .C1(new_n860), .C2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT102), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n860), .A2(new_n864), .ZN(new_n867));
  INV_X1    g442(.A(new_n821), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n865), .A2(new_n869), .ZN(G311));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n868), .ZN(G150));
  XNOR2_X1  g446(.A(KEYINPUT103), .B(G860), .ZN(new_n872));
  NAND2_X1  g447(.A1(G80), .A2(G543), .ZN(new_n873));
  INV_X1    g448(.A(G67), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n502), .B2(new_n874), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n503), .A2(G93), .B1(new_n875), .B2(new_n500), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n506), .A2(G55), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n872), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n546), .A2(new_n547), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n546), .A2(new_n876), .A3(new_n547), .A4(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT38), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n617), .A2(G559), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n872), .B1(new_n888), .B2(KEYINPUT39), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(G145));
  OAI21_X1  g466(.A(new_n781), .B1(new_n722), .B2(new_n728), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n721), .A2(KEYINPUT93), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(new_n724), .A3(new_n727), .A4(new_n782), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n480), .A2(G130), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n478), .A2(G142), .ZN(new_n897));
  OR3_X1    g472(.A1(new_n465), .A2(KEYINPUT106), .A3(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(KEYINPUT106), .B1(new_n465), .B2(G118), .ZN(new_n899));
  OR2_X1    g474(.A1(G106), .A2(G2105), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n898), .A2(G2104), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n638), .A2(new_n845), .A3(new_n847), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n638), .B1(new_n845), .B2(new_n847), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n638), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n848), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n902), .A3(new_n904), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n497), .A2(KEYINPUT104), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n488), .A2(new_n493), .A3(new_n912), .A4(new_n496), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n765), .A3(new_n767), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n768), .A2(new_n911), .A3(new_n913), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n907), .A2(new_n910), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n907), .A2(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n892), .B(new_n894), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n892), .A2(new_n894), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n917), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(KEYINPUT107), .A3(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(new_n483), .B(G160), .Z(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(new_n653), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G37), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n920), .A2(new_n929), .A3(KEYINPUT107), .A4(new_n923), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g507(.A1(new_n881), .A2(G868), .ZN(new_n933));
  XNOR2_X1  g508(.A(G290), .B(G288), .ZN(new_n934));
  INV_X1    g509(.A(new_n598), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n935), .A2(G166), .A3(new_n596), .ZN(new_n936));
  OAI21_X1  g511(.A(G303), .B1(new_n597), .B2(new_n598), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n936), .A2(new_n937), .A3(new_n934), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT109), .B1(new_n943), .B2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n943), .A2(new_n938), .A3(KEYINPUT42), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n884), .ZN(new_n949));
  NOR3_X1   g524(.A1(new_n630), .A2(new_n631), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n617), .A2(new_n626), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT86), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n884), .B1(new_n952), .B2(new_n629), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g529(.A1(new_n506), .A2(G54), .B1(new_n609), .B2(G651), .ZN(new_n955));
  INV_X1    g530(.A(new_n616), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT10), .B1(new_n503), .B2(G92), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n955), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g533(.A1(G299), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n615), .A2(new_n616), .ZN(new_n960));
  AOI22_X1  g535(.A1(new_n574), .A2(new_n562), .B1(new_n960), .B2(new_n955), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n954), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  INV_X1    g540(.A(new_n953), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n952), .A2(new_n629), .A3(new_n884), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n962), .A4(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT41), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n959), .A2(new_n961), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n617), .A2(new_n574), .A3(new_n562), .ZN(new_n972));
  NAND2_X1  g547(.A1(G299), .A2(new_n958), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT41), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n975), .B1(new_n950), .B2(new_n953), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n964), .A2(new_n965), .A3(new_n969), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n969), .A2(new_n976), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n967), .B1(new_n954), .B2(new_n962), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n948), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n977), .B(new_n980), .C1(new_n946), .C2(new_n947), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n933), .B1(new_n984), .B2(G868), .ZN(G295));
  AOI21_X1  g560(.A(new_n933), .B1(new_n984), .B2(G868), .ZN(G331));
  NAND3_X1  g561(.A1(G171), .A2(new_n577), .A3(new_n579), .ZN(new_n987));
  NAND2_X1  g562(.A1(G168), .A2(G301), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(KEYINPUT112), .A3(new_n949), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n987), .A2(new_n884), .A3(new_n988), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n884), .B1(new_n988), .B2(new_n987), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n989), .A2(new_n949), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(new_n991), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n995), .A2(new_n962), .B1(new_n975), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n945), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(KEYINPUT113), .B(new_n928), .C1(new_n945), .C2(new_n998), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n962), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n996), .A2(new_n992), .A3(new_n991), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n990), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n970), .B1(new_n959), .B2(new_n961), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n972), .A2(new_n973), .A3(KEYINPUT41), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n987), .A2(new_n884), .A3(new_n988), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n1005), .B(new_n1006), .C1(new_n1007), .C2(new_n994), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n944), .B(new_n942), .C1(new_n1004), .C2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT113), .B1(new_n1010), .B2(new_n928), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT43), .B(new_n999), .C1(new_n1001), .C2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1013));
  OAI22_X1  g588(.A1(new_n995), .A2(new_n1013), .B1(new_n1002), .B2(new_n997), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n944), .A3(new_n942), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n999), .A2(new_n1015), .A3(new_n928), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n1019));
  NAND3_X1  g594(.A1(new_n1012), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n1017), .B(new_n999), .C1(new_n1001), .C2(new_n1011), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n1016), .B2(KEYINPUT43), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1020), .A2(new_n1024), .ZN(G397));
  INV_X1    g600(.A(KEYINPUT124), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(G166), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1384), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n497), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT50), .ZN(new_n1034));
  INV_X1    g609(.A(G40), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n468), .A2(new_n471), .A3(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT115), .B(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n497), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1034), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G2090), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT45), .B1(new_n497), .B2(new_n1032), .ZN(new_n1041));
  INV_X1    g616(.A(G125), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n475), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n470), .ZN(new_n1044));
  OAI21_X1  g619(.A(G2105), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n635), .A2(G137), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1045), .A2(G40), .A3(new_n460), .A4(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1041), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n911), .A2(KEYINPUT45), .A3(new_n1032), .A4(new_n913), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1971), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1031), .B(G8), .C1(new_n1040), .C2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1033), .A2(new_n1047), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(new_n1028), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n582), .A2(new_n583), .A3(G1976), .A4(new_n584), .ZN(new_n1054));
  INV_X1    g629(.A(G1976), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT52), .B1(G288), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n489), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1058), .B1(new_n473), .B2(new_n474), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n491), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1060), .A2(new_n465), .B1(new_n495), .B2(new_n494), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1384), .B1(new_n1061), .B2(new_n488), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1036), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1063), .A2(G8), .A3(new_n1054), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT49), .ZN(new_n1067));
  INV_X1    g642(.A(G1981), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n587), .A2(new_n595), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n595), .B2(new_n586), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n595), .A2(new_n586), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G1981), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n587), .A2(new_n595), .A3(new_n1068), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1073), .A2(KEYINPUT49), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1071), .A2(new_n1075), .A3(new_n1053), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1051), .A2(new_n1066), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1062), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1081), .B(new_n1036), .C1(new_n1062), .C2(new_n1037), .ZN(new_n1082));
  OAI22_X1  g657(.A1(new_n1079), .A2(G1971), .B1(new_n1082), .B2(G2090), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1031), .B1(new_n1083), .B2(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1026), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1053), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1087), .B1(new_n1088), .B2(new_n1067), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1086), .B1(new_n1089), .B2(new_n1075), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1082), .A2(G2090), .ZN(new_n1091));
  OAI21_X1  g666(.A(G8), .B1(new_n1091), .B2(new_n1050), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1031), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1090), .A2(new_n1094), .A3(KEYINPUT124), .A4(new_n1051), .ZN(new_n1095));
  INV_X1    g670(.A(G2078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1048), .A2(new_n1049), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1097), .A2(new_n1098), .B1(new_n754), .B2(new_n1039), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1036), .B(KEYINPUT118), .C1(new_n1062), .C2(KEYINPUT45), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT119), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1062), .B2(KEYINPUT45), .ZN(new_n1105));
  AND4_X1   g680(.A1(new_n1104), .A2(new_n497), .A3(KEYINPUT45), .A4(new_n1032), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1096), .A2(KEYINPUT53), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1099), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  AND4_X1   g685(.A1(G171), .A2(new_n1085), .A3(new_n1095), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(G1966), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1039), .B2(G2084), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1047), .B1(new_n1062), .B2(new_n1037), .ZN(new_n1115));
  INV_X1    g690(.A(G2084), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1115), .A2(KEYINPUT120), .A3(new_n1116), .A4(new_n1034), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(G8), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT51), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n529), .A2(G8), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n807), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(new_n1114), .A3(new_n1117), .ZN(new_n1126));
  OAI211_X1 g701(.A(KEYINPUT51), .B(G8), .C1(new_n1126), .C2(new_n529), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1122), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1118), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1121), .B1(new_n1129), .B2(new_n1125), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT62), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1133), .B(new_n1130), .C1(new_n1122), .C2(new_n1127), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1111), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(G1348), .B1(new_n1115), .B2(new_n1034), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1063), .A2(G2067), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n617), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1036), .B1(new_n1033), .B2(KEYINPUT50), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1062), .A2(new_n1037), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n817), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT56), .B(G2072), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1048), .A2(new_n1049), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT57), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n562), .A2(new_n574), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n572), .A2(new_n573), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n571), .A2(G651), .A3(new_n567), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n557), .A2(new_n558), .A3(new_n561), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT57), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1142), .A2(new_n1144), .A3(new_n1146), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1151), .A2(new_n1146), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g731(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1156), .A2(new_n1152), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g736(.A(KEYINPUT122), .B(KEYINPUT61), .C1(new_n1156), .C2(new_n1152), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT58), .B(G1341), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1078), .A2(G1996), .B1(new_n1052), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n548), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(new_n548), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n958), .A2(KEYINPUT60), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1171), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1172));
  INV_X1    g747(.A(G2067), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1052), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1062), .A2(new_n1080), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1038), .A2(new_n1036), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g752(.A(new_n958), .B(new_n1174), .C1(new_n1177), .C2(G1348), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1138), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1172), .B1(new_n1179), .B2(KEYINPUT60), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1156), .A2(KEYINPUT61), .A3(new_n1152), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1170), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1157), .B1(new_n1163), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1184));
  NOR2_X1   g759(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT54), .ZN(new_n1186));
  NOR2_X1   g761(.A1(G301), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1188), .ZN(new_n1189));
  AND2_X1   g764(.A1(new_n1189), .A2(new_n1099), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1049), .A2(KEYINPUT53), .A3(new_n1096), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n911), .A2(new_n1032), .A3(new_n913), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT45), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1047), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1191), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1196), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1197));
  AOI22_X1  g772(.A1(new_n1190), .A2(new_n1197), .B1(new_n1110), .B2(new_n1188), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1085), .A2(new_n1198), .A3(new_n1095), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1183), .A2(new_n1184), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT121), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1119), .B2(G286), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1126), .A2(KEYINPUT121), .A3(G8), .A4(new_n580), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(G8), .B1(new_n1040), .B2(new_n1050), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1093), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1206), .A2(KEYINPUT63), .A3(new_n1051), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1066), .A2(new_n1076), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1208), .A2(KEYINPUT116), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT116), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1066), .A2(new_n1076), .A3(new_n1210), .ZN(new_n1211));
  AOI21_X1  g786(.A(new_n1207), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1204), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1090), .A2(new_n1094), .A3(new_n1051), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n1214), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1213), .B1(KEYINPUT63), .B2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1076), .A2(new_n1055), .A3(new_n831), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1087), .B1(new_n1217), .B2(new_n1074), .ZN(new_n1218));
  INV_X1    g793(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1211), .ZN(new_n1220));
  AOI21_X1  g795(.A(new_n1210), .B1(new_n1066), .B2(new_n1076), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1219), .B(KEYINPUT117), .C1(new_n1222), .C2(new_n1051), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT117), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1051), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1224), .B1(new_n1225), .B2(new_n1218), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  NAND4_X1  g802(.A1(new_n1135), .A2(new_n1200), .A3(new_n1216), .A4(new_n1227), .ZN(new_n1228));
  AND3_X1   g803(.A1(new_n1193), .A2(new_n1194), .A3(new_n1036), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n768), .B(G2067), .ZN(new_n1230));
  XNOR2_X1  g805(.A(new_n1230), .B(KEYINPUT114), .ZN(new_n1231));
  INV_X1    g806(.A(G1996), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n781), .B(new_n1232), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n848), .A2(new_n853), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n849), .A2(new_n852), .ZN(new_n1235));
  NAND4_X1  g810(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .A4(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g811(.A(G290), .B(G1986), .ZN(new_n1237));
  OAI21_X1  g812(.A(new_n1229), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g813(.A1(new_n1228), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1231), .A2(new_n782), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1229), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1242));
  XNOR2_X1  g817(.A(new_n1242), .B(KEYINPUT46), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  XOR2_X1   g819(.A(new_n1244), .B(KEYINPUT47), .Z(new_n1245));
  NAND2_X1  g820(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1246));
  OAI22_X1  g821(.A1(new_n1246), .A2(new_n1235), .B1(G2067), .B2(new_n768), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1247), .A2(new_n1229), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1236), .A2(new_n1229), .ZN(new_n1249));
  NOR2_X1   g824(.A1(G290), .A2(G1986), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1229), .A2(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g826(.A(new_n1251), .B(KEYINPUT125), .ZN(new_n1252));
  INV_X1    g827(.A(KEYINPUT48), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1249), .A2(new_n1254), .ZN(new_n1255));
  NOR2_X1   g830(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1256));
  OAI21_X1  g831(.A(new_n1248), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g832(.A1(new_n1245), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g833(.A1(new_n1239), .A2(new_n1258), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g834(.A1(new_n693), .A2(new_n695), .A3(G319), .ZN(new_n1261));
  INV_X1    g835(.A(KEYINPUT126), .ZN(new_n1262));
  NAND2_X1  g836(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND4_X1  g837(.A1(new_n693), .A2(new_n695), .A3(KEYINPUT126), .A4(G319), .ZN(new_n1264));
  NAND3_X1  g838(.A1(new_n1263), .A2(new_n672), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g839(.A1(new_n1265), .A2(KEYINPUT127), .ZN(new_n1266));
  INV_X1    g840(.A(KEYINPUT127), .ZN(new_n1267));
  NAND4_X1  g841(.A1(new_n1263), .A2(new_n1267), .A3(new_n672), .A4(new_n1264), .ZN(new_n1268));
  NAND2_X1  g842(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AND3_X1   g843(.A1(new_n931), .A2(new_n1269), .A3(new_n713), .ZN(new_n1270));
  AND3_X1   g844(.A1(new_n1270), .A2(new_n1018), .A3(new_n1012), .ZN(G308));
  NAND3_X1  g845(.A1(new_n1270), .A2(new_n1018), .A3(new_n1012), .ZN(G225));
endmodule


