//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1304, new_n1305, new_n1306, new_n1307, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(G77), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT69), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n212), .A2(new_n213), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n209), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT70), .ZN(new_n220));
  INV_X1    g0020(.A(KEYINPUT1), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT71), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n209), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  INV_X1    g0026(.A(G50), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT66), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n227), .B1(new_n202), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n228), .B2(new_n202), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT67), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT68), .Z(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n226), .B1(new_n221), .B2(new_n220), .C1(new_n232), .C2(new_n236), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n223), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT72), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  INV_X1    g0043(.A(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT2), .B(G226), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n242), .B(new_n247), .ZN(G358));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n233), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT74), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT75), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(G58), .ZN(new_n260));
  INV_X1    g0060(.A(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT74), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n260), .A2(KEYINPUT8), .A3(new_n262), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n261), .A2(KEYINPUT75), .A3(KEYINPUT8), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n234), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G150), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n234), .A2(new_n270), .ZN(new_n271));
  OAI22_X1  g0071(.A1(new_n203), .A2(new_n234), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n257), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  OR2_X1    g0073(.A1(KEYINPUT73), .A2(G1), .ZN(new_n274));
  NAND2_X1  g0074(.A1(KEYINPUT73), .A2(G1), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(G13), .A3(G20), .A4(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n227), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n275), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(new_n234), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT76), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT76), .B1(new_n280), .B2(new_n234), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n257), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n285), .A2(new_n227), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n270), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  AOI21_X1  g0093(.A(G1698), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G222), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT3), .B(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G223), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(G1698), .ZN(new_n298));
  OAI221_X1 g0098(.A(new_n295), .B1(new_n204), .B2(new_n296), .C1(new_n297), .C2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  INV_X1    g0102(.A(new_n233), .ZN(new_n303));
  NAND2_X1  g0103(.A1(G33), .A2(G41), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G41), .ZN(new_n306));
  INV_X1    g0106(.A(G45), .ZN(new_n307));
  AOI21_X1  g0107(.A(G1), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(KEYINPUT73), .A2(G1), .ZN(new_n310));
  NOR2_X1   g0110(.A1(KEYINPUT73), .A2(G1), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(G41), .A2(G45), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n300), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G226), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n301), .A2(new_n309), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n290), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n318), .A2(G190), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT78), .B(G200), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n289), .A2(KEYINPUT9), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT9), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(new_n279), .B2(new_n288), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n333), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n331), .A2(new_n333), .A3(new_n328), .A4(new_n325), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT10), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n324), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(G1698), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n296), .A2(G232), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G107), .ZN(new_n340));
  INV_X1    g0140(.A(G238), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n339), .B1(new_n340), .B2(new_n296), .C1(new_n298), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n300), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n304), .A2(G1), .A3(G13), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n308), .A2(new_n345), .A3(G274), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n315), .B2(G244), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n344), .B1(new_n343), .B2(new_n347), .ZN(new_n350));
  OAI21_X1  g0150(.A(G190), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n350), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n352), .A2(new_n327), .A3(new_n348), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n285), .A2(new_n204), .A3(new_n287), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT8), .B(G58), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n271), .B1(new_n234), .B2(new_n204), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n267), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n257), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G77), .B2(new_n276), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n354), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n351), .A2(new_n353), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n319), .B1(new_n349), .B2(new_n350), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n352), .A2(new_n321), .A3(new_n348), .ZN(new_n364));
  INV_X1    g0164(.A(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n337), .A2(new_n362), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT14), .ZN(new_n368));
  OAI211_X1 g0168(.A(G238), .B(new_n345), .C1(new_n280), .C2(new_n313), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G97), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(G226), .A2(G1698), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n244), .B2(G1698), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n371), .B1(new_n373), .B2(new_n296), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n309), .B(new_n369), .C1(new_n374), .C2(new_n345), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  INV_X1    g0176(.A(G226), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n338), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n244), .A2(G1698), .ZN(new_n379));
  AND2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n300), .B1(new_n383), .B2(new_n371), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n384), .A2(new_n385), .A3(new_n309), .A4(new_n369), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n376), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n368), .B1(new_n387), .B2(G169), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT79), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n375), .A2(KEYINPUT79), .A3(KEYINPUT13), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n391), .A2(G179), .A3(new_n386), .A4(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n387), .A2(new_n368), .A3(G169), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n234), .A2(G33), .A3(G77), .ZN(new_n396));
  INV_X1    g0196(.A(G68), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(G20), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n396), .B(new_n398), .C1(new_n271), .C2(new_n227), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n257), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT11), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT11), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n402), .A3(new_n257), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT12), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n277), .A2(new_n405), .A3(new_n397), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT12), .B1(new_n276), .B2(G68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n287), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n404), .B(new_n408), .C1(new_n285), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n395), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n387), .B2(G200), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n391), .A2(G190), .A3(new_n386), .A4(new_n392), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT80), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n409), .A2(new_n265), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n418), .A2(new_n285), .B1(new_n276), .B2(new_n265), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  INV_X1    g0220(.A(G159), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n271), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT74), .B(G58), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n202), .B1(new_n423), .B2(new_n397), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n422), .B1(new_n424), .B2(G20), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT7), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n296), .B2(G20), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n380), .A2(new_n381), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT7), .A3(new_n234), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n397), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT81), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n425), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT7), .B1(new_n428), .B2(new_n234), .ZN(new_n433));
  NOR4_X1   g0233(.A1(new_n380), .A2(new_n381), .A3(new_n426), .A4(G20), .ZN(new_n434));
  OAI21_X1  g0234(.A(G68), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n420), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n422), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n258), .A2(G58), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n262), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n201), .B1(new_n440), .B2(G68), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n438), .B1(new_n441), .B2(new_n234), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n442), .A2(new_n430), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n286), .B1(new_n443), .B2(KEYINPUT16), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n419), .B1(new_n437), .B2(new_n444), .ZN(new_n445));
  OAI211_X1 g0245(.A(G232), .B(new_n345), .C1(new_n280), .C2(new_n313), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n309), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n297), .A2(new_n338), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n377), .A2(G1698), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n448), .B(new_n449), .C1(new_n380), .C2(new_n381), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G87), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n345), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n321), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(new_n300), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(new_n319), .A3(new_n446), .A4(new_n309), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT82), .ZN(new_n457));
  AND3_X1   g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n453), .B2(new_n456), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT18), .B1(new_n445), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n419), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n346), .B1(new_n315), .B2(G232), .ZN(new_n463));
  INV_X1    g0263(.A(G190), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n455), .ZN(new_n465));
  INV_X1    g0265(.A(G200), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n466), .B1(new_n447), .B2(new_n452), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n442), .B1(KEYINPUT81), .B2(new_n435), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n430), .A2(new_n431), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT16), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n435), .A2(new_n425), .A3(KEYINPUT16), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n257), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n462), .B(new_n468), .C1(new_n471), .C2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT17), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(G169), .B1(new_n463), .B2(new_n455), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n447), .A2(G179), .A3(new_n452), .ZN(new_n478));
  OAI21_X1  g0278(.A(KEYINPUT82), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT18), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(new_n470), .A3(new_n425), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n473), .B1(new_n420), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n481), .B(new_n482), .C1(new_n485), .C2(new_n419), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n468), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n461), .A2(new_n476), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n367), .A2(new_n417), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n296), .A2(G264), .A3(G1698), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n296), .A2(G257), .A3(new_n338), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n428), .A2(G303), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n300), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT84), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(new_n306), .A3(KEYINPUT5), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT5), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n499), .B1(KEYINPUT84), .B2(G41), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NOR3_X1   g0302(.A1(new_n310), .A2(new_n311), .A3(new_n307), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n305), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n503), .A2(new_n498), .A3(new_n500), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(G270), .A3(new_n345), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n496), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G200), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n312), .A2(G33), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(new_n286), .A3(G116), .A4(new_n276), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n277), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n256), .A2(new_n233), .B1(G20), .B2(new_n511), .ZN(new_n514));
  AOI21_X1  g0314(.A(G20), .B1(G33), .B2(G283), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n270), .A2(G97), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT86), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT86), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT20), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT20), .B(new_n514), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n513), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n508), .B(new_n523), .C1(new_n464), .C2(new_n507), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT21), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n507), .A2(G169), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(new_n523), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n496), .A2(G179), .A3(new_n504), .A4(new_n506), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n522), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(new_n510), .A3(new_n512), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n531), .A2(KEYINPUT21), .A3(G169), .A4(new_n507), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n524), .A2(new_n527), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n271), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G77), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT6), .ZN(new_n537));
  INV_X1    g0337(.A(G97), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n537), .A2(new_n538), .A3(G107), .ZN(new_n539));
  XNOR2_X1  g0339(.A(G97), .B(G107), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n539), .B1(new_n537), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n536), .B1(new_n541), .B2(new_n234), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n340), .B1(new_n427), .B2(new_n429), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n257), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n509), .A2(new_n286), .A3(G97), .A4(new_n276), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n277), .A2(new_n538), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n274), .A2(G45), .A3(new_n275), .ZN(new_n549));
  OAI211_X1 g0349(.A(G257), .B(new_n345), .C1(new_n501), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n504), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(new_n338), .C1(new_n380), .C2(new_n381), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n296), .A2(KEYINPUT4), .A3(G244), .A4(new_n338), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G283), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n296), .A2(G250), .A3(G1698), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n551), .B1(new_n300), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(G190), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n300), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT83), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n563), .A3(new_n300), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n551), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n548), .B(new_n560), .C1(new_n565), .C2(new_n466), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n504), .A2(new_n550), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n561), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n568), .A2(new_n321), .B1(new_n544), .B2(new_n547), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n558), .A2(new_n563), .A3(new_n300), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n563), .B1(new_n558), .B2(new_n300), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n319), .B(new_n567), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n300), .B1(new_n502), .B2(new_n503), .ZN(new_n575));
  OAI211_X1 g0375(.A(G257), .B(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n576));
  OAI211_X1 g0376(.A(G250), .B(new_n338), .C1(new_n380), .C2(new_n381), .ZN(new_n577));
  INV_X1    g0377(.A(G294), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n577), .C1(new_n270), .C2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n575), .A2(G264), .B1(new_n579), .B2(new_n300), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n319), .A3(new_n504), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n300), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n505), .A2(G264), .A3(new_n345), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n504), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n321), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n234), .B(G87), .C1(new_n380), .C2(new_n381), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT87), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT22), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(KEYINPUT22), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n296), .A2(new_n234), .A3(G87), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT23), .B1(new_n234), .B2(G107), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT23), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n593), .A2(new_n340), .A3(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n234), .A2(G33), .A3(G116), .ZN(new_n595));
  NAND2_X1  g0395(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n592), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT88), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n602), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n591), .A2(new_n604), .A3(new_n598), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n286), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n276), .A2(G107), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n607), .A2(KEYINPUT25), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(KEYINPUT25), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n287), .B1(G33), .B2(new_n312), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(G107), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n581), .B(new_n585), .C1(new_n606), .C2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n604), .B1(new_n591), .B2(new_n598), .ZN(new_n614));
  AOI211_X1 g0414(.A(new_n602), .B(new_n597), .C1(new_n588), .C2(new_n590), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n257), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(G200), .B1(new_n580), .B2(new_n504), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n584), .A2(G190), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n616), .B(new_n611), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(G244), .B(G1698), .C1(new_n380), .C2(new_n381), .ZN(new_n620));
  OAI211_X1 g0420(.A(G238), .B(new_n338), .C1(new_n380), .C2(new_n381), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n620), .B(new_n621), .C1(new_n270), .C2(new_n511), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n300), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n503), .A2(new_n305), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n549), .A2(G250), .A3(new_n345), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n627), .A2(new_n464), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n270), .A2(new_n511), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n294), .B2(G238), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n345), .B1(new_n631), .B2(new_n620), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n624), .A2(new_n625), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n327), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT19), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n234), .B1(new_n370), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(G87), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n637), .A2(new_n538), .A3(new_n340), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n234), .B(G68), .C1(new_n380), .C2(new_n381), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n635), .B1(new_n267), .B2(new_n538), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n257), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n277), .A2(new_n357), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n509), .A2(new_n286), .A3(G87), .A4(new_n276), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n629), .A2(new_n634), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n633), .B1(new_n300), .B2(new_n622), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT85), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n319), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n623), .A2(new_n626), .A3(new_n319), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(KEYINPUT85), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n627), .A2(new_n321), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n409), .A2(new_n509), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n643), .B(new_n644), .C1(new_n654), .C2(new_n357), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n650), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n613), .A2(new_n619), .A3(new_n647), .A4(new_n656), .ZN(new_n657));
  NOR4_X1   g0457(.A1(new_n491), .A2(new_n534), .A3(new_n574), .A4(new_n657), .ZN(G372));
  AND2_X1   g0458(.A1(new_n461), .A2(new_n486), .ZN(new_n659));
  INV_X1    g0459(.A(new_n366), .ZN(new_n660));
  AOI22_X1  g0460(.A1(new_n660), .A2(new_n415), .B1(new_n411), .B2(new_n395), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n476), .A2(new_n487), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n659), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n334), .A2(new_n336), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n324), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n647), .A2(new_n656), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n667), .A2(new_n668), .A3(new_n573), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n653), .A2(new_n651), .A3(new_n655), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n634), .A2(new_n646), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n628), .B1(new_n671), .B2(KEYINPUT89), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n634), .A2(new_n646), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n670), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT90), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n573), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n569), .A2(new_n572), .A3(KEYINPUT90), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n669), .B1(new_n679), .B2(new_n668), .ZN(new_n680));
  INV_X1    g0480(.A(new_n670), .ZN(new_n681));
  INV_X1    g0481(.A(new_n613), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n527), .A2(new_n533), .A3(new_n532), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n326), .B1(new_n623), .B2(new_n626), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n686));
  OAI21_X1  g0486(.A(KEYINPUT89), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(new_n629), .A3(new_n674), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n566), .A2(new_n573), .A3(new_n619), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n681), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n680), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n666), .B1(new_n491), .B2(new_n692), .ZN(G369));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n234), .A2(G13), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT91), .B1(new_n280), .B2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT27), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT91), .ZN(new_n699));
  INV_X1    g0499(.A(new_n696), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n312), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n697), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G213), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n280), .A2(KEYINPUT91), .A3(new_n696), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n699), .B1(new_n312), .B2(new_n700), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT27), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(KEYINPUT92), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT92), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(KEYINPUT27), .C1(new_n704), .C2(new_n705), .ZN(new_n709));
  AOI211_X1 g0509(.A(new_n695), .B(new_n703), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n683), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n616), .A2(new_n611), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n710), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n613), .A2(new_n714), .A3(new_n619), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n713), .A2(new_n710), .A3(new_n581), .A4(new_n585), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT94), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n719), .A3(new_n716), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n712), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n613), .A2(new_n710), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n694), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n712), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n715), .A2(new_n719), .A3(new_n716), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n719), .B1(new_n715), .B2(new_n716), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n722), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n727), .A2(KEYINPUT95), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n718), .A2(new_n720), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  XOR2_X1   g0532(.A(KEYINPUT93), .B(G330), .Z(new_n733));
  NOR2_X1   g0533(.A1(new_n711), .A2(new_n523), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n534), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n683), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n733), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n732), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n730), .A2(new_n740), .ZN(G399));
  NOR2_X1   g0541(.A1(new_n638), .A2(G116), .ZN(new_n742));
  INV_X1    g0542(.A(new_n224), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n742), .B(G1), .C1(G41), .C2(new_n743), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT96), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n743), .A2(G41), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n745), .B1(new_n231), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT28), .Z(new_n748));
  AOI21_X1  g0548(.A(G179), .B1(new_n623), .B2(new_n626), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n749), .A2(new_n507), .A3(new_n584), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AND4_X1   g0552(.A1(new_n583), .A2(new_n582), .A3(new_n623), .A4(new_n626), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n529), .A2(new_n753), .A3(new_n559), .A4(KEYINPUT30), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n648), .A2(new_n580), .A3(new_n567), .A4(new_n561), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n756), .B2(new_n528), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n752), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  XOR2_X1   g0558(.A(KEYINPUT97), .B(KEYINPUT31), .Z(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n758), .A2(new_n710), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(KEYINPUT31), .B1(new_n758), .B2(new_n710), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AND4_X1   g0563(.A1(new_n613), .A2(new_n619), .A3(new_n647), .A4(new_n656), .ZN(new_n764));
  INV_X1    g0564(.A(new_n574), .ZN(new_n765));
  INV_X1    g0565(.A(new_n534), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n711), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n733), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT98), .ZN(new_n769));
  INV_X1    g0569(.A(new_n689), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n613), .A2(new_n527), .A3(new_n532), .A4(new_n533), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n670), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND4_X1  g0572(.A1(new_n675), .A2(new_n677), .A3(KEYINPUT26), .A4(new_n678), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n668), .B1(new_n667), .B2(new_n573), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n769), .B1(new_n776), .B2(new_n711), .ZN(new_n777));
  AOI211_X1 g0577(.A(KEYINPUT98), .B(new_n710), .C1(new_n772), .C2(new_n775), .ZN(new_n778));
  OAI21_X1  g0578(.A(KEYINPUT29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(KEYINPUT29), .B1(new_n691), .B2(new_n711), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n768), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n748), .B1(new_n782), .B2(G1), .ZN(G364));
  OAI21_X1  g0583(.A(G1), .B1(new_n696), .B2(new_n307), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n746), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT99), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n787), .A2(G13), .A3(G33), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n787), .B1(G13), .B2(G33), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G20), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n233), .B1(G20), .B2(new_n321), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  XOR2_X1   g0594(.A(new_n794), .B(KEYINPUT100), .Z(new_n795));
  XOR2_X1   g0595(.A(new_n795), .B(KEYINPUT101), .Z(new_n796));
  NOR2_X1   g0596(.A1(new_n743), .A2(new_n296), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n254), .B2(G45), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(new_n232), .B2(G45), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n743), .A2(new_n428), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n801), .A2(G355), .B1(new_n511), .B2(new_n743), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n796), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n234), .A2(new_n319), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n804), .A2(new_n464), .A3(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G317), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(KEYINPUT33), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n807), .A2(KEYINPUT33), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NOR3_X1   g0610(.A1(new_n464), .A2(G179), .A3(G200), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n234), .ZN(new_n812));
  INV_X1    g0612(.A(G326), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n804), .A2(G190), .A3(G200), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n810), .B1(new_n578), .B2(new_n812), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n234), .A2(G179), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n327), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n464), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(G303), .ZN(new_n819));
  NOR2_X1   g0619(.A1(G190), .A2(G200), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n804), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n296), .B1(new_n822), .B2(G311), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n816), .A2(new_n820), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n234), .A2(new_n319), .A3(new_n464), .A4(G200), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G329), .A2(new_n825), .B1(new_n826), .B2(G322), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n819), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n817), .A2(G190), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n815), .B(new_n828), .C1(G283), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n825), .A2(G159), .ZN(new_n831));
  INV_X1    g0631(.A(new_n814), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n831), .A2(KEYINPUT32), .B1(new_n832), .B2(G50), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n428), .B1(new_n822), .B2(G77), .ZN(new_n834));
  INV_X1    g0634(.A(new_n826), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n834), .C1(new_n423), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n818), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n637), .ZN(new_n838));
  INV_X1    g0638(.A(new_n829), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n839), .A2(new_n340), .ZN(new_n840));
  INV_X1    g0640(.A(new_n812), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(G97), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n842), .B1(new_n397), .B2(new_n805), .C1(new_n831), .C2(KEYINPUT32), .ZN(new_n843));
  NOR4_X1   g0643(.A1(new_n836), .A2(new_n838), .A3(new_n840), .A4(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n830), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n786), .B(new_n803), .C1(new_n793), .C2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n735), .A2(new_n736), .A3(new_n792), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n735), .A2(new_n733), .A3(new_n736), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n738), .A2(new_n849), .A3(new_n786), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(G396));
  AND4_X1   g0652(.A1(new_n365), .A2(new_n363), .A3(new_n364), .A4(new_n711), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n365), .A2(new_n710), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n362), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n366), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n692), .B2(new_n710), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n711), .C1(new_n680), .C2(new_n690), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n768), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n785), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n790), .A2(new_n793), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n786), .B1(new_n204), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n793), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n829), .A2(G87), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n867), .B1(new_n868), .B2(new_n824), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT102), .Z(new_n870));
  OAI221_X1 g0670(.A(new_n428), .B1(new_n511), .B2(new_n821), .C1(new_n835), .C2(new_n578), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n832), .A2(G303), .ZN(new_n872));
  INV_X1    g0672(.A(G283), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n842), .B(new_n872), .C1(new_n873), .C2(new_n805), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n871), .B(new_n874), .C1(G107), .C2(new_n818), .ZN(new_n875));
  INV_X1    g0675(.A(G132), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n296), .B1(new_n824), .B2(new_n876), .C1(new_n812), .C2(new_n423), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n839), .A2(new_n397), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n877), .B(new_n878), .C1(G50), .C2(new_n818), .ZN(new_n879));
  AOI22_X1  g0679(.A1(G159), .A2(new_n822), .B1(new_n826), .B2(G143), .ZN(new_n880));
  INV_X1    g0680(.A(G137), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n880), .B1(new_n881), .B2(new_n814), .C1(new_n269), .C2(new_n805), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT34), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n870), .A2(new_n875), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  OAI221_X1 g0684(.A(new_n865), .B1(new_n866), .B2(new_n884), .C1(new_n856), .C2(new_n791), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n863), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(G384));
  INV_X1    g0687(.A(new_n541), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n511), .B(new_n236), .C1(new_n888), .C2(KEYINPUT35), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(KEYINPUT35), .B2(new_n888), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT36), .Z(new_n891));
  OAI211_X1 g0691(.A(new_n231), .B(G77), .C1(new_n397), .C2(new_n423), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(G50), .B2(new_n397), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n312), .A2(G13), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n412), .A2(new_n710), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n445), .B2(new_n460), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT37), .B1(new_n445), .B2(new_n468), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n481), .B(KEYINPUT104), .C1(new_n485), .C2(new_n419), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n703), .B1(new_n707), .B2(new_n709), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n485), .B2(new_n419), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n898), .A2(new_n899), .A3(new_n900), .A4(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n420), .B1(new_n442), .B2(new_n430), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n419), .B1(new_n444), .B2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n901), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n460), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n474), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT37), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n488), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n910), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n474), .B1(new_n445), .B2(new_n460), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n445), .A2(new_n906), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n903), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT105), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n488), .A2(new_n920), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n921), .A2(new_n903), .A3(KEYINPUT105), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n918), .B1(new_n927), .B2(new_n914), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n896), .B(new_n917), .C1(new_n928), .C2(KEYINPUT39), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n659), .A2(new_n901), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n710), .A2(new_n411), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n413), .A2(new_n414), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n932), .B1(new_n395), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT103), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n392), .A2(new_n386), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT79), .B1(new_n375), .B2(KEYINPUT13), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n936), .A2(new_n319), .A3(new_n937), .ZN(new_n938));
  AOI211_X1 g0738(.A(KEYINPUT14), .B(new_n321), .C1(new_n376), .C2(new_n386), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n938), .A2(new_n388), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n411), .ZN(new_n941));
  OAI211_X1 g0741(.A(new_n415), .B(new_n931), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT103), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n943), .B(new_n932), .C1(new_n395), .C2(new_n933), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n935), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n853), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n859), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n915), .A2(new_n916), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n930), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT106), .B1(new_n929), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n779), .A2(new_n490), .A3(new_n781), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n666), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n953), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n760), .B1(new_n758), .B2(new_n710), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n767), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n960), .A2(new_n945), .A3(new_n856), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n949), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n945), .A3(new_n856), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n926), .A2(new_n925), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT105), .B1(new_n921), .B2(new_n903), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n914), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n964), .B1(new_n967), .B2(new_n916), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n963), .B1(new_n968), .B2(new_n962), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n490), .A2(new_n960), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n969), .B(new_n970), .Z(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(new_n733), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n956), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n312), .B2(new_n700), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n956), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n895), .B1(new_n974), .B2(new_n975), .ZN(G367));
  NOR2_X1   g0776(.A1(new_n711), .A2(new_n548), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n574), .A2(new_n977), .B1(new_n573), .B2(new_n711), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n978), .A2(KEYINPUT109), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(KEYINPUT109), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(KEYINPUT42), .B1(new_n981), .B2(new_n727), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n682), .B1(new_n979), .B2(new_n980), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n983), .A2(new_n573), .ZN(new_n984));
  OAI211_X1 g0784(.A(KEYINPUT110), .B(new_n982), .C1(new_n984), .C2(new_n710), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT110), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT42), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n979), .A2(new_n980), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n987), .B1(new_n988), .B2(new_n721), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n710), .B1(new_n983), .B2(new_n573), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n986), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n987), .A3(new_n721), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n985), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n710), .A2(new_n686), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n681), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT107), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n675), .A2(new_n994), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT108), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT108), .B1(new_n996), .B2(new_n997), .ZN(new_n1001));
  NOR3_X1   g0801(.A1(new_n1000), .A2(KEYINPUT43), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(KEYINPUT43), .B2(new_n998), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n985), .A2(new_n991), .A3(new_n992), .A4(new_n1002), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1006), .B1(new_n740), .B2(new_n981), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1004), .A2(new_n739), .A3(new_n988), .A4(new_n1005), .ZN(new_n1008));
  XOR2_X1   g0808(.A(new_n746), .B(KEYINPUT41), .Z(new_n1009));
  NOR3_X1   g0809(.A1(new_n721), .A2(new_n694), .A3(new_n722), .ZN(new_n1010));
  AOI21_X1  g0810(.A(KEYINPUT95), .B1(new_n727), .B2(new_n728), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n988), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n730), .A2(KEYINPUT45), .A3(new_n988), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT44), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n730), .B2(new_n988), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n723), .A2(KEYINPUT44), .A3(new_n729), .A4(new_n981), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1016), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n739), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n718), .A2(new_n720), .A3(new_n712), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n727), .A2(new_n1023), .A3(new_n737), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n737), .B1(new_n727), .B2(new_n1023), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT29), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n773), .A2(new_n774), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n711), .B1(new_n1028), .B2(new_n690), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(KEYINPUT98), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n776), .A2(new_n769), .A3(new_n711), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n861), .B(new_n1026), .C1(new_n1032), .C2(new_n780), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1016), .A2(new_n1020), .A3(new_n740), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1022), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1009), .B1(new_n1036), .B2(new_n782), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1007), .B(new_n1008), .C1(new_n1037), .C2(new_n784), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n241), .A2(new_n797), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n224), .B2(new_n357), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n296), .B1(new_n826), .B2(G303), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n873), .B2(new_n821), .C1(new_n807), .C2(new_n824), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G97), .B2(new_n829), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n805), .A2(new_n578), .B1(new_n814), .B2(new_n868), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G107), .B2(new_n841), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT46), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n837), .B2(new_n511), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n818), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n296), .B1(new_n824), .B2(new_n881), .ZN(new_n1050));
  INV_X1    g0850(.A(G143), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n812), .A2(new_n397), .B1(new_n814), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1050), .B(new_n1052), .C1(G150), .C2(new_n826), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n829), .A2(G77), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(new_n423), .C2(new_n837), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n805), .A2(new_n421), .B1(new_n821), .B2(new_n227), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT111), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1049), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT47), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n785), .B1(new_n795), .B2(new_n1040), .C1(new_n1059), .C2(new_n866), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT112), .Z(new_n1061));
  NAND3_X1  g0861(.A1(new_n996), .A2(new_n792), .A3(new_n997), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1038), .A2(new_n1063), .ZN(G387));
  INV_X1    g0864(.A(new_n742), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n801), .A2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(G107), .B2(new_n224), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n247), .A2(G45), .ZN(new_n1068));
  AOI211_X1 g0868(.A(G45), .B(new_n1065), .C1(G68), .C2(G77), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n355), .A2(G50), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1070), .B(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n798), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1067), .B1(new_n1068), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n818), .A2(G77), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n269), .B2(new_n824), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n812), .A2(new_n357), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n296), .B1(new_n397), .B2(new_n821), .C1(new_n835), .C2(new_n227), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G159), .C2(new_n832), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1076), .A2(KEYINPUT114), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n829), .A2(G97), .B1(new_n265), .B2(new_n806), .ZN(new_n1082));
  AND4_X1   g0882(.A1(new_n1077), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n428), .B1(new_n824), .B2(new_n813), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G303), .A2(new_n822), .B1(new_n826), .B2(G317), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n832), .A2(G322), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(new_n868), .C2(new_n805), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(new_n818), .A2(G294), .B1(G283), .B2(new_n841), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(KEYINPUT49), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n1084), .B(new_n1094), .C1(G116), .C2(new_n829), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1083), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n785), .B1(new_n796), .B2(new_n1074), .C1(new_n1097), .C2(new_n866), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n732), .B2(new_n792), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n784), .B2(new_n1026), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n782), .A2(new_n1026), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1033), .A2(new_n746), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(G393));
  AND3_X1   g0903(.A1(new_n1016), .A2(new_n1020), .A3(new_n740), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n740), .B1(new_n1016), .B2(new_n1020), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n981), .A2(new_n792), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n251), .A2(new_n797), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n538), .B2(new_n224), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n785), .B1(new_n795), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n812), .A2(new_n204), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n296), .B1(new_n824), .B2(new_n1051), .C1(new_n355), .C2(new_n821), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n1111), .B(new_n1112), .C1(G50), .C2(new_n806), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n835), .A2(new_n421), .B1(new_n814), .B2(new_n269), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT51), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n818), .A2(G68), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1115), .A3(new_n867), .A4(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n296), .B(new_n840), .C1(G322), .C2(new_n825), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n835), .A2(new_n868), .B1(new_n814), .B2(new_n807), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT52), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1118), .B(new_n1120), .C1(new_n873), .C2(new_n837), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n812), .A2(new_n511), .B1(new_n821), .B2(new_n578), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G303), .B2(new_n806), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT115), .Z(new_n1124));
  OAI21_X1  g0924(.A(new_n1117), .B1(new_n1121), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1110), .B1(new_n1125), .B2(new_n793), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1106), .A2(new_n784), .B1(new_n1107), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1033), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1128), .A2(new_n1036), .A3(new_n746), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(G390));
  INV_X1    g0930(.A(KEYINPUT118), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1030), .A2(new_n1031), .A3(new_n947), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n855), .A2(new_n366), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(new_n1133), .A3(new_n945), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n928), .A2(new_n896), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT39), .B1(new_n967), .B2(new_n916), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n917), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1137), .A2(new_n1138), .B1(new_n896), .B2(new_n948), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n768), .A2(new_n856), .A3(new_n945), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n917), .B1(new_n928), .B2(KEYINPUT39), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n948), .A2(new_n896), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1142), .A2(new_n1143), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1144));
  NOR4_X1   g0944(.A1(new_n657), .A2(new_n574), .A3(new_n534), .A4(new_n710), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n529), .A2(new_n753), .A3(new_n559), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n755), .B1(new_n750), .B2(new_n751), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n711), .B1(new_n1147), .B2(new_n754), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n959), .B1(new_n1148), .B2(new_n760), .ZN(new_n1149));
  OAI21_X1  g0949(.A(G330), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n942), .A2(new_n944), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n940), .A2(new_n415), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n943), .B1(new_n1152), .B2(new_n932), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n856), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(KEYINPUT116), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G330), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n758), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1157), .A2(new_n957), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n1158), .B2(new_n767), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT116), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n856), .A4(new_n945), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1155), .A2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1141), .B1(new_n1144), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n859), .A2(new_n947), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n945), .B1(new_n768), .B2(new_n856), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT117), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1155), .B(new_n1161), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n946), .B1(new_n1150), .B2(new_n857), .ZN(new_n1171));
  AND2_X1   g0971(.A1(new_n1171), .A2(new_n1140), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n490), .A2(new_n1159), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n954), .A2(new_n1175), .A3(new_n666), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1174), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1131), .B(new_n746), .C1(new_n1163), .C2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1163), .A2(new_n1177), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n746), .B1(new_n1163), .B2(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT118), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1142), .A2(new_n790), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n786), .B1(new_n266), .B2(new_n864), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n818), .A2(G150), .ZN(new_n1185));
  XOR2_X1   g0985(.A(new_n1185), .B(KEYINPUT53), .Z(new_n1186));
  INV_X1    g0986(.A(G128), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n812), .A2(new_n421), .B1(new_n814), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n296), .B1(new_n835), .B2(new_n876), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1188), .B(new_n1189), .C1(G125), .C2(new_n825), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1186), .B(new_n1190), .C1(new_n227), .C2(new_n839), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT54), .B(G143), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n805), .A2(new_n881), .B1(new_n821), .B2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1193), .B(KEYINPUT119), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1111), .B1(G283), .B2(new_n832), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n340), .B2(new_n805), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n296), .B1(new_n826), .B2(G116), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n538), .B2(new_n821), .C1(new_n578), .C2(new_n824), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(new_n838), .A2(new_n1196), .A3(new_n878), .A4(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n1191), .A2(new_n1194), .B1(KEYINPUT120), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(KEYINPUT120), .B2(new_n1199), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1183), .B(new_n1184), .C1(new_n866), .C2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n784), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1202), .B1(new_n1163), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT121), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  OAI211_X1 g1006(.A(KEYINPUT121), .B(new_n1202), .C1(new_n1163), .C2(new_n1203), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(new_n1180), .A2(new_n1182), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(G378));
  INV_X1    g1009(.A(new_n337), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n289), .A2(new_n906), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n337), .B1(new_n289), .B2(new_n906), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n790), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n864), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n785), .B1(new_n1220), .B2(G50), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n829), .A2(new_n440), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n296), .A2(G41), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n825), .A2(G283), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1075), .A2(new_n1222), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT123), .Z(new_n1226));
  OAI22_X1  g1026(.A1(new_n835), .A2(new_n340), .B1(new_n357), .B2(new_n821), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G68), .B2(new_n841), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G97), .A2(new_n806), .B1(new_n832), .B2(G116), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1226), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  AOI211_X1 g1033(.A(G50), .B(new_n1223), .C1(new_n270), .C2(new_n306), .ZN(new_n1234));
  XOR2_X1   g1034(.A(new_n1234), .B(KEYINPUT122), .Z(new_n1235));
  OAI22_X1  g1035(.A1(new_n835), .A2(new_n1187), .B1(new_n821), .B2(new_n881), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G132), .B2(new_n806), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G150), .A2(new_n841), .B1(new_n832), .B2(G125), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1237), .B(new_n1238), .C1(new_n837), .C2(new_n1192), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  AOI211_X1 g1040(.A(G33), .B(G41), .C1(new_n825), .C2(G124), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n839), .B2(new_n421), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1239), .B2(KEYINPUT59), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1235), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1232), .A2(new_n1233), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1221), .B1(new_n1245), .B2(new_n793), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1219), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n969), .A2(G330), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT124), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1217), .A2(new_n1249), .A3(new_n1218), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n929), .A2(new_n950), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT106), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n950), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n969), .A2(new_n1250), .A3(G330), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1252), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n969), .A2(G330), .A3(new_n1250), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1250), .B1(new_n969), .B2(G330), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n1259), .A2(new_n1260), .B1(new_n951), .B2(new_n952), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1247), .B1(new_n1262), .B2(new_n1203), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n954), .A2(new_n666), .A3(new_n1175), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1162), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n768), .A2(new_n856), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n946), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT117), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1162), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1273), .A2(new_n1164), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(new_n1265), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1265), .B1(new_n1268), .B2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1258), .A2(new_n1261), .A3(KEYINPUT57), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n746), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1176), .B1(new_n1163), .B2(new_n1274), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT57), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1264), .B1(new_n1278), .B2(new_n1281), .ZN(G375));
  OAI21_X1  g1082(.A(new_n785), .B1(new_n1220), .B2(G68), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1078), .B1(G116), .B2(new_n806), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n578), .B2(new_n814), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n818), .A2(G97), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n296), .B1(new_n826), .B2(G283), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(G107), .A2(new_n822), .B1(new_n825), .B2(G303), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1054), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n818), .A2(G159), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n428), .B1(new_n822), .B2(G150), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(G128), .A2(new_n825), .B1(new_n826), .B2(G137), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1222), .A2(new_n1290), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n832), .A2(G132), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n1294), .B1(new_n227), .B2(new_n812), .C1(new_n805), .C2(new_n1192), .ZN(new_n1295));
  OAI22_X1  g1095(.A1(new_n1285), .A2(new_n1289), .B1(new_n1293), .B2(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1283), .B1(new_n1296), .B2(new_n793), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1297), .B1(new_n945), .B2(new_n791), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1298), .B1(new_n1274), .B2(new_n1203), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(new_n1275), .A2(new_n1009), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1274), .A2(new_n1265), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1302), .ZN(G381));
  XNOR2_X1  g1103(.A(G375), .B(KEYINPUT125), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n851), .B(new_n1100), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1305));
  OR2_X1    g1105(.A1(G384), .A2(new_n1305), .ZN(new_n1306));
  NOR4_X1   g1106(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1208), .A3(new_n1307), .ZN(G407));
  NAND4_X1  g1108(.A1(new_n1304), .A2(G213), .A3(new_n695), .A4(new_n1208), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(G407), .A3(G213), .ZN(G409));
  NAND3_X1  g1110(.A1(new_n1182), .A2(new_n1179), .A3(new_n1178), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1276), .A2(new_n1262), .A3(new_n1009), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n1311), .B(new_n1312), .C1(new_n1313), .C2(new_n1263), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1314), .B1(G375), .B2(new_n1208), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n695), .A2(G213), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1274), .A2(KEYINPUT60), .A3(new_n1265), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n746), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1177), .A2(KEYINPUT60), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1301), .B2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n886), .B1(new_n1320), .B2(new_n1299), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1318), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1319), .A2(new_n1301), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1299), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(G384), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1315), .A2(new_n1316), .A3(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT62), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n695), .A2(G213), .A3(G2897), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1321), .A2(new_n1325), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1331), .B1(new_n1321), .B2(new_n1325), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1330), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1315), .A2(new_n1336), .A3(new_n1327), .A4(new_n1316), .ZN(new_n1337));
  XOR2_X1   g1137(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1338));
  NAND4_X1  g1138(.A1(new_n1329), .A2(new_n1335), .A3(new_n1337), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1036), .A2(new_n782), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1009), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1340), .B1(new_n1343), .B2(new_n1203), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1063), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(G393), .A2(G396), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1305), .ZN(new_n1347));
  AND3_X1   g1147(.A1(new_n1127), .A2(new_n1129), .A3(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1347), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1349));
  OAI22_X1  g1149(.A1(new_n1344), .A2(new_n1345), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1347), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(G390), .A2(new_n1351), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1127), .A2(new_n1129), .A3(new_n1347), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1352), .A2(new_n1038), .A3(new_n1063), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1339), .A2(new_n1355), .ZN(new_n1356));
  INV_X1    g1156(.A(KEYINPUT61), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1350), .A2(new_n1357), .A3(new_n1354), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT126), .ZN(new_n1359));
  XNOR2_X1  g1159(.A(new_n1358), .B(new_n1359), .ZN(new_n1360));
  NAND4_X1  g1160(.A1(new_n1315), .A2(KEYINPUT63), .A3(new_n1316), .A4(new_n1327), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1328), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT63), .ZN(new_n1363));
  AOI21_X1  g1163(.A(new_n1363), .B1(new_n1330), .B2(new_n1334), .ZN(new_n1364));
  OAI211_X1 g1164(.A(new_n1360), .B(new_n1361), .C1(new_n1362), .C2(new_n1364), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1356), .A2(new_n1365), .ZN(G405));
  OR2_X1    g1166(.A1(G375), .A2(new_n1208), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(G375), .A2(new_n1208), .ZN(new_n1368));
  AND3_X1   g1168(.A1(new_n1367), .A2(new_n1326), .A3(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1326), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1370));
  OR3_X1    g1170(.A1(new_n1369), .A2(new_n1370), .A3(new_n1355), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1355), .B1(new_n1369), .B2(new_n1370), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1371), .A2(new_n1372), .ZN(G402));
endmodule


