//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  AOI21_X1  g007(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(G107), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n189), .B(new_n192), .C1(new_n194), .C2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n191), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT65), .A2(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT65), .A2(G146), .ZN(new_n201));
  OAI21_X1  g015(.A(G143), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n202), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n202), .A2(KEYINPUT70), .A3(new_n205), .A4(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n202), .A2(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT1), .B1(new_n214), .B2(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G128), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n199), .B1(new_n212), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT84), .B1(new_n218), .B2(KEYINPUT10), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT10), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n210), .A2(new_n211), .B1(new_n213), .B2(new_n216), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n199), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G137), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n225), .A2(G134), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT11), .B1(new_n227), .B2(G137), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n225), .A3(G134), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n226), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  OR2_X1    g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n231), .A2(new_n234), .A3(new_n232), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n234), .B1(new_n231), .B2(new_n232), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n233), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n203), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT65), .A2(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n214), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT66), .B1(new_n203), .B2(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT64), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT0), .A3(G128), .ZN(new_n248));
  OR2_X1    g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n246), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n240), .A2(KEYINPUT66), .A3(new_n214), .A4(new_n241), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n244), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT67), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n244), .A2(new_n250), .A3(KEYINPUT67), .A4(new_n251), .ZN(new_n255));
  INV_X1    g069(.A(new_n245), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT65), .B(G146), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n204), .B1(new_n257), .B2(G143), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n254), .A2(new_n255), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT83), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(new_n262), .A3(G101), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n196), .A2(KEYINPUT4), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n190), .B1(new_n191), .B2(G104), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n191), .A2(G104), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n189), .B1(new_n267), .B2(new_n192), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n260), .B(new_n263), .C1(new_n264), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n261), .A2(G101), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n196), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(new_n257), .B2(G143), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n244), .B(new_n251), .C1(new_n274), .C2(new_n206), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n212), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n199), .A2(new_n221), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n259), .A2(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AND3_X1   g092(.A1(new_n224), .A2(new_n238), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n238), .B1(new_n224), .B2(new_n278), .ZN(new_n280));
  INV_X1    g094(.A(G953), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT72), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G953), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G227), .ZN(new_n286));
  XNOR2_X1  g100(.A(G110), .B(G140), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n286), .B(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g103(.A1(new_n279), .A2(new_n280), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n212), .A2(new_n275), .A3(new_n199), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n291), .B1(new_n199), .B2(new_n222), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n231), .A2(new_n232), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(KEYINPUT68), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n231), .A2(new_n234), .A3(new_n232), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT85), .B1(new_n296), .B2(new_n233), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT12), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n212), .A2(new_n275), .A3(new_n199), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n297), .B(KEYINPUT12), .C1(new_n300), .C2(new_n218), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n224), .A2(new_n238), .A3(new_n278), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n288), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n188), .B1(new_n290), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n187), .B1(new_n305), .B2(G469), .ZN(new_n306));
  INV_X1    g120(.A(G469), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT87), .ZN(new_n308));
  OAI211_X1 g122(.A(new_n308), .B(new_n289), .C1(new_n279), .C2(new_n280), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n302), .A2(new_n288), .A3(new_n303), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(KEYINPUT70), .B1(new_n258), .B2(new_n207), .ZN(new_n312));
  INV_X1    g126(.A(new_n211), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n217), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n199), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n220), .B1(new_n316), .B2(new_n221), .ZN(new_n317));
  INV_X1    g131(.A(new_n223), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n278), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n237), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n303), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n308), .B1(new_n321), .B2(new_n289), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n307), .B(new_n188), .C1(new_n311), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n306), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G952), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  INV_X1    g140(.A(G234), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  AOI211_X1 g144(.A(new_n188), .B(new_n285), .C1(G234), .C2(G237), .ZN(new_n331));
  XOR2_X1   g145(.A(KEYINPUT21), .B(G898), .Z(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(G214), .B1(G237), .B2(G902), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(KEYINPUT88), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n254), .A2(new_n255), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n258), .A2(new_n256), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(KEYINPUT89), .A3(G125), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n343));
  INV_X1    g157(.A(G125), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n259), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n212), .A2(new_n344), .A3(new_n275), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(G224), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G953), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n342), .A2(new_n345), .A3(new_n351), .A4(new_n346), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G119), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G116), .ZN(new_n355));
  INV_X1    g169(.A(G116), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G119), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT71), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT2), .B(G113), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n272), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g177(.A(G110), .B(G122), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n355), .A2(new_n357), .A3(KEYINPUT5), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(G113), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n367));
  OAI22_X1  g181(.A1(new_n366), .A2(new_n367), .B1(new_n360), .B2(new_n358), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(new_n199), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n364), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n364), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n361), .B1(new_n269), .B2(new_n271), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n372), .B1(new_n373), .B2(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(KEYINPUT6), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT6), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n376), .B(new_n372), .C1(new_n373), .C2(new_n369), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n353), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT91), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n346), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n346), .A2(new_n380), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n342), .A2(new_n345), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT7), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n349), .B1(KEYINPUT92), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(KEYINPUT92), .B2(new_n384), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n358), .A2(new_n360), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n367), .B1(new_n365), .B2(KEYINPUT90), .ZN(new_n389));
  OR2_X1    g203(.A1(new_n365), .A2(KEYINPUT90), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n391), .A2(new_n199), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n364), .B(KEYINPUT8), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n392), .B(new_n393), .C1(new_n315), .C2(new_n368), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n371), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n387), .B(new_n395), .C1(new_n384), .C2(new_n352), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n379), .A2(new_n396), .A3(new_n188), .ZN(new_n397));
  OAI21_X1  g211(.A(G210), .B1(G237), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(G902), .B1(new_n353), .B2(new_n378), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n398), .A3(new_n396), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n338), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G221), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n404), .B1(new_n406), .B2(new_n188), .ZN(new_n407));
  INV_X1    g221(.A(new_n301), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(new_n298), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n289), .B1(new_n279), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n320), .A2(new_n288), .A3(new_n303), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n307), .B1(new_n412), .B2(new_n188), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n407), .B1(new_n413), .B2(new_n187), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n324), .A2(new_n403), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G122), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G116), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n356), .A2(G122), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n191), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT98), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n417), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n418), .A2(KEYINPUT14), .ZN(new_n423));
  OAI21_X1  g237(.A(G107), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT96), .B1(new_n214), .B2(G128), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT96), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n206), .A3(G143), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n426), .A2(new_n428), .B1(G128), .B2(new_n214), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G134), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT13), .B1(new_n426), .B2(new_n428), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n227), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n429), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n428), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n214), .A2(G128), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n227), .B2(new_n433), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n419), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n191), .B1(new_n417), .B2(new_n418), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT97), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT97), .ZN(new_n446));
  AOI211_X1 g260(.A(new_n446), .B(new_n443), .C1(new_n435), .C2(new_n439), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n432), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G217), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n405), .A2(new_n449), .A3(G953), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n434), .A2(new_n429), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n438), .A2(new_n433), .A3(new_n227), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n444), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n446), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n440), .A2(KEYINPUT97), .A3(new_n444), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n450), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n458), .A3(new_n432), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n451), .A2(new_n459), .A3(new_n188), .ZN(new_n460));
  INV_X1    g274(.A(G478), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT15), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n462), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n451), .A2(new_n459), .A3(new_n188), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n285), .A2(G214), .A3(new_n328), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(new_n214), .ZN(new_n468));
  AOI21_X1  g282(.A(G237), .B1(new_n282), .B2(new_n284), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(G143), .A3(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT18), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(new_n232), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT94), .ZN(new_n476));
  XNOR2_X1  g290(.A(G125), .B(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n257), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G125), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n344), .A2(G140), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G146), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n476), .B1(new_n478), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n478), .A2(new_n483), .A3(new_n476), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n472), .A2(new_n475), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND4_X1   g301(.A1(G143), .A2(new_n285), .A3(G214), .A4(new_n328), .ZN(new_n488));
  AOI21_X1  g302(.A(G143), .B1(new_n469), .B2(G214), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT93), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n490), .A2(new_n491), .A3(new_n473), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n232), .B1(new_n468), .B2(new_n470), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT93), .B1(new_n493), .B2(KEYINPUT18), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n487), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n477), .A2(KEYINPUT16), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT16), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n479), .A3(G125), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n203), .ZN(new_n500));
  OAI211_X1 g314(.A(G146), .B(new_n498), .C1(new_n482), .C2(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(KEYINPUT78), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT78), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n503), .A3(new_n203), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n502), .A2(new_n504), .B1(new_n493), .B2(KEYINPUT17), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n468), .A2(new_n232), .A3(new_n470), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n490), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G113), .B(G122), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(G104), .ZN(new_n511));
  XOR2_X1   g325(.A(new_n511), .B(KEYINPUT95), .Z(new_n512));
  AND3_X1   g326(.A1(new_n495), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n495), .B2(new_n509), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n188), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G475), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT20), .ZN(new_n518));
  INV_X1    g332(.A(new_n486), .ZN(new_n519));
  OAI22_X1  g333(.A1(new_n471), .A2(new_n474), .B1(new_n519), .B2(new_n484), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n491), .B1(new_n490), .B2(new_n473), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n493), .A2(KEYINPUT93), .A3(KEYINPUT18), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n482), .B(KEYINPUT19), .ZN(new_n524));
  INV_X1    g338(.A(new_n257), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n501), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n490), .B2(new_n507), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n511), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n495), .A2(new_n509), .A3(new_n512), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G475), .A2(G902), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n518), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  AOI211_X1 g347(.A(KEYINPUT20), .B(new_n533), .C1(new_n528), .C2(new_n529), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n517), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n415), .A2(new_n466), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n449), .B1(G234), .B2(new_n188), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT23), .B1(new_n354), .B2(G128), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT23), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n206), .A3(G119), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G110), .ZN(new_n542));
  OAI211_X1 g356(.A(new_n541), .B(new_n542), .C1(G119), .C2(new_n206), .ZN(new_n543));
  XNOR2_X1  g357(.A(G119), .B(G128), .ZN(new_n544));
  OR2_X1    g358(.A1(KEYINPUT24), .A2(G110), .ZN(new_n545));
  NAND2_X1  g359(.A1(KEYINPUT24), .A2(G110), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(KEYINPUT76), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT76), .ZN(new_n548));
  AND2_X1   g362(.A1(KEYINPUT24), .A2(G110), .ZN(new_n549));
  NOR2_X1   g363(.A1(KEYINPUT24), .A2(G110), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n543), .B1(new_n552), .B2(KEYINPUT79), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT79), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n554), .B(new_n544), .C1(new_n547), .C2(new_n551), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT80), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n544), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n549), .A2(new_n550), .A3(new_n548), .ZN(new_n558));
  AOI21_X1  g372(.A(KEYINPUT76), .B1(new_n545), .B2(new_n546), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n554), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT80), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n552), .A2(KEYINPUT79), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .A4(new_n543), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n501), .A2(new_n478), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n541), .B1(G119), .B2(new_n206), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT77), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n542), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n568), .B2(new_n567), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n547), .A2(new_n551), .A3(new_n544), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n570), .A2(new_n504), .A3(new_n502), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT82), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT22), .B(G137), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT81), .ZN(new_n578));
  INV_X1    g392(.A(new_n285), .ZN(new_n579));
  NOR3_X1   g393(.A1(new_n579), .A2(new_n404), .A3(new_n327), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n578), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n574), .A2(new_n576), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n566), .A2(new_n572), .A3(new_n575), .A4(new_n581), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(KEYINPUT25), .B1(new_n585), .B2(new_n188), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT25), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n587), .B(G902), .C1(new_n583), .C2(new_n584), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n537), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n537), .A2(G902), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n339), .A2(new_n340), .A3(new_n237), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n227), .A2(G137), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n227), .A2(G137), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n595), .B1(KEYINPUT69), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(KEYINPUT69), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n232), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n294), .B2(new_n295), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n276), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n594), .A2(new_n361), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n469), .A2(G210), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n604), .B(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT73), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n594), .A2(new_n601), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT30), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n594), .A2(KEYINPUT30), .A3(new_n601), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n362), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT73), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n602), .A2(new_n614), .A3(new_n606), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n608), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT31), .ZN(new_n617));
  INV_X1    g431(.A(new_n606), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT28), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n362), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n619), .B1(new_n620), .B2(new_n602), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n602), .A2(new_n619), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n618), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT31), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n608), .A2(new_n613), .A3(new_n625), .A4(new_n615), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n617), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(G472), .A2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT32), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT75), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT75), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(new_n631), .A3(KEYINPUT32), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT32), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n627), .A2(new_n628), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n611), .A2(new_n362), .A3(new_n612), .ZN(new_n636));
  INV_X1    g450(.A(new_n602), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n618), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT29), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n361), .B1(new_n594), .B2(new_n601), .ZN(new_n640));
  OAI21_X1  g454(.A(KEYINPUT28), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n622), .A3(new_n606), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT74), .B1(new_n621), .B2(new_n623), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT74), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n618), .A2(new_n639), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n643), .A2(new_n648), .A3(new_n188), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n634), .A2(new_n635), .B1(new_n649), .B2(G472), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n593), .B1(new_n633), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n536), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G101), .ZN(G3));
  AND2_X1   g467(.A1(new_n324), .A2(new_n414), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n627), .A2(new_n188), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(G472), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n656), .A2(new_n635), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n654), .A2(new_n592), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n400), .A2(new_n402), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n460), .A2(new_n461), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n458), .A2(KEYINPUT100), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  OAI21_X1  g476(.A(KEYINPUT99), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n458), .B1(new_n457), .B2(new_n432), .ZN(new_n664));
  AOI211_X1 g478(.A(new_n450), .B(new_n431), .C1(new_n455), .C2(new_n456), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n663), .B1(KEYINPUT99), .B2(new_n662), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n451), .A2(new_n459), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n188), .A2(G478), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n660), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n535), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n659), .A2(new_n673), .A3(new_n336), .A4(new_n335), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n658), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT34), .B(G104), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  NAND2_X1  g491(.A1(new_n659), .A2(new_n336), .ZN(new_n678));
  INV_X1    g492(.A(new_n535), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n335), .A3(new_n466), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n658), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT35), .B(G107), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G9));
  NOR2_X1   g497(.A1(new_n581), .A2(KEYINPUT36), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n573), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n590), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n589), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n535), .A2(new_n466), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n656), .A2(new_n687), .A3(new_n635), .A4(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n415), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT37), .B(G110), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NAND2_X1  g506(.A1(new_n633), .A2(new_n650), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n589), .A2(new_n686), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n678), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n466), .B(new_n517), .C1(new_n532), .C2(new_n534), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n330), .B1(new_n331), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n693), .A2(new_n654), .A3(new_n695), .A4(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G128), .ZN(G30));
  XOR2_X1   g515(.A(new_n698), .B(KEYINPUT39), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n654), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n616), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n606), .B1(new_n620), .B2(new_n602), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n188), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n635), .A2(new_n634), .B1(G472), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n687), .B1(new_n633), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n659), .B(KEYINPUT38), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(new_n336), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n535), .A2(new_n466), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n705), .A2(new_n710), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n698), .ZN(new_n718));
  AND3_X1   g532(.A1(new_n535), .A2(new_n671), .A3(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n693), .A2(new_n654), .A3(new_n695), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G146), .ZN(G48));
  OAI21_X1  g535(.A(new_n188), .B1(new_n311), .B2(new_n322), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  INV_X1    g537(.A(new_n407), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n323), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n674), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n651), .A2(new_n726), .A3(KEYINPUT101), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT101), .B1(new_n651), .B2(new_n726), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT41), .B(G113), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  AOI21_X1  g545(.A(new_n713), .B1(new_n400), .B2(new_n402), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(new_n723), .A3(new_n323), .A4(new_n724), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n650), .B2(new_n633), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n593), .A2(new_n680), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G116), .ZN(G18));
  NAND4_X1  g551(.A1(new_n734), .A2(new_n335), .A3(new_n688), .A4(new_n687), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G119), .ZN(G21));
  INV_X1    g553(.A(new_n714), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n732), .A2(new_n335), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n725), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n617), .A2(new_n626), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n606), .B1(new_n644), .B2(new_n646), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n628), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n592), .A2(new_n656), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AND4_X1   g562(.A1(new_n656), .A2(new_n687), .A3(new_n719), .A4(new_n745), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n723), .A2(new_n323), .A3(new_n724), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n749), .A2(KEYINPUT102), .A3(new_n750), .A4(new_n732), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT102), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n656), .A2(new_n687), .A3(new_n719), .A4(new_n745), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n752), .B1(new_n733), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G125), .ZN(G27));
  INV_X1    g570(.A(KEYINPUT103), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n290), .B2(new_n304), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n411), .A2(KEYINPUT103), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(G469), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n307), .A2(new_n188), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n323), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n401), .A2(new_n398), .A3(new_n396), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n398), .B1(new_n401), .B2(new_n396), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n764), .A2(new_n765), .A3(new_n713), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n763), .A2(new_n766), .A3(new_n724), .ZN(new_n767));
  INV_X1    g581(.A(new_n719), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(KEYINPUT42), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n693), .A3(new_n592), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n635), .A2(new_n634), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n649), .A2(G472), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n629), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n592), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n763), .A2(new_n766), .A3(new_n724), .A4(new_n719), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT42), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G131), .ZN(G33));
  NAND3_X1  g592(.A1(new_n651), .A2(new_n699), .A3(new_n767), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G134), .ZN(G36));
  NOR2_X1   g594(.A1(new_n290), .A2(new_n757), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n781), .B1(new_n757), .B2(new_n412), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(KEYINPUT45), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n412), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(G469), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT46), .B(new_n762), .C1(new_n783), .C2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT104), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n762), .B1(new_n783), .B2(new_n786), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT46), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n782), .A2(KEYINPUT45), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(G469), .A3(new_n785), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(KEYINPUT104), .A3(KEYINPUT46), .A4(new_n762), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n789), .A2(new_n792), .A3(new_n795), .A4(new_n323), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n724), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n657), .A2(new_n694), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n679), .A2(new_n800), .A3(new_n671), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n535), .A2(KEYINPUT105), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n535), .A2(KEYINPUT105), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n671), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n801), .B1(new_n804), .B2(KEYINPUT43), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n799), .A2(KEYINPUT44), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT44), .B1(new_n799), .B2(new_n805), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n400), .A2(new_n402), .A3(new_n336), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n798), .A2(new_n702), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(KEYINPUT106), .B(G137), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(G39));
  INV_X1    g626(.A(KEYINPUT47), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n796), .B2(new_n724), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n796), .A2(new_n813), .A3(new_n724), .ZN(new_n816));
  NOR4_X1   g630(.A1(new_n693), .A2(new_n592), .A3(new_n808), .A4(new_n768), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G140), .ZN(G42));
  NAND2_X1  g633(.A1(new_n724), .A2(new_n337), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n711), .A2(new_n804), .A3(new_n820), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n633), .A2(new_n592), .A3(new_n709), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n723), .A2(new_n323), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n821), .A2(new_n822), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n672), .A2(new_n696), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n592), .A2(new_n656), .A3(new_n828), .A4(new_n635), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n415), .B1(new_n829), .B2(new_n689), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n651), .B2(new_n536), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n324), .A2(new_n414), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n832), .B1(new_n650), .B2(new_n633), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n688), .A2(new_n766), .A3(new_n687), .A4(new_n718), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n833), .A2(new_n834), .B1(new_n749), .B2(new_n767), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n777), .A2(new_n779), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n734), .A2(new_n735), .B1(new_n746), .B2(new_n742), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n837), .B(new_n738), .C1(new_n727), .C2(new_n728), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n763), .A2(new_n724), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n732), .A2(new_n740), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n698), .B(KEYINPUT107), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n710), .A2(new_n840), .A3(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n755), .A2(new_n700), .A3(new_n720), .A4(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n700), .A2(new_n720), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT52), .A3(new_n755), .A4(new_n844), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n839), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT53), .B1(new_n839), .B2(new_n850), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT108), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n839), .A2(new_n850), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT108), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n827), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT111), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n856), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n839), .A2(new_n850), .A3(KEYINPUT53), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n827), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n725), .A2(new_n329), .A3(new_n808), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n864), .A2(new_n805), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n656), .A3(new_n687), .A4(new_n745), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n535), .A2(new_n671), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n822), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n805), .A2(new_n330), .A3(new_n746), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n870), .A2(new_n713), .A3(new_n712), .A4(new_n750), .ZN(new_n871));
  NOR2_X1   g685(.A1(KEYINPUT110), .A2(KEYINPUT50), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT109), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n823), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n823), .A2(new_n876), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n878), .A2(new_n724), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n815), .B2(new_n816), .ZN(new_n881));
  INV_X1    g695(.A(new_n870), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n882), .A2(new_n808), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n875), .B(KEYINPUT51), .C1(new_n881), .C2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n865), .A2(new_n592), .A3(new_n773), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT48), .Z(new_n887));
  NAND3_X1  g701(.A1(new_n822), .A2(new_n864), .A3(new_n673), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n326), .B(new_n888), .C1(new_n882), .C2(new_n733), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n816), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n814), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n883), .B1(new_n893), .B2(new_n880), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT51), .B1(new_n894), .B2(new_n875), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n858), .A2(new_n859), .A3(new_n863), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n325), .A2(new_n281), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT112), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n860), .A2(new_n855), .A3(new_n861), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n851), .B1(new_n852), .B2(KEYINPUT108), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n862), .B1(new_n903), .B2(new_n827), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n859), .B1(new_n904), .B2(new_n896), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n826), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(KEYINPUT113), .B(new_n826), .C1(new_n900), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(G75));
  INV_X1    g724(.A(KEYINPUT115), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n853), .A2(new_n857), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n353), .B(new_n378), .ZN(new_n915));
  XOR2_X1   g729(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n916));
  XNOR2_X1  g730(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n913), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n285), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n918), .B1(new_n913), .B2(new_n914), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n911), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n923), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n925), .A2(KEYINPUT115), .A3(new_n921), .A4(new_n919), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n924), .A2(new_n926), .ZN(G51));
  NOR3_X1   g741(.A1(new_n903), .A2(new_n188), .A3(new_n794), .ZN(new_n928));
  XNOR2_X1  g742(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n761), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n903), .A2(new_n827), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT54), .B1(new_n901), .B2(new_n902), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n311), .A2(new_n322), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n928), .B1(new_n935), .B2(KEYINPUT117), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n933), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n920), .B1(new_n936), .B2(new_n938), .ZN(G54));
  NAND4_X1  g753(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n940));
  INV_X1    g754(.A(new_n530), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n920), .ZN(G60));
  XNOR2_X1  g758(.A(new_n669), .B(KEYINPUT118), .ZN(new_n945));
  INV_X1    g759(.A(new_n904), .ZN(new_n946));
  NAND2_X1  g760(.A1(G478), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT59), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n945), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n931), .A2(new_n932), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n945), .A2(new_n948), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n920), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT60), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n912), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n585), .B(KEYINPUT119), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT120), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n912), .A2(new_n685), .A3(new_n954), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n958), .A2(KEYINPUT61), .A3(new_n921), .A4(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n957), .A2(KEYINPUT120), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n921), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n955), .B2(new_n956), .ZN(new_n963));
  OAI22_X1  g777(.A1(new_n960), .A2(new_n961), .B1(new_n963), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g778(.A(new_n831), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n838), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n579), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT121), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n333), .B2(new_n348), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(G898), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n378), .B1(new_n971), .B2(new_n579), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT122), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n970), .B(new_n973), .ZN(G69));
  AOI21_X1  g788(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n703), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n651), .A3(new_n766), .A4(new_n828), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n818), .A2(new_n810), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n848), .A2(new_n755), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n716), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT62), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n980), .A2(new_n716), .A3(KEYINPUT62), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n285), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT125), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n611), .A2(new_n612), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n524), .B(KEYINPUT123), .Z(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT124), .Z(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n987), .A2(new_n988), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n579), .B1(new_n979), .B2(new_n985), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT125), .B1(new_n995), .B2(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n579), .A2(G900), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n980), .A2(new_n777), .A3(new_n779), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n774), .A2(new_n841), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n798), .A2(new_n702), .A3(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1000), .A2(new_n810), .A3(new_n818), .A4(new_n1002), .ZN(new_n1003));
  OAI211_X1 g817(.A(new_n991), .B(new_n999), .C1(new_n1003), .C2(new_n579), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n997), .A2(new_n998), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n998), .B1(new_n997), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n976), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n997), .A2(new_n1004), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n997), .A2(new_n998), .A3(new_n1004), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1009), .A2(new_n975), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1007), .A2(new_n1011), .ZN(G72));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  INV_X1    g828(.A(new_n966), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1003), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1016), .A2(new_n602), .A3(new_n618), .A4(new_n613), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n638), .A2(new_n616), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1014), .B(new_n1018), .C1(new_n851), .C2(new_n852), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1017), .A2(new_n921), .A3(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n606), .B1(new_n636), .B2(new_n637), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1014), .B1(new_n986), .B2(new_n1015), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1020), .B1(new_n1024), .B2(new_n1025), .ZN(G57));
endmodule


