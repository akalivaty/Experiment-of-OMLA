//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT68), .B(KEYINPUT27), .Z(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(new_n198), .B2(G146), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n196), .A2(KEYINPUT64), .A3(G143), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n194), .B1(new_n197), .B2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n200), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT11), .ZN(new_n208));
  INV_X1    g022(.A(G134), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G137), .ZN(new_n210));
  INV_X1    g024(.A(G137), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT11), .A3(G134), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G137), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n210), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n209), .A2(G137), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n211), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT66), .B1(new_n207), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G119), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G116), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT65), .B(G116), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n223), .B1(new_n224), .B2(G119), .ZN(new_n225));
  XOR2_X1   g039(.A(KEYINPUT2), .B(G113), .Z(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT65), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n231), .A3(G119), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n226), .A2(new_n232), .A3(new_n222), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g048(.A1(new_n215), .A2(new_n218), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n195), .A2(new_n197), .A3(new_n199), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n198), .A2(G146), .ZN(new_n237));
  OAI21_X1  g051(.A(KEYINPUT64), .B1(new_n196), .B2(G143), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n201), .A2(new_n198), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n236), .B1(new_n240), .B2(new_n205), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n197), .A2(new_n199), .A3(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n245), .B1(new_n204), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n210), .A2(new_n212), .A3(new_n214), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n215), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n220), .A2(new_n234), .A3(new_n243), .A4(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n235), .A2(new_n241), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n234), .B1(new_n256), .B2(new_n252), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n234), .A2(new_n252), .A3(new_n256), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n193), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT30), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n252), .A2(new_n264), .A3(new_n256), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n220), .A2(new_n243), .A3(new_n252), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(KEYINPUT30), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n263), .B1(new_n267), .B2(new_n234), .ZN(new_n268));
  INV_X1    g082(.A(new_n234), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n243), .A2(new_n252), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n264), .B1(new_n270), .B2(new_n220), .ZN(new_n271));
  OAI211_X1 g085(.A(KEYINPUT67), .B(new_n269), .C1(new_n271), .C2(new_n265), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  INV_X1    g087(.A(new_n193), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n273), .B1(new_n254), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n253), .A2(new_n193), .A3(KEYINPUT69), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n268), .A2(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n262), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n276), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n266), .A2(KEYINPUT30), .ZN(new_n284));
  INV_X1    g098(.A(new_n265), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT67), .B1(new_n286), .B2(new_n269), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n263), .B(new_n234), .C1(new_n284), .C2(new_n285), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n281), .B(new_n283), .C1(new_n287), .C2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n279), .B1(new_n282), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT72), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n187), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(G472), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n255), .A2(new_n260), .A3(new_n193), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n254), .B1(new_n268), .B2(new_n272), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n193), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n266), .A2(new_n269), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n253), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(KEYINPUT28), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n259), .A2(new_n258), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n274), .A2(new_n297), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n295), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n268), .A2(new_n272), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n283), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n261), .B1(new_n310), .B2(KEYINPUT31), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n280), .B1(new_n277), .B2(new_n281), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n293), .A2(new_n187), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n308), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n294), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT82), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT82), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n197), .A2(new_n321), .A3(KEYINPUT1), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(G128), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n197), .A2(new_n199), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n200), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n326));
  INV_X1    g140(.A(G104), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n326), .B1(new_n327), .B2(G107), .ZN(new_n328));
  INV_X1    g142(.A(G107), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT3), .A3(G104), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(KEYINPUT80), .A2(G101), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT80), .A2(G101), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT79), .B1(new_n329), .B2(G104), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n327), .A3(G107), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n334), .A3(new_n335), .A4(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT81), .B1(new_n329), .B2(G104), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n340), .A2(new_n327), .A3(G107), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n329), .A2(G104), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G101), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n318), .B1(new_n325), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n251), .A2(KEYINPUT84), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT84), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n250), .A2(new_n348), .A3(new_n215), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT4), .ZN(new_n351));
  INV_X1    g165(.A(new_n331), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n335), .A2(new_n337), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n351), .B(G101), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n355));
  INV_X1    g169(.A(G101), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n335), .A2(new_n337), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(new_n331), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n248), .B(new_n354), .C1(new_n355), .C2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n241), .A2(KEYINPUT10), .A3(new_n338), .A4(new_n344), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n346), .A2(new_n350), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G953), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(G227), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT78), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  XOR2_X1   g179(.A(new_n364), .B(new_n365), .Z(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n345), .A2(new_n207), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n345), .B2(new_n325), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT85), .B1(new_n250), .B2(new_n215), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n370), .A2(KEYINPUT12), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n369), .A2(new_n251), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n251), .ZN(new_n373));
  INV_X1    g187(.A(new_n371), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n367), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n346), .A2(new_n359), .A3(new_n360), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n378));
  AND3_X1   g192(.A1(new_n377), .A2(new_n378), .A3(new_n251), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n377), .B2(new_n251), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n361), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n366), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n376), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XOR2_X1   g197(.A(KEYINPUT88), .B(G469), .Z(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n383), .A2(G902), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G902), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n369), .A2(new_n251), .A3(new_n371), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n371), .B1(new_n369), .B2(new_n251), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n361), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n382), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n361), .A2(new_n366), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n379), .B2(new_n380), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n391), .A2(KEYINPUT87), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT87), .B1(new_n391), .B2(new_n393), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n386), .B1(new_n396), .B2(G469), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT98), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n229), .A2(new_n231), .A3(G122), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n228), .A2(G122), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G107), .B1(new_n399), .B2(new_n400), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n198), .A2(G128), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n194), .A2(G143), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G134), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n405), .A2(new_n406), .A3(new_n209), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n399), .A2(new_n329), .A3(new_n401), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n224), .A2(KEYINPUT14), .A3(G122), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n413), .A2(KEYINPUT98), .A3(G107), .A4(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n404), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT13), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n417), .B1(new_n194), .B2(G143), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n194), .A2(G143), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT97), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(KEYINPUT13), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NOR3_X1   g236(.A1(new_n418), .A2(KEYINPUT97), .A3(new_n419), .ZN(new_n423));
  OAI21_X1  g237(.A(G134), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n399), .A2(new_n401), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(G107), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n411), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(new_n409), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT9), .B(G234), .ZN(new_n429));
  INV_X1    g243(.A(G217), .ZN(new_n430));
  NOR3_X1   g244(.A1(new_n429), .A2(new_n430), .A3(G953), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n416), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(KEYINPUT99), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT99), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n416), .A2(new_n428), .A3(new_n434), .A4(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n416), .A2(new_n428), .ZN(new_n436));
  INV_X1    g250(.A(new_n431), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n433), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT100), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n387), .ZN(new_n441));
  INV_X1    g255(.A(G478), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(KEYINPUT15), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n443), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n439), .A2(new_n440), .A3(new_n387), .A4(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g261(.A(G113), .B(G122), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(new_n327), .ZN(new_n449));
  INV_X1    g263(.A(G237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n362), .A3(G214), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G143), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n189), .B(G214), .C1(new_n452), .C2(G143), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT18), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n213), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(G140), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G125), .ZN(new_n461));
  INV_X1    g275(.A(G125), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(G146), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n463), .A3(new_n196), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n454), .B(new_n455), .C1(new_n457), .C2(new_n213), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n459), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n456), .A2(G131), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT17), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n454), .A2(new_n455), .A3(new_n213), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n213), .B1(new_n454), .B2(new_n455), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT17), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT16), .ZN(new_n477));
  OR3_X1    g291(.A1(new_n462), .A2(KEYINPUT16), .A3(G140), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(G146), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT75), .ZN(new_n480));
  AOI21_X1  g294(.A(G146), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT75), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(new_n478), .A3(new_n483), .A4(G146), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n449), .B(new_n469), .C1(new_n476), .C2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n477), .A2(G146), .A3(new_n478), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n481), .B1(new_n488), .B2(new_n483), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n473), .A2(new_n489), .A3(new_n480), .A4(new_n475), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n449), .B1(new_n490), .B2(new_n469), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n387), .B1(new_n487), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(G475), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT19), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT19), .B1(new_n461), .B2(new_n463), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n196), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n454), .A2(new_n455), .A3(new_n213), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n496), .B(new_n479), .C1(new_n497), .C2(new_n474), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(KEYINPUT94), .A3(new_n469), .ZN(new_n499));
  INV_X1    g313(.A(new_n449), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT94), .B1(new_n498), .B2(new_n469), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n486), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT20), .ZN(new_n504));
  INV_X1    g318(.A(G475), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n387), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT95), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n504), .B1(new_n503), .B2(new_n507), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n493), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT96), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT96), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n493), .B(new_n512), .C1(new_n508), .C2(new_n509), .ZN(new_n513));
  NAND2_X1  g327(.A1(G234), .A2(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(G952), .A3(new_n362), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT21), .B(G898), .Z(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(G902), .A3(G953), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n447), .A2(new_n511), .A3(new_n513), .A4(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G221), .B1(new_n429), .B2(G902), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n397), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(G217), .A2(G902), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n430), .B2(G234), .ZN(new_n524));
  XOR2_X1   g338(.A(new_n524), .B(KEYINPUT73), .Z(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n194), .A2(G119), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n221), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT24), .B(G110), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n532), .A3(KEYINPUT74), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(new_n529), .B2(new_n531), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n536));
  INV_X1    g350(.A(new_n527), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n536), .B(new_n528), .C1(new_n537), .C2(KEYINPUT23), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n533), .A2(new_n535), .B1(G110), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n485), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n538), .A2(G110), .B1(new_n532), .B2(new_n530), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n479), .A3(new_n466), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n362), .A2(G221), .A3(G234), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n542), .A3(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n526), .B1(new_n550), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT76), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n525), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n550), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(KEYINPUT25), .A3(new_n387), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(KEYINPUT76), .A3(new_n551), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n525), .A2(new_n387), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT77), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n232), .A2(KEYINPUT5), .A3(new_n222), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n222), .A2(KEYINPUT5), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(G113), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n225), .A2(new_n226), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n569), .A2(new_n570), .A3(new_n338), .A4(new_n344), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n354), .B1(new_n227), .B2(new_n233), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n355), .A2(new_n358), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G122), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n575), .B(new_n571), .C1(new_n572), .C2(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(KEYINPUT6), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT6), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n574), .A2(new_n580), .A3(new_n576), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n462), .B(new_n236), .C1(new_n240), .C2(new_n205), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n582), .B1(new_n248), .B2(new_n462), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n362), .A2(G224), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n583), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n579), .A2(new_n581), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT89), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n575), .B(KEYINPUT8), .Z(new_n591));
  AOI22_X1  g405(.A1(new_n569), .A2(new_n570), .B1(new_n338), .B2(new_n344), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT90), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(G113), .B1(new_n222), .B2(KEYINPUT5), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n225), .B2(KEYINPUT5), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n345), .B1(new_n596), .B2(new_n233), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n597), .A2(new_n571), .A3(KEYINPUT90), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n590), .B1(new_n594), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT7), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n585), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n583), .A2(new_n601), .ZN(new_n602));
  OAI221_X1 g416(.A(new_n582), .B1(new_n600), .B2(new_n585), .C1(new_n248), .C2(new_n462), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n578), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n594), .A2(new_n590), .A3(new_n598), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n579), .A2(KEYINPUT89), .A3(new_n581), .A4(new_n586), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n589), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT92), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n589), .A2(new_n608), .A3(new_n614), .A4(new_n609), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n589), .A2(new_n608), .A3(new_n612), .A4(new_n609), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n566), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n317), .A2(new_n522), .A3(new_n564), .A4(new_n618), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(new_n334), .Z(G3));
  NOR2_X1   g434(.A1(new_n291), .A2(G902), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n621), .A2(new_n295), .B1(new_n293), .B2(new_n291), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n377), .A2(new_n251), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n377), .A2(new_n378), .A3(new_n251), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n366), .B1(new_n626), .B2(new_n361), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n387), .B(new_n384), .C1(new_n627), .C2(new_n376), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT87), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n375), .A2(new_n372), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n366), .B1(new_n630), .B2(new_n361), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n367), .B1(new_n624), .B2(new_n625), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n391), .A2(KEYINPUT87), .A3(new_n393), .ZN(new_n634));
  AOI21_X1  g448(.A(G902), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(G469), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n628), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n564), .A2(new_n637), .A3(new_n520), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT101), .B1(new_n622), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n290), .A2(new_n282), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n293), .B1(new_n640), .B2(new_n311), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n314), .A2(new_n387), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n641), .B1(new_n642), .B2(G472), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n397), .A2(new_n563), .A3(new_n521), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT101), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n610), .A2(new_n613), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n566), .B1(new_n648), .B2(new_n617), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT33), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n436), .B2(new_n437), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n439), .A2(new_n650), .B1(new_n432), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n442), .A2(G902), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n439), .A2(new_n387), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n652), .A2(new_n653), .B1(new_n442), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n511), .B2(new_n513), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n649), .A2(new_n518), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n649), .A2(KEYINPUT102), .A3(new_n518), .A4(new_n656), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n647), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NAND2_X1  g478(.A1(new_n444), .A2(new_n446), .ZN(new_n665));
  INV_X1    g479(.A(new_n491), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n486), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n505), .B1(new_n667), .B2(new_n387), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n503), .A2(new_n507), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT20), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n503), .A2(new_n504), .A3(new_n507), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n668), .A2(KEYINPUT103), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n668), .A2(KEYINPUT103), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n518), .B(KEYINPUT104), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n665), .A2(new_n672), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n649), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n647), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT35), .B(G107), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  NOR2_X1   g494(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n543), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n540), .A2(new_n542), .A3(new_n681), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n560), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT105), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n554), .B2(new_n557), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n643), .A2(new_n522), .A3(new_n618), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT37), .B(G110), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(KEYINPUT106), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n689), .B(new_n691), .ZN(G12));
  OAI21_X1  g506(.A(new_n515), .B1(new_n517), .B2(G900), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT107), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n665), .A2(new_n672), .A3(new_n673), .A4(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n649), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n397), .A2(new_n521), .A3(new_n687), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n649), .A2(new_n696), .A3(KEYINPUT108), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n317), .A2(new_n699), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  NAND2_X1  g517(.A1(new_n302), .A2(new_n274), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n310), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n295), .B1(new_n705), .B2(new_n387), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n314), .B2(new_n315), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n294), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT109), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n294), .A2(new_n707), .A3(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT38), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n616), .A2(new_n713), .A3(new_n617), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n713), .B1(new_n616), .B2(new_n617), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT110), .B(KEYINPUT39), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n694), .B(new_n716), .Z(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n637), .A2(new_n520), .A3(new_n718), .ZN(new_n719));
  OAI22_X1  g533(.A1(new_n714), .A2(new_n715), .B1(new_n719), .B2(KEYINPUT40), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n511), .A2(new_n513), .B1(new_n446), .B2(new_n444), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n565), .A3(new_n687), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n719), .B2(KEYINPUT40), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n712), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT111), .B(G143), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G45));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n511), .A2(new_n513), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n654), .A2(new_n442), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n439), .A2(new_n650), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n651), .A2(new_n432), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n653), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n730), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AND4_X1   g549(.A1(new_n728), .A2(new_n729), .A3(new_n735), .A4(new_n695), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n728), .B1(new_n656), .B2(new_n695), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n317), .A3(new_n649), .A4(new_n700), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  INV_X1    g554(.A(new_n661), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n563), .B1(new_n294), .B2(new_n316), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n383), .B2(G902), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n743), .A2(new_n628), .A3(new_n520), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT41), .B(G113), .Z(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NOR2_X1   g562(.A1(new_n745), .A2(new_n676), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n228), .ZN(G18));
  AND2_X1   g564(.A1(new_n744), .A2(new_n649), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n519), .A2(new_n687), .ZN(new_n752));
  INV_X1    g566(.A(new_n308), .ZN(new_n753));
  INV_X1    g567(.A(new_n315), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n753), .B1(new_n291), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n293), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT32), .B1(new_n314), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n751), .B(new_n752), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  NAND2_X1  g573(.A1(new_n649), .A2(new_n722), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n743), .A2(new_n628), .A3(new_n520), .A4(new_n674), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n193), .B1(new_n303), .B2(new_n304), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n763), .B1(new_n310), .B2(KEYINPUT31), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n293), .B1(new_n640), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT113), .B(G472), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n765), .B1(new_n642), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n762), .A2(new_n767), .A3(new_n564), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G122), .ZN(G24));
  NAND4_X1  g583(.A1(new_n738), .A2(new_n688), .A3(new_n767), .A4(new_n751), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G125), .ZN(G27));
  AOI22_X1  g585(.A1(new_n626), .A2(new_n392), .B1(new_n390), .B2(new_n382), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n772), .B2(G902), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n521), .B1(new_n628), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n617), .A2(new_n565), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n616), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT114), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n616), .A2(new_n774), .A3(KEYINPUT114), .A4(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n742), .A3(new_n738), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT115), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT42), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n784), .A3(new_n742), .A4(new_n738), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n738), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n783), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n317), .A2(new_n564), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT116), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n742), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n788), .A2(new_n790), .A3(new_n780), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G131), .ZN(G33));
  NAND3_X1  g609(.A1(new_n780), .A2(new_n742), .A3(new_n696), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G134), .ZN(G36));
  NAND3_X1  g611(.A1(new_n735), .A2(new_n511), .A3(new_n513), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT43), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT43), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n688), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT44), .B1(new_n802), .B2(new_n622), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n801), .A2(new_n643), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n616), .A2(new_n775), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n394), .A2(new_n395), .ZN(new_n809));
  OAI211_X1 g623(.A(KEYINPUT117), .B(G469), .C1(new_n809), .C2(KEYINPUT45), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n633), .B2(new_n634), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(new_n636), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n772), .A2(KEYINPUT45), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(G469), .A2(G902), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT46), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n808), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n386), .B1(new_n817), .B2(new_n818), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n815), .A2(KEYINPUT118), .A3(KEYINPUT46), .A4(new_n816), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n819), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n807), .A2(new_n520), .A3(new_n718), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NOR4_X1   g638(.A1(new_n787), .A2(new_n317), .A3(new_n564), .A4(new_n806), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n822), .A2(KEYINPUT47), .A3(new_n520), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT47), .B1(new_n822), .B2(new_n520), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NOR4_X1   g643(.A1(new_n563), .A2(new_n798), .A3(new_n566), .A4(new_n521), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n743), .A2(new_n628), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT119), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n832), .B2(KEYINPUT49), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n833), .B1(KEYINPUT49), .B2(new_n832), .ZN(new_n834));
  INV_X1    g648(.A(new_n712), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n714), .A2(new_n715), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n515), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n799), .A2(new_n838), .A3(new_n800), .ZN(new_n839));
  INV_X1    g653(.A(new_n766), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n314), .B2(new_n387), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n839), .A2(new_n563), .A3(new_n765), .A4(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n831), .A2(new_n565), .A3(new_n521), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(KEYINPUT50), .A3(new_n836), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT50), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n799), .A2(new_n800), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n846), .A2(new_n564), .A3(new_n838), .A4(new_n767), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n836), .A2(new_n843), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n841), .A2(new_n687), .A3(new_n765), .ZN(new_n850));
  NOR4_X1   g664(.A1(new_n839), .A2(new_n521), .A3(new_n831), .A4(new_n806), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n844), .A2(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n806), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n564), .A2(new_n853), .A3(new_n838), .A4(new_n744), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n835), .A2(KEYINPUT122), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n854), .A2(new_n710), .A3(new_n711), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n729), .A2(new_n735), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n832), .A2(new_n520), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n826), .A2(new_n827), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n842), .A2(new_n853), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n861), .B(KEYINPUT51), .C1(new_n863), .C2(new_n864), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n790), .A2(new_n792), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n851), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n855), .A2(new_n858), .A3(new_n656), .ZN(new_n872));
  INV_X1    g686(.A(G952), .ZN(new_n873));
  AOI211_X1 g687(.A(new_n873), .B(G953), .C1(new_n842), .C2(new_n751), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n867), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n780), .A2(new_n738), .A3(new_n850), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n672), .A2(new_n673), .A3(new_n695), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n806), .A2(new_n665), .A3(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n317), .A3(new_n700), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n796), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n796), .A2(new_n878), .A3(KEYINPUT120), .A4(new_n881), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n794), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n745), .B1(new_n741), .B2(new_n676), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n619), .A2(new_n689), .A3(new_n768), .A4(new_n758), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n694), .B(KEYINPUT121), .Z(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AOI211_X1 g706(.A(new_n686), .B(new_n892), .C1(new_n554), .C2(new_n557), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n649), .A2(new_n893), .A3(new_n774), .A4(new_n722), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n708), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n739), .A2(new_n770), .A3(new_n702), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT52), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(new_n708), .B2(new_n894), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n739), .A2(new_n770), .A3(new_n898), .A4(new_n702), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n729), .A2(new_n735), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n511), .A2(new_n665), .A3(new_n513), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n903), .A2(new_n618), .A3(new_n674), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n904), .A2(new_n639), .A3(new_n646), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n890), .A2(new_n897), .A3(new_n899), .A4(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT53), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n887), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI22_X1  g722(.A1(new_n884), .A2(new_n885), .B1(new_n786), .B2(new_n793), .ZN(new_n909));
  AND4_X1   g723(.A1(new_n619), .A2(new_n689), .A3(new_n768), .A4(new_n758), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n742), .B(new_n744), .C1(new_n661), .C2(new_n677), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n899), .A3(new_n905), .A4(new_n911), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n896), .A2(KEYINPUT52), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n909), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n877), .B1(new_n908), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n907), .B1(new_n887), .B2(new_n906), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n909), .A2(new_n914), .A3(KEYINPUT53), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(KEYINPUT54), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n876), .B1(new_n916), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n837), .B1(new_n920), .B2(new_n921), .ZN(G75));
  NAND2_X1  g736(.A1(new_n873), .A2(G953), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT123), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n579), .A2(new_n581), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n586), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT55), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n917), .A2(new_n918), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n929), .A2(G210), .A3(G902), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n930), .B2(KEYINPUT56), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n387), .B1(new_n917), .B2(new_n918), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(G210), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT56), .ZN(new_n934));
  INV_X1    g748(.A(new_n928), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n925), .B1(new_n931), .B2(new_n936), .ZN(G51));
  INV_X1    g751(.A(new_n815), .ZN(new_n938));
  OAI211_X1 g752(.A(G902), .B(new_n938), .C1(new_n908), .C2(new_n915), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n932), .B2(new_n938), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n816), .B(KEYINPUT57), .Z(new_n944));
  NAND3_X1  g758(.A1(new_n916), .A2(new_n919), .A3(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n383), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n925), .B1(new_n943), .B2(new_n947), .ZN(G54));
  NAND4_X1  g762(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n949), .A2(new_n503), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n503), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n925), .B1(new_n950), .B2(new_n951), .ZN(G60));
  XNOR2_X1  g766(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n442), .A2(new_n387), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n916), .A2(new_n919), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n733), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n916), .A2(new_n652), .A3(new_n919), .A4(new_n955), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n957), .A2(new_n924), .A3(new_n958), .ZN(G63));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n523), .B(KEYINPUT60), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n917), .B2(new_n918), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n683), .A2(new_n684), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n924), .B1(new_n962), .B2(new_n555), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n962), .A2(new_n555), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(KEYINPUT61), .A3(new_n924), .A4(new_n964), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(G66));
  AOI21_X1  g784(.A(new_n362), .B1(new_n516), .B2(G224), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n890), .A2(new_n905), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n973), .B2(new_n362), .ZN(new_n974));
  INV_X1    g788(.A(G898), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n926), .B1(new_n975), .B2(G953), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n974), .B(new_n976), .ZN(G69));
  OR2_X1    g791(.A1(new_n494), .A2(new_n495), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n286), .B(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n362), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n739), .A2(new_n702), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT62), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n725), .A2(new_n982), .A3(new_n983), .A4(new_n770), .ZN(new_n984));
  OR4_X1    g798(.A1(new_n789), .A2(new_n719), .A3(new_n806), .A4(new_n902), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n823), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n986), .A2(new_n828), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n725), .A2(new_n982), .A3(new_n770), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT126), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT126), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(new_n991), .A3(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n981), .B1(new_n987), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n822), .A2(new_n520), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n869), .A2(new_n649), .A3(new_n722), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n718), .B(new_n995), .C1(new_n996), .C2(new_n807), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n982), .A2(new_n770), .A3(new_n796), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n998), .B1(new_n786), .B2(new_n793), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n997), .A2(new_n362), .A3(new_n828), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G900), .A2(G953), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n980), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n362), .B1(G227), .B2(G900), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n994), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1005));
  NAND2_X1  g819(.A1(G227), .A2(G900), .ZN(new_n1006));
  AND4_X1   g820(.A1(G953), .A2(new_n1005), .A3(new_n1006), .A4(new_n979), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n1004), .A2(new_n1007), .ZN(G72));
  NAND4_X1  g822(.A1(new_n993), .A2(new_n986), .A3(new_n828), .A4(new_n972), .ZN(new_n1009));
  NAND2_X1  g823(.A1(G472), .A2(G902), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT63), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n299), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n193), .A3(new_n1013), .ZN(new_n1014));
  AND4_X1   g828(.A1(new_n828), .A2(new_n997), .A3(new_n972), .A4(new_n999), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1011), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n274), .B(new_n299), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1014), .A2(new_n924), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1013), .A2(new_n274), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1016), .B1(new_n1019), .B2(new_n310), .ZN(new_n1020));
  AND3_X1   g834(.A1(new_n929), .A2(KEYINPUT127), .A3(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(KEYINPUT127), .B1(new_n929), .B2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1018), .A2(new_n1023), .ZN(G57));
endmodule


