

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  INV_X1 U323 ( .A(n586), .ZN(n480) );
  XNOR2_X1 U324 ( .A(KEYINPUT38), .B(n484), .ZN(n520) );
  XOR2_X1 U325 ( .A(n492), .B(KEYINPUT28), .Z(n544) );
  XNOR2_X1 U326 ( .A(n447), .B(n325), .ZN(n540) );
  NOR2_X1 U327 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U328 ( .A(n389), .B(KEYINPUT32), .ZN(n390) );
  XNOR2_X1 U329 ( .A(n391), .B(n390), .ZN(n393) );
  XOR2_X1 U330 ( .A(G15GAT), .B(G1GAT), .Z(n371) );
  NAND2_X1 U331 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U332 ( .A(n317), .B(n316), .ZN(n319) );
  XNOR2_X1 U333 ( .A(n319), .B(n318), .ZN(n324) );
  XOR2_X1 U334 ( .A(n399), .B(n398), .Z(n578) );
  NOR2_X1 U335 ( .A1(n475), .A2(n451), .ZN(n548) );
  INV_X1 U336 ( .A(G36GAT), .ZN(n485) );
  XNOR2_X1 U337 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U338 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U339 ( .A(n485), .B(KEYINPUT108), .ZN(n486) );
  XNOR2_X1 U340 ( .A(n498), .B(n497), .ZN(G1349GAT) );
  XNOR2_X1 U341 ( .A(n487), .B(n486), .ZN(G1329GAT) );
  XNOR2_X1 U342 ( .A(G148GAT), .B(KEYINPUT72), .ZN(n291) );
  XNOR2_X1 U343 ( .A(n291), .B(KEYINPUT73), .ZN(n292) );
  XOR2_X1 U344 ( .A(n292), .B(G204GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(G78GAT), .B(G106GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n382) );
  XOR2_X1 U347 ( .A(KEYINPUT90), .B(G218GAT), .Z(n296) );
  XNOR2_X1 U348 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U350 ( .A(G197GAT), .B(n297), .Z(n443) );
  XNOR2_X1 U351 ( .A(n382), .B(n443), .ZN(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n299) );
  XOR2_X1 U353 ( .A(G141GAT), .B(G22GAT), .Z(n369) );
  XOR2_X1 U354 ( .A(KEYINPUT78), .B(G162GAT), .Z(n363) );
  XNOR2_X1 U355 ( .A(n369), .B(n363), .ZN(n298) );
  XNOR2_X1 U356 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U357 ( .A(n300), .B(KEYINPUT22), .Z(n307) );
  XOR2_X1 U358 ( .A(G155GAT), .B(KEYINPUT91), .Z(n302) );
  XNOR2_X1 U359 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n428) );
  XOR2_X1 U361 ( .A(KEYINPUT89), .B(n428), .Z(n304) );
  NAND2_X1 U362 ( .A1(G228GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U363 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U364 ( .A(G50GAT), .B(n305), .ZN(n306) );
  XNOR2_X1 U365 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n492) );
  INV_X1 U367 ( .A(n544), .ZN(n475) );
  XOR2_X1 U368 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n311) );
  XNOR2_X1 U369 ( .A(KEYINPUT88), .B(G183GAT), .ZN(n310) );
  XNOR2_X1 U370 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U371 ( .A(KEYINPUT17), .B(n312), .Z(n447) );
  XOR2_X1 U372 ( .A(KEYINPUT87), .B(G176GAT), .Z(n314) );
  NAND2_X1 U373 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U374 ( .A(n314), .B(n313), .ZN(n317) );
  XNOR2_X1 U375 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n315), .B(G127GAT), .ZN(n429) );
  INV_X1 U377 ( .A(n429), .ZN(n316) );
  XOR2_X1 U378 ( .A(G190GAT), .B(G134GAT), .Z(n353) );
  XOR2_X1 U379 ( .A(G120GAT), .B(G71GAT), .Z(n395) );
  XNOR2_X1 U380 ( .A(n353), .B(n395), .ZN(n318) );
  XOR2_X1 U381 ( .A(KEYINPUT20), .B(G99GAT), .Z(n321) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(G15GAT), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U384 ( .A(G169GAT), .B(n322), .ZN(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U386 ( .A(KEYINPUT84), .B(KEYINPUT81), .Z(n327) );
  XNOR2_X1 U387 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n332) );
  XNOR2_X1 U389 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n328), .B(KEYINPUT13), .ZN(n392) );
  XOR2_X1 U391 ( .A(n392), .B(G71GAT), .Z(n330) );
  XNOR2_X1 U392 ( .A(n371), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U395 ( .A(G155GAT), .B(G78GAT), .Z(n334) );
  XNOR2_X1 U396 ( .A(G22GAT), .B(G127GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U398 ( .A(KEYINPUT83), .B(G64GAT), .Z(n336) );
  XNOR2_X1 U399 ( .A(G8GAT), .B(G211GAT), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U401 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U402 ( .A(KEYINPUT85), .B(KEYINPUT82), .Z(n340) );
  NAND2_X1 U403 ( .A1(G231GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U405 ( .A(KEYINPUT15), .B(n341), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U407 ( .A(n345), .B(n344), .Z(n582) );
  INV_X1 U408 ( .A(n582), .ZN(n479) );
  XNOR2_X1 U409 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n346), .B(G29GAT), .ZN(n347) );
  XOR2_X1 U411 ( .A(n347), .B(KEYINPUT8), .Z(n349) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(G50GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n349), .B(n348), .ZN(n380) );
  XOR2_X1 U414 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n351) );
  XNOR2_X1 U415 ( .A(G218GAT), .B(KEYINPUT79), .ZN(n350) );
  XNOR2_X1 U416 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U417 ( .A(n352), .B(KEYINPUT80), .Z(n355) );
  XNOR2_X1 U418 ( .A(n353), .B(G106GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U420 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n357) );
  NAND2_X1 U421 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U422 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U423 ( .A(n359), .B(n358), .Z(n365) );
  XOR2_X1 U424 ( .A(KEYINPUT74), .B(G92GAT), .Z(n361) );
  XNOR2_X1 U425 ( .A(G99GAT), .B(KEYINPUT75), .ZN(n360) );
  XNOR2_X1 U426 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U427 ( .A(G85GAT), .B(n362), .Z(n381) );
  XNOR2_X1 U428 ( .A(n363), .B(n381), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(n380), .B(n366), .Z(n499) );
  INV_X1 U431 ( .A(n499), .ZN(n568) );
  XOR2_X1 U432 ( .A(KEYINPUT46), .B(KEYINPUT114), .Z(n401) );
  XOR2_X1 U433 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n368) );
  XNOR2_X1 U434 ( .A(KEYINPUT66), .B(KEYINPUT67), .ZN(n367) );
  XNOR2_X1 U435 ( .A(n368), .B(n367), .ZN(n370) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U437 ( .A(n371), .B(KEYINPUT30), .Z(n373) );
  NAND2_X1 U438 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U439 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U440 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U441 ( .A(G169GAT), .B(G8GAT), .Z(n438) );
  XOR2_X1 U442 ( .A(n376), .B(n438), .Z(n378) );
  XNOR2_X1 U443 ( .A(G113GAT), .B(G197GAT), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X2 U445 ( .A(n380), .B(n379), .Z(n575) );
  XNOR2_X1 U446 ( .A(n382), .B(n381), .ZN(n399) );
  INV_X1 U447 ( .A(KEYINPUT33), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n383), .A2(KEYINPUT71), .ZN(n386) );
  INV_X1 U449 ( .A(KEYINPUT71), .ZN(n384) );
  NAND2_X1 U450 ( .A1(n384), .A2(KEYINPUT33), .ZN(n385) );
  NAND2_X1 U451 ( .A1(n386), .A2(n385), .ZN(n388) );
  XNOR2_X1 U452 ( .A(KEYINPUT31), .B(KEYINPUT77), .ZN(n387) );
  XNOR2_X1 U453 ( .A(n388), .B(n387), .ZN(n391) );
  AND2_X1 U454 ( .A1(G230GAT), .A2(G233GAT), .ZN(n389) );
  XOR2_X1 U455 ( .A(n393), .B(n392), .Z(n397) );
  XNOR2_X1 U456 ( .A(G176GAT), .B(G64GAT), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n394), .B(KEYINPUT76), .ZN(n439) );
  XNOR2_X1 U458 ( .A(n395), .B(n439), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U460 ( .A(KEYINPUT41), .B(n578), .ZN(n522) );
  INV_X1 U461 ( .A(n522), .ZN(n555) );
  NAND2_X1 U462 ( .A1(n575), .A2(n555), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  NOR2_X1 U464 ( .A1(n568), .A2(n402), .ZN(n403) );
  NAND2_X1 U465 ( .A1(n479), .A2(n403), .ZN(n404) );
  XNOR2_X1 U466 ( .A(KEYINPUT47), .B(n404), .ZN(n405) );
  XNOR2_X1 U467 ( .A(n405), .B(KEYINPUT115), .ZN(n410) );
  XOR2_X1 U468 ( .A(n568), .B(KEYINPUT36), .Z(n586) );
  NOR2_X1 U469 ( .A1(n479), .A2(n586), .ZN(n406) );
  XOR2_X1 U470 ( .A(KEYINPUT45), .B(n406), .Z(n407) );
  NOR2_X1 U471 ( .A1(n578), .A2(n407), .ZN(n408) );
  XOR2_X1 U472 ( .A(KEYINPUT69), .B(n575), .Z(n563) );
  INV_X1 U473 ( .A(n563), .ZN(n483) );
  NAND2_X1 U474 ( .A1(n408), .A2(n483), .ZN(n409) );
  NAND2_X1 U475 ( .A1(n410), .A2(n409), .ZN(n412) );
  XOR2_X1 U476 ( .A(KEYINPUT116), .B(KEYINPUT48), .Z(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n488) );
  XOR2_X1 U478 ( .A(G85GAT), .B(G162GAT), .Z(n414) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(G134GAT), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n418) );
  XOR2_X1 U481 ( .A(G57GAT), .B(G148GAT), .Z(n416) );
  XNOR2_X1 U482 ( .A(G141GAT), .B(G120GAT), .ZN(n415) );
  XNOR2_X1 U483 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U484 ( .A(n418), .B(n417), .Z(n423) );
  XOR2_X1 U485 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n420) );
  NAND2_X1 U486 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U487 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U488 ( .A(KEYINPUT1), .B(n421), .ZN(n422) );
  XNOR2_X1 U489 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U490 ( .A(KEYINPUT6), .B(KEYINPUT92), .Z(n425) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U493 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U495 ( .A(n431), .B(n430), .ZN(n536) );
  XOR2_X1 U496 ( .A(G92GAT), .B(G204GAT), .Z(n433) );
  XNOR2_X1 U497 ( .A(G36GAT), .B(G190GAT), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U499 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n435) );
  XNOR2_X1 U500 ( .A(KEYINPUT94), .B(KEYINPUT95), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U502 ( .A(n437), .B(n436), .Z(n445) );
  XOR2_X1 U503 ( .A(n439), .B(n438), .Z(n441) );
  NAND2_X1 U504 ( .A1(G226GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U507 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U508 ( .A(n447), .B(n446), .ZN(n538) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n538), .ZN(n466) );
  NOR2_X1 U510 ( .A1(n536), .A2(n466), .ZN(n473) );
  INV_X1 U511 ( .A(n473), .ZN(n448) );
  NOR2_X1 U512 ( .A1(n488), .A2(n448), .ZN(n449) );
  XNOR2_X1 U513 ( .A(n449), .B(KEYINPUT117), .ZN(n552) );
  NOR2_X1 U514 ( .A1(n540), .A2(n552), .ZN(n450) );
  XOR2_X1 U515 ( .A(KEYINPUT118), .B(n450), .Z(n451) );
  NAND2_X1 U516 ( .A1(n548), .A2(n555), .ZN(n455) );
  XOR2_X1 U517 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n453) );
  INV_X1 U518 ( .A(G120GAT), .ZN(n452) );
  XNOR2_X1 U519 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U520 ( .A(n455), .B(n454), .ZN(G1341GAT) );
  NAND2_X1 U521 ( .A1(n548), .A2(n582), .ZN(n459) );
  XOR2_X1 U522 ( .A(KEYINPUT50), .B(KEYINPUT120), .Z(n457) );
  INV_X1 U523 ( .A(G127GAT), .ZN(n456) );
  XNOR2_X1 U524 ( .A(n459), .B(n458), .ZN(G1342GAT) );
  NOR2_X1 U525 ( .A1(n540), .A2(n538), .ZN(n460) );
  NOR2_X1 U526 ( .A1(n492), .A2(n460), .ZN(n463) );
  XNOR2_X1 U527 ( .A(KEYINPUT25), .B(KEYINPUT102), .ZN(n461) );
  XNOR2_X1 U528 ( .A(n461), .B(KEYINPUT101), .ZN(n462) );
  XNOR2_X1 U529 ( .A(n463), .B(n462), .ZN(n469) );
  XOR2_X1 U530 ( .A(KEYINPUT99), .B(KEYINPUT26), .Z(n465) );
  NAND2_X1 U531 ( .A1(n492), .A2(n540), .ZN(n464) );
  XNOR2_X1 U532 ( .A(n465), .B(n464), .ZN(n573) );
  NOR2_X1 U533 ( .A1(n466), .A2(n573), .ZN(n467) );
  XNOR2_X1 U534 ( .A(KEYINPUT100), .B(n467), .ZN(n468) );
  XNOR2_X1 U535 ( .A(KEYINPUT103), .B(n470), .ZN(n471) );
  NAND2_X1 U536 ( .A1(n471), .A2(n536), .ZN(n472) );
  XOR2_X1 U537 ( .A(KEYINPUT104), .B(n472), .Z(n478) );
  NAND2_X1 U538 ( .A1(n473), .A2(n540), .ZN(n474) );
  NOR2_X1 U539 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U540 ( .A(n476), .B(KEYINPUT98), .ZN(n477) );
  NOR2_X1 U541 ( .A1(n478), .A2(n477), .ZN(n503) );
  OR2_X1 U542 ( .A1(n503), .A2(n481), .ZN(n482) );
  XNOR2_X1 U543 ( .A(KEYINPUT37), .B(n482), .ZN(n535) );
  NOR2_X1 U544 ( .A1(n483), .A2(n578), .ZN(n505) );
  NAND2_X1 U545 ( .A1(n535), .A2(n505), .ZN(n484) );
  NOR2_X1 U546 ( .A1(n520), .A2(n538), .ZN(n487) );
  NOR2_X1 U547 ( .A1(n488), .A2(n538), .ZN(n489) );
  XNOR2_X1 U548 ( .A(n489), .B(KEYINPUT54), .ZN(n490) );
  NAND2_X1 U549 ( .A1(n490), .A2(n536), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n491), .B(KEYINPUT64), .ZN(n574) );
  NOR2_X1 U551 ( .A1(n492), .A2(n574), .ZN(n493) );
  XNOR2_X1 U552 ( .A(n493), .B(KEYINPUT55), .ZN(n494) );
  NOR2_X2 U553 ( .A1(n540), .A2(n494), .ZN(n567) );
  NAND2_X1 U554 ( .A1(n567), .A2(n555), .ZN(n498) );
  XOR2_X1 U555 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n496) );
  XNOR2_X1 U556 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n495) );
  NAND2_X1 U557 ( .A1(n582), .A2(n499), .ZN(n500) );
  XNOR2_X1 U558 ( .A(n500), .B(KEYINPUT16), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(KEYINPUT86), .ZN(n502) );
  NOR2_X1 U560 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U561 ( .A(KEYINPUT105), .B(n504), .Z(n523) );
  NAND2_X1 U562 ( .A1(n505), .A2(n523), .ZN(n512) );
  NOR2_X1 U563 ( .A1(n536), .A2(n512), .ZN(n507) );
  XNOR2_X1 U564 ( .A(KEYINPUT34), .B(KEYINPUT106), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U566 ( .A(G1GAT), .B(n508), .Z(G1324GAT) );
  NOR2_X1 U567 ( .A1(n538), .A2(n512), .ZN(n509) );
  XOR2_X1 U568 ( .A(G8GAT), .B(n509), .Z(G1325GAT) );
  NOR2_X1 U569 ( .A1(n540), .A2(n512), .ZN(n511) );
  XNOR2_X1 U570 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  NOR2_X1 U572 ( .A1(n544), .A2(n512), .ZN(n513) );
  XOR2_X1 U573 ( .A(G22GAT), .B(n513), .Z(G1327GAT) );
  NOR2_X1 U574 ( .A1(n536), .A2(n520), .ZN(n516) );
  XOR2_X1 U575 ( .A(G29GAT), .B(KEYINPUT107), .Z(n514) );
  XNOR2_X1 U576 ( .A(KEYINPUT39), .B(n514), .ZN(n515) );
  XNOR2_X1 U577 ( .A(n516), .B(n515), .ZN(G1328GAT) );
  NOR2_X1 U578 ( .A1(n520), .A2(n540), .ZN(n518) );
  XNOR2_X1 U579 ( .A(KEYINPUT40), .B(KEYINPUT109), .ZN(n517) );
  XNOR2_X1 U580 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U581 ( .A(G43GAT), .B(n519), .ZN(G1330GAT) );
  NOR2_X1 U582 ( .A1(n544), .A2(n520), .ZN(n521) );
  XOR2_X1 U583 ( .A(G50GAT), .B(n521), .Z(G1331GAT) );
  NOR2_X1 U584 ( .A1(n575), .A2(n522), .ZN(n534) );
  NAND2_X1 U585 ( .A1(n523), .A2(n534), .ZN(n529) );
  NOR2_X1 U586 ( .A1(n536), .A2(n529), .ZN(n524) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n524), .Z(n525) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(n525), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n538), .A2(n529), .ZN(n526) );
  XOR2_X1 U590 ( .A(KEYINPUT110), .B(n526), .Z(n527) );
  XNOR2_X1 U591 ( .A(G64GAT), .B(n527), .ZN(G1333GAT) );
  NOR2_X1 U592 ( .A1(n540), .A2(n529), .ZN(n528) );
  XOR2_X1 U593 ( .A(G71GAT), .B(n528), .Z(G1334GAT) );
  NOR2_X1 U594 ( .A1(n529), .A2(n544), .ZN(n533) );
  XOR2_X1 U595 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n531) );
  XNOR2_X1 U596 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1335GAT) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n543) );
  NOR2_X1 U600 ( .A1(n536), .A2(n543), .ZN(n537) );
  XOR2_X1 U601 ( .A(G85GAT), .B(n537), .Z(G1336GAT) );
  NOR2_X1 U602 ( .A1(n538), .A2(n543), .ZN(n539) );
  XOR2_X1 U603 ( .A(G92GAT), .B(n539), .Z(G1337GAT) );
  NOR2_X1 U604 ( .A1(n540), .A2(n543), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1338GAT) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U608 ( .A(KEYINPUT44), .B(n545), .Z(n546) );
  XNOR2_X1 U609 ( .A(G106GAT), .B(n546), .ZN(G1339GAT) );
  NAND2_X1 U610 ( .A1(n563), .A2(n548), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G113GAT), .B(n547), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT121), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U613 ( .A1(n548), .A2(n568), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U615 ( .A(G134GAT), .B(n551), .Z(G1343GAT) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(KEYINPUT122), .ZN(n554) );
  NOR2_X1 U617 ( .A1(n573), .A2(n552), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n575), .A2(n560), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U621 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n582), .A2(n560), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U626 ( .A(G162GAT), .B(KEYINPUT123), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n568), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n567), .ZN(n564) );
  XNOR2_X1 U630 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT125), .Z(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n582), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT60), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(n572), .Z(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n584) );
  NAND2_X1 U641 ( .A1(n584), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n580) );
  NAND2_X1 U644 ( .A1(n584), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U646 ( .A(G204GAT), .B(n581), .Z(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U649 ( .A(KEYINPUT62), .ZN(n588) );
  INV_X1 U650 ( .A(n584), .ZN(n585) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

