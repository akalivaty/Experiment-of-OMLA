

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775;

  XNOR2_X1 U365 ( .A(n574), .B(n387), .ZN(n708) );
  INV_X1 U366 ( .A(G116), .ZN(n504) );
  XNOR2_X2 U367 ( .A(n543), .B(KEYINPUT16), .ZN(n430) );
  XNOR2_X2 U368 ( .A(n512), .B(n511), .ZN(n543) );
  INV_X1 U369 ( .A(n343), .ZN(n345) );
  NAND2_X1 U370 ( .A1(n436), .A2(n435), .ZN(n343) );
  XNOR2_X2 U371 ( .A(n386), .B(n555), .ZN(n712) );
  INV_X1 U372 ( .A(G953), .ZN(n762) );
  AND2_X2 U373 ( .A1(n408), .A2(n355), .ZN(n419) );
  NAND2_X2 U374 ( .A1(n612), .A2(n606), .ZN(n607) );
  XNOR2_X2 U375 ( .A(KEYINPUT69), .B(G119), .ZN(n508) );
  XNOR2_X2 U376 ( .A(n431), .B(G143), .ZN(n492) );
  XNOR2_X2 U377 ( .A(G128), .B(KEYINPUT79), .ZN(n431) );
  XNOR2_X2 U378 ( .A(KEYINPUT3), .B(G113), .ZN(n510) );
  INV_X1 U379 ( .A(n695), .ZN(n402) );
  NOR2_X1 U380 ( .A1(G953), .A2(G237), .ZN(n513) );
  NAND2_X1 U381 ( .A1(n426), .A2(n679), .ZN(n733) );
  INV_X1 U382 ( .A(n672), .ZN(n670) );
  NOR2_X1 U383 ( .A1(n682), .A2(n632), .ZN(n425) );
  XNOR2_X1 U384 ( .A(n760), .B(G146), .ZN(n521) );
  XOR2_X1 U385 ( .A(G146), .B(G125), .Z(n537) );
  BUF_X1 U386 ( .A(n740), .Z(n745) );
  NAND2_X1 U387 ( .A1(n750), .A2(n425), .ZN(n424) );
  AND2_X1 U388 ( .A1(n394), .A2(n393), .ZN(n392) );
  NOR2_X1 U389 ( .A1(n642), .A2(n396), .ZN(n390) );
  XNOR2_X1 U390 ( .A(n578), .B(n577), .ZN(n772) );
  AND2_X1 U391 ( .A1(n374), .A2(n372), .ZN(n371) );
  XNOR2_X1 U392 ( .A(n473), .B(KEYINPUT104), .ZN(n672) );
  XNOR2_X1 U393 ( .A(n541), .B(n493), .ZN(n760) );
  XNOR2_X1 U394 ( .A(n507), .B(n508), .ZN(n512) );
  XNOR2_X1 U395 ( .A(n492), .B(KEYINPUT4), .ZN(n541) );
  XNOR2_X1 U396 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U397 ( .A(n494), .B(G107), .ZN(n542) );
  XNOR2_X1 U398 ( .A(n537), .B(n404), .ZN(n479) );
  XNOR2_X1 U399 ( .A(G104), .B(G110), .ZN(n494) );
  NAND2_X1 U400 ( .A1(n356), .A2(n588), .ZN(n682) );
  AND2_X1 U401 ( .A1(n609), .A2(n616), .ZN(n610) );
  XNOR2_X2 U402 ( .A(n576), .B(n575), .ZN(n616) );
  NOR2_X1 U403 ( .A1(G902), .A2(G237), .ZN(n526) );
  XNOR2_X1 U404 ( .A(n409), .B(KEYINPUT83), .ZN(n579) );
  NAND2_X1 U405 ( .A1(n773), .A2(n608), .ZN(n395) );
  INV_X1 U406 ( .A(KEYINPUT38), .ZN(n387) );
  AND2_X1 U407 ( .A1(n670), .A2(n568), .ZN(n570) );
  XNOR2_X1 U408 ( .A(n569), .B(KEYINPUT105), .ZN(n599) );
  NAND2_X1 U409 ( .A1(n434), .A2(n433), .ZN(n432) );
  NOR2_X1 U410 ( .A1(n774), .A2(n437), .ZN(n433) );
  AND2_X1 U411 ( .A1(n442), .A2(n441), .ZN(n440) );
  NAND2_X1 U412 ( .A1(n581), .A2(n443), .ZN(n441) );
  NAND2_X1 U413 ( .A1(n391), .A2(n390), .ZN(n389) );
  XNOR2_X1 U414 ( .A(G128), .B(KEYINPUT23), .ZN(n480) );
  XNOR2_X1 U415 ( .A(n479), .B(n478), .ZN(n759) );
  XNOR2_X1 U416 ( .A(G902), .B(KEYINPUT15), .ZN(n631) );
  XNOR2_X1 U417 ( .A(n357), .B(n444), .ZN(n356) );
  OR2_X1 U418 ( .A1(n635), .A2(G902), .ZN(n525) );
  XNOR2_X1 U419 ( .A(n560), .B(n353), .ZN(n593) );
  NAND2_X1 U420 ( .A1(n403), .A2(n459), .ZN(n552) );
  OR2_X1 U421 ( .A1(n736), .A2(n378), .ZN(n377) );
  AND2_X1 U422 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U423 ( .A1(G469), .A2(n459), .ZN(n378) );
  XOR2_X1 U424 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n454) );
  XNOR2_X1 U425 ( .A(n399), .B(n549), .ZN(n583) );
  NAND2_X1 U426 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U427 ( .A1(n366), .A2(n349), .ZN(n361) );
  AND2_X1 U428 ( .A1(n365), .A2(n364), .ZN(n363) );
  NOR2_X1 U429 ( .A1(n619), .A2(n350), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n598), .B(KEYINPUT22), .ZN(n604) );
  XNOR2_X1 U431 ( .A(n460), .B(G478), .ZN(n564) );
  INV_X1 U432 ( .A(KEYINPUT44), .ZN(n396) );
  INV_X1 U433 ( .A(KEYINPUT68), .ZN(n443) );
  INV_X1 U434 ( .A(KEYINPUT91), .ZN(n509) );
  NAND2_X1 U435 ( .A1(n506), .A2(n505), .ZN(n507) );
  NAND2_X1 U436 ( .A1(n359), .A2(n358), .ZN(n357) );
  NAND2_X1 U437 ( .A1(n345), .A2(n432), .ZN(n358) );
  NAND2_X1 U438 ( .A1(n439), .A2(n344), .ZN(n438) );
  INV_X1 U439 ( .A(KEYINPUT48), .ZN(n444) );
  NAND2_X1 U440 ( .A1(n732), .A2(G902), .ZN(n380) );
  XNOR2_X1 U441 ( .A(G134), .B(G131), .ZN(n493) );
  XOR2_X1 U442 ( .A(G137), .B(G140), .Z(n495) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n529) );
  INV_X1 U444 ( .A(KEYINPUT109), .ZN(n555) );
  NAND2_X1 U445 ( .A1(n708), .A2(n707), .ZN(n386) );
  NAND2_X1 U446 ( .A1(n571), .A2(n574), .ZN(n366) );
  OR2_X1 U447 ( .A1(n695), .A2(n694), .ZN(n691) );
  INV_X1 U448 ( .A(KEYINPUT6), .ZN(n405) );
  XNOR2_X1 U449 ( .A(n481), .B(n412), .ZN(n483) );
  XNOR2_X1 U450 ( .A(n480), .B(n413), .ZN(n412) );
  INV_X1 U451 ( .A(KEYINPUT95), .ZN(n413) );
  XNOR2_X1 U452 ( .A(G119), .B(G110), .ZN(n482) );
  INV_X1 U453 ( .A(KEYINPUT10), .ZN(n404) );
  XOR2_X1 U454 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n462) );
  NAND2_X1 U455 ( .A1(n427), .A2(n632), .ZN(n418) );
  NAND2_X1 U456 ( .A1(n631), .A2(KEYINPUT64), .ZN(n422) );
  NAND2_X1 U457 ( .A1(n428), .A2(n421), .ZN(n420) );
  NAND2_X1 U458 ( .A1(KEYINPUT64), .A2(KEYINPUT2), .ZN(n421) );
  INV_X1 U459 ( .A(KEYINPUT75), .ZN(n423) );
  AND2_X1 U460 ( .A1(n373), .A2(n406), .ZN(n372) );
  INV_X1 U461 ( .A(n611), .ZN(n406) );
  XOR2_X1 U462 ( .A(KEYINPUT108), .B(KEYINPUT30), .Z(n528) );
  AND2_X1 U463 ( .A1(n593), .A2(n554), .ZN(n561) );
  XNOR2_X1 U464 ( .A(n384), .B(n383), .ZN(n562) );
  INV_X1 U465 ( .A(KEYINPUT28), .ZN(n383) );
  AND2_X1 U466 ( .A1(n571), .A2(n557), .ZN(n385) );
  XNOR2_X1 U467 ( .A(n470), .B(n415), .ZN(n563) );
  XNOR2_X1 U468 ( .A(n471), .B(n651), .ZN(n415) );
  NAND2_X1 U469 ( .A1(n593), .A2(n450), .ZN(n429) );
  INV_X1 U470 ( .A(KEYINPUT97), .ZN(n501) );
  NAND2_X1 U471 ( .A1(n402), .A2(n401), .ZN(n400) );
  XNOR2_X1 U472 ( .A(n411), .B(n455), .ZN(n458) );
  XNOR2_X1 U473 ( .A(n457), .B(n456), .ZN(n411) );
  INV_X1 U474 ( .A(KEYINPUT40), .ZN(n550) );
  INV_X1 U475 ( .A(KEYINPUT111), .ZN(n577) );
  AND2_X1 U476 ( .A1(n562), .A2(n561), .ZN(n669) );
  NOR2_X1 U477 ( .A1(n604), .A2(n600), .ZN(n602) );
  XNOR2_X1 U478 ( .A(n608), .B(G110), .ZN(G12) );
  NOR2_X1 U479 ( .A1(n581), .A2(n443), .ZN(n344) );
  INV_X1 U480 ( .A(KEYINPUT64), .ZN(n427) );
  INV_X1 U481 ( .A(n694), .ZN(n401) );
  NOR2_X1 U482 ( .A1(n573), .A2(n572), .ZN(n346) );
  AND2_X1 U483 ( .A1(n407), .A2(n620), .ZN(n347) );
  NAND2_X2 U484 ( .A1(n379), .A2(n377), .ZN(n576) );
  INV_X1 U485 ( .A(G902), .ZN(n459) );
  AND2_X1 U486 ( .A1(n711), .A2(n561), .ZN(n348) );
  XOR2_X1 U487 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n349) );
  XNOR2_X1 U488 ( .A(KEYINPUT70), .B(KEYINPUT34), .ZN(n350) );
  XOR2_X1 U489 ( .A(n594), .B(KEYINPUT0), .Z(n351) );
  XNOR2_X1 U490 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n352) );
  XOR2_X1 U491 ( .A(n559), .B(KEYINPUT19), .Z(n353) );
  AND2_X1 U492 ( .A1(n428), .A2(KEYINPUT64), .ZN(n354) );
  NAND2_X1 U493 ( .A1(n422), .A2(n420), .ZN(n355) );
  NAND2_X1 U494 ( .A1(n440), .A2(n438), .ZN(n359) );
  NAND2_X1 U495 ( .A1(n363), .A2(n360), .ZN(n367) );
  INV_X1 U496 ( .A(n573), .ZN(n362) );
  NAND2_X1 U497 ( .A1(n366), .A2(n349), .ZN(n364) );
  NAND2_X1 U498 ( .A1(n573), .A2(n349), .ZN(n365) );
  NAND2_X1 U499 ( .A1(n367), .A2(n616), .ZN(n578) );
  INV_X1 U500 ( .A(n574), .ZN(n368) );
  NAND2_X1 U501 ( .A1(n407), .A2(n369), .ZN(n399) );
  AND2_X1 U502 ( .A1(n548), .A2(n620), .ZN(n369) );
  NAND2_X1 U503 ( .A1(n347), .A2(n445), .ZN(n668) );
  NAND2_X1 U504 ( .A1(n371), .A2(n370), .ZN(n397) );
  NAND2_X1 U505 ( .A1(n718), .A2(n350), .ZN(n370) );
  NAND2_X1 U506 ( .A1(n619), .A2(n350), .ZN(n373) );
  NAND2_X1 U507 ( .A1(n376), .A2(n375), .ZN(n374) );
  INV_X1 U508 ( .A(n718), .ZN(n376) );
  XNOR2_X2 U509 ( .A(n410), .B(n352), .ZN(n718) );
  NAND2_X1 U510 ( .A1(n736), .A2(n732), .ZN(n381) );
  NAND2_X1 U511 ( .A1(n570), .A2(n382), .ZN(n573) );
  NAND2_X1 U512 ( .A1(n610), .A2(n382), .ZN(n410) );
  NOR2_X2 U513 ( .A1(n604), .A2(n382), .ZN(n612) );
  XNOR2_X2 U514 ( .A(n621), .B(n405), .ZN(n382) );
  NAND2_X1 U515 ( .A1(n348), .A2(n562), .ZN(n580) );
  NAND2_X1 U516 ( .A1(n599), .A2(n385), .ZN(n384) );
  XNOR2_X2 U517 ( .A(n388), .B(n545), .ZN(n645) );
  XNOR2_X1 U518 ( .A(n388), .B(KEYINPUT125), .ZN(n756) );
  XNOR2_X2 U519 ( .A(n430), .B(n544), .ZN(n388) );
  NAND2_X1 U520 ( .A1(n603), .A2(n695), .ZN(n608) );
  XNOR2_X2 U521 ( .A(n607), .B(KEYINPUT32), .ZN(n773) );
  NAND2_X1 U522 ( .A1(n392), .A2(n389), .ZN(n627) );
  INV_X1 U523 ( .A(n395), .ZN(n391) );
  NAND2_X1 U524 ( .A1(n395), .A2(n396), .ZN(n393) );
  NAND2_X1 U525 ( .A1(n642), .A2(n396), .ZN(n394) );
  XNOR2_X2 U526 ( .A(n397), .B(KEYINPUT35), .ZN(n642) );
  XNOR2_X2 U527 ( .A(n398), .B(KEYINPUT42), .ZN(n775) );
  NOR2_X2 U528 ( .A1(n706), .A2(n556), .ZN(n398) );
  NOR2_X1 U529 ( .A1(n400), .A2(n576), .ZN(n502) );
  INV_X1 U530 ( .A(n746), .ZN(n403) );
  XNOR2_X1 U531 ( .A(n527), .B(n528), .ZN(n407) );
  NAND2_X1 U532 ( .A1(n630), .A2(n354), .ZN(n408) );
  NAND2_X1 U533 ( .A1(n583), .A2(n670), .ZN(n551) );
  NAND2_X1 U534 ( .A1(n447), .A2(n668), .ZN(n409) );
  NAND2_X1 U535 ( .A1(n419), .A2(n417), .ZN(n426) );
  NOR2_X2 U536 ( .A1(n680), .A2(n682), .ZN(n630) );
  XNOR2_X2 U537 ( .A(n629), .B(n628), .ZN(n680) );
  NAND2_X1 U538 ( .A1(n774), .A2(n437), .ZN(n435) );
  XNOR2_X2 U539 ( .A(n551), .B(n550), .ZN(n774) );
  XNOR2_X1 U540 ( .A(n488), .B(n487), .ZN(n746) );
  NAND2_X1 U541 ( .A1(n775), .A2(n437), .ZN(n436) );
  XNOR2_X2 U542 ( .A(n414), .B(KEYINPUT41), .ZN(n706) );
  NOR2_X2 U543 ( .A1(n712), .A2(n710), .ZN(n414) );
  XNOR2_X1 U544 ( .A(n416), .B(n469), .ZN(n653) );
  XNOR2_X1 U545 ( .A(n479), .B(n449), .ZN(n416) );
  NAND2_X1 U546 ( .A1(n582), .A2(n443), .ZN(n442) );
  OR2_X1 U547 ( .A1(n630), .A2(n418), .ZN(n417) );
  XNOR2_X2 U548 ( .A(n424), .B(n423), .ZN(n679) );
  INV_X1 U549 ( .A(n680), .ZN(n750) );
  INV_X1 U550 ( .A(n631), .ZN(n428) );
  INV_X1 U551 ( .A(n597), .ZN(n619) );
  NAND2_X1 U552 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X2 U553 ( .A(n429), .B(n351), .ZN(n597) );
  XNOR2_X2 U554 ( .A(n525), .B(n524), .ZN(n569) );
  INV_X1 U555 ( .A(n775), .ZN(n434) );
  INV_X1 U556 ( .A(KEYINPUT46), .ZN(n437) );
  INV_X1 U557 ( .A(n582), .ZN(n439) );
  NAND2_X1 U558 ( .A1(n580), .A2(KEYINPUT47), .ZN(n447) );
  NOR2_X1 U559 ( .A1(n446), .A2(n611), .ZN(n445) );
  NAND2_X1 U560 ( .A1(n574), .A2(n557), .ZN(n446) );
  XNOR2_X1 U561 ( .A(n468), .B(n467), .ZN(n469) );
  AND2_X1 U562 ( .A1(G210), .A2(n546), .ZN(n448) );
  XOR2_X1 U563 ( .A(n462), .B(n461), .Z(n449) );
  OR2_X1 U564 ( .A1(n592), .A2(n591), .ZN(n450) );
  INV_X1 U565 ( .A(n495), .ZN(n478) );
  XNOR2_X1 U566 ( .A(n539), .B(n538), .ZN(n540) );
  AND2_X1 U567 ( .A1(n595), .A2(n401), .ZN(n596) );
  XNOR2_X1 U568 ( .A(n485), .B(n484), .ZN(n488) );
  INV_X1 U569 ( .A(KEYINPUT63), .ZN(n640) );
  XOR2_X1 U570 ( .A(KEYINPUT7), .B(G107), .Z(n452) );
  XNOR2_X1 U571 ( .A(G116), .B(G122), .ZN(n451) );
  XNOR2_X1 U572 ( .A(n452), .B(n451), .ZN(n457) );
  XOR2_X1 U573 ( .A(G134), .B(KEYINPUT9), .Z(n456) );
  NAND2_X1 U574 ( .A1(G234), .A2(n762), .ZN(n453) );
  XNOR2_X1 U575 ( .A(n454), .B(n453), .ZN(n486) );
  NAND2_X1 U576 ( .A1(G217), .A2(n486), .ZN(n455) );
  XNOR2_X1 U577 ( .A(n492), .B(n458), .ZN(n741) );
  NAND2_X1 U578 ( .A1(n741), .A2(n459), .ZN(n460) );
  INV_X1 U579 ( .A(n564), .ZN(n472) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(KEYINPUT103), .ZN(n471) );
  NAND2_X1 U581 ( .A1(G214), .A2(n513), .ZN(n461) );
  XOR2_X1 U582 ( .A(G104), .B(G122), .Z(n464) );
  XNOR2_X1 U583 ( .A(G113), .B(G143), .ZN(n463) );
  XNOR2_X1 U584 ( .A(n464), .B(n463), .ZN(n468) );
  XOR2_X1 U585 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n466) );
  XNOR2_X1 U586 ( .A(G131), .B(G140), .ZN(n465) );
  XNOR2_X1 U587 ( .A(n466), .B(n465), .ZN(n467) );
  NOR2_X1 U588 ( .A1(G902), .A2(n653), .ZN(n470) );
  INV_X1 U589 ( .A(G475), .ZN(n651) );
  NAND2_X1 U590 ( .A1(n472), .A2(n563), .ZN(n473) );
  XOR2_X1 U591 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n476) );
  NAND2_X1 U592 ( .A1(G234), .A2(n631), .ZN(n474) );
  XNOR2_X1 U593 ( .A(KEYINPUT20), .B(n474), .ZN(n489) );
  NAND2_X1 U594 ( .A1(G217), .A2(n489), .ZN(n475) );
  XNOR2_X1 U595 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U596 ( .A(KEYINPUT25), .B(n477), .ZN(n553) );
  INV_X1 U597 ( .A(n759), .ZN(n485) );
  XOR2_X1 U598 ( .A(KEYINPUT24), .B(KEYINPUT94), .Z(n481) );
  XNOR2_X1 U599 ( .A(n483), .B(n482), .ZN(n484) );
  NAND2_X1 U600 ( .A1(n486), .A2(G221), .ZN(n487) );
  XNOR2_X2 U601 ( .A(n553), .B(n552), .ZN(n695) );
  XOR2_X1 U602 ( .A(KEYINPUT21), .B(KEYINPUT96), .Z(n491) );
  NAND2_X1 U603 ( .A1(n489), .A2(G221), .ZN(n490) );
  XOR2_X1 U604 ( .A(n491), .B(n490), .Z(n694) );
  XNOR2_X1 U605 ( .A(G101), .B(KEYINPUT78), .ZN(n499) );
  XOR2_X1 U606 ( .A(n542), .B(n495), .Z(n497) );
  NAND2_X1 U607 ( .A1(G227), .A2(n762), .ZN(n496) );
  XNOR2_X1 U608 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U609 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U610 ( .A(n521), .B(n500), .ZN(n736) );
  INV_X1 U611 ( .A(G469), .ZN(n732) );
  XNOR2_X1 U612 ( .A(n502), .B(n501), .ZN(n620) );
  INV_X1 U613 ( .A(G101), .ZN(n503) );
  NAND2_X1 U614 ( .A1(n503), .A2(G116), .ZN(n506) );
  NAND2_X1 U615 ( .A1(n504), .A2(G101), .ZN(n505) );
  NAND2_X1 U616 ( .A1(n513), .A2(G210), .ZN(n516) );
  INV_X1 U617 ( .A(KEYINPUT5), .ZN(n514) );
  XNOR2_X1 U618 ( .A(n514), .B(G137), .ZN(n515) );
  XNOR2_X1 U619 ( .A(n516), .B(n515), .ZN(n518) );
  XNOR2_X1 U620 ( .A(KEYINPUT74), .B(KEYINPUT98), .ZN(n517) );
  XNOR2_X1 U621 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U622 ( .A(n543), .B(n519), .ZN(n520) );
  XNOR2_X1 U623 ( .A(n521), .B(n520), .ZN(n635) );
  XNOR2_X1 U624 ( .A(G472), .B(KEYINPUT99), .ZN(n523) );
  INV_X1 U625 ( .A(KEYINPUT71), .ZN(n522) );
  XNOR2_X1 U626 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U627 ( .A(n526), .B(KEYINPUT73), .ZN(n546) );
  NAND2_X1 U628 ( .A1(G214), .A2(n546), .ZN(n707) );
  NAND2_X1 U629 ( .A1(n599), .A2(n707), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n529), .B(KEYINPUT14), .ZN(n530) );
  XNOR2_X1 U631 ( .A(KEYINPUT72), .B(n530), .ZN(n531) );
  NAND2_X1 U632 ( .A1(G952), .A2(n531), .ZN(n725) );
  NOR2_X1 U633 ( .A1(G953), .A2(n725), .ZN(n592) );
  NAND2_X1 U634 ( .A1(G902), .A2(n531), .ZN(n532) );
  XOR2_X1 U635 ( .A(KEYINPUT92), .B(n532), .Z(n533) );
  NAND2_X1 U636 ( .A1(G953), .A2(n533), .ZN(n589) );
  XNOR2_X1 U637 ( .A(KEYINPUT106), .B(n589), .ZN(n534) );
  NOR2_X1 U638 ( .A1(G900), .A2(n534), .ZN(n535) );
  NOR2_X1 U639 ( .A1(n592), .A2(n535), .ZN(n566) );
  INV_X1 U640 ( .A(n566), .ZN(n557) );
  NAND2_X1 U641 ( .A1(G224), .A2(n762), .ZN(n536) );
  XNOR2_X1 U642 ( .A(n537), .B(n536), .ZN(n539) );
  XNOR2_X1 U643 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n538) );
  XNOR2_X1 U644 ( .A(n541), .B(n540), .ZN(n545) );
  XOR2_X1 U645 ( .A(n542), .B(G122), .Z(n544) );
  NAND2_X1 U646 ( .A1(n645), .A2(n631), .ZN(n547) );
  XNOR2_X2 U647 ( .A(n547), .B(n448), .ZN(n558) );
  BUF_X2 U648 ( .A(n558), .Z(n574) );
  AND2_X1 U649 ( .A1(n557), .A2(n708), .ZN(n548) );
  XOR2_X1 U650 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n549) );
  XOR2_X1 U651 ( .A(n553), .B(n552), .Z(n605) );
  NOR2_X1 U652 ( .A1(n605), .A2(n694), .ZN(n571) );
  INV_X1 U653 ( .A(n576), .ZN(n554) );
  NAND2_X1 U654 ( .A1(n562), .A2(n554), .ZN(n556) );
  NOR2_X1 U655 ( .A1(n563), .A2(n564), .ZN(n595) );
  INV_X1 U656 ( .A(n595), .ZN(n710) );
  NAND2_X1 U657 ( .A1(n563), .A2(n564), .ZN(n611) );
  NAND2_X1 U658 ( .A1(n558), .A2(n707), .ZN(n560) );
  INV_X1 U659 ( .A(KEYINPUT66), .ZN(n559) );
  INV_X1 U660 ( .A(n563), .ZN(n565) );
  AND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n664) );
  INV_X1 U662 ( .A(n664), .ZN(n674) );
  NAND2_X1 U663 ( .A1(n672), .A2(n674), .ZN(n711) );
  INV_X1 U664 ( .A(n707), .ZN(n567) );
  NOR2_X1 U665 ( .A1(n567), .A2(n566), .ZN(n568) );
  INV_X1 U666 ( .A(n569), .ZN(n621) );
  INV_X1 U667 ( .A(n571), .ZN(n572) );
  INV_X1 U668 ( .A(KEYINPUT1), .ZN(n575) );
  NAND2_X1 U669 ( .A1(n579), .A2(n772), .ZN(n582) );
  NOR2_X1 U670 ( .A1(KEYINPUT47), .A2(n580), .ZN(n581) );
  NAND2_X1 U671 ( .A1(n583), .A2(n664), .ZN(n677) );
  INV_X1 U672 ( .A(n616), .ZN(n690) );
  NAND2_X1 U673 ( .A1(n690), .A2(n346), .ZN(n584) );
  XNOR2_X1 U674 ( .A(n584), .B(KEYINPUT43), .ZN(n585) );
  NAND2_X1 U675 ( .A1(n585), .A2(n368), .ZN(n586) );
  XNOR2_X1 U676 ( .A(KEYINPUT107), .B(n586), .ZN(n770) );
  INV_X1 U677 ( .A(n770), .ZN(n587) );
  AND2_X1 U678 ( .A1(n677), .A2(n587), .ZN(n588) );
  NOR2_X1 U679 ( .A1(G898), .A2(n589), .ZN(n590) );
  XOR2_X1 U680 ( .A(KEYINPUT93), .B(n590), .Z(n591) );
  INV_X1 U681 ( .A(KEYINPUT67), .ZN(n594) );
  OR2_X1 U682 ( .A1(n616), .A2(n599), .ZN(n600) );
  INV_X1 U683 ( .A(KEYINPUT65), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n602), .B(n601), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n690), .A2(n605), .ZN(n606) );
  INV_X1 U686 ( .A(n691), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n612), .B(KEYINPUT88), .ZN(n614) );
  NOR2_X1 U688 ( .A1(n616), .A2(n695), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n614), .A2(n613), .ZN(n658) );
  NOR2_X1 U690 ( .A1(n569), .A2(n691), .ZN(n615) );
  NAND2_X1 U691 ( .A1(n616), .A2(n615), .ZN(n701) );
  NOR2_X1 U692 ( .A1(n619), .A2(n701), .ZN(n618) );
  XNOR2_X1 U693 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n618), .B(n617), .ZN(n675) );
  INV_X1 U695 ( .A(n620), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n597), .A2(n623), .ZN(n660) );
  NAND2_X1 U698 ( .A1(n675), .A2(n660), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n624), .A2(n711), .ZN(n625) );
  AND2_X1 U700 ( .A1(n658), .A2(n625), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n629) );
  XOR2_X1 U702 ( .A(KEYINPUT86), .B(KEYINPUT45), .Z(n628) );
  INV_X1 U703 ( .A(KEYINPUT2), .ZN(n632) );
  INV_X2 U704 ( .A(n733), .ZN(n740) );
  NAND2_X1 U705 ( .A1(n740), .A2(G472), .ZN(n637) );
  XNOR2_X1 U706 ( .A(KEYINPUT90), .B(KEYINPUT112), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(KEYINPUT62), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U709 ( .A(n637), .B(n636), .ZN(n639) );
  INV_X1 U710 ( .A(G952), .ZN(n638) );
  AND2_X1 U711 ( .A1(n638), .A2(G953), .ZN(n749) );
  NOR2_X2 U712 ( .A1(n639), .A2(n749), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(G57) );
  XOR2_X1 U714 ( .A(n642), .B(G122), .Z(G24) );
  NAND2_X1 U715 ( .A1(n740), .A2(G210), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT81), .B(KEYINPUT54), .Z(n643) );
  XNOR2_X1 U717 ( .A(n643), .B(KEYINPUT55), .ZN(n644) );
  XNOR2_X1 U718 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U719 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U720 ( .A1(n648), .A2(n749), .ZN(n650) );
  XOR2_X1 U721 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n649) );
  XNOR2_X1 U722 ( .A(n650), .B(n649), .ZN(G51) );
  NOR2_X1 U723 ( .A1(n733), .A2(n651), .ZN(n655) );
  XOR2_X1 U724 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n656), .A2(n749), .ZN(n657) );
  XNOR2_X1 U728 ( .A(n657), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U729 ( .A(G101), .B(n658), .ZN(G3) );
  NOR2_X1 U730 ( .A1(n660), .A2(n672), .ZN(n659) );
  XOR2_X1 U731 ( .A(G104), .B(n659), .Z(G6) );
  NOR2_X1 U732 ( .A1(n660), .A2(n674), .ZN(n662) );
  XNOR2_X1 U733 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n661) );
  XNOR2_X1 U734 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(G107), .B(n663), .ZN(G9) );
  XOR2_X1 U736 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n666) );
  NAND2_X1 U737 ( .A1(n669), .A2(n664), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U739 ( .A(G128), .B(n667), .Z(G30) );
  XNOR2_X1 U740 ( .A(G143), .B(n668), .ZN(G45) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U742 ( .A(n671), .B(G146), .ZN(G48) );
  NOR2_X1 U743 ( .A1(n672), .A2(n675), .ZN(n673) );
  XOR2_X1 U744 ( .A(G113), .B(n673), .Z(G15) );
  NOR2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U746 ( .A(G116), .B(n676), .Z(G18) );
  XNOR2_X1 U747 ( .A(G134), .B(n677), .ZN(G36) );
  XOR2_X1 U748 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n731) );
  NOR2_X1 U749 ( .A1(n706), .A2(n718), .ZN(n678) );
  NOR2_X1 U750 ( .A1(n678), .A2(G953), .ZN(n729) );
  INV_X1 U751 ( .A(n679), .ZN(n689) );
  XOR2_X1 U752 ( .A(KEYINPUT2), .B(KEYINPUT82), .Z(n684) );
  NAND2_X1 U753 ( .A1(n680), .A2(n684), .ZN(n681) );
  XOR2_X1 U754 ( .A(KEYINPUT85), .B(n681), .Z(n686) );
  BUF_X1 U755 ( .A(n682), .Z(n683) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U758 ( .A(KEYINPUT80), .B(n687), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n727) );
  NAND2_X1 U760 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n692), .B(KEYINPUT50), .ZN(n693) );
  XNOR2_X1 U762 ( .A(KEYINPUT115), .B(n693), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U764 ( .A(n696), .B(KEYINPUT49), .ZN(n697) );
  XNOR2_X1 U765 ( .A(KEYINPUT114), .B(n697), .ZN(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n700), .A2(n569), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U769 ( .A(n703), .B(KEYINPUT51), .ZN(n704) );
  XNOR2_X1 U770 ( .A(n704), .B(KEYINPUT116), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n706), .A2(n705), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n710), .A2(n709), .ZN(n716) );
  INV_X1 U774 ( .A(n711), .ZN(n713) );
  NOR2_X1 U775 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U776 ( .A(KEYINPUT117), .B(n714), .Z(n715) );
  NOR2_X1 U777 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U778 ( .A(n717), .B(KEYINPUT118), .ZN(n719) );
  NOR2_X1 U779 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U781 ( .A(KEYINPUT119), .B(n722), .Z(n723) );
  XNOR2_X1 U782 ( .A(n723), .B(KEYINPUT52), .ZN(n724) );
  NOR2_X1 U783 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U784 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U786 ( .A(n731), .B(n730), .ZN(G75) );
  NOR2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n738) );
  XNOR2_X1 U788 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n734), .B(KEYINPUT57), .ZN(n735) );
  XNOR2_X1 U790 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U791 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U792 ( .A1(n749), .A2(n739), .ZN(G54) );
  NAND2_X1 U793 ( .A1(n745), .A2(G478), .ZN(n743) );
  XOR2_X1 U794 ( .A(KEYINPUT124), .B(n741), .Z(n742) );
  XNOR2_X1 U795 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n749), .A2(n744), .ZN(G63) );
  NAND2_X1 U797 ( .A1(n745), .A2(G217), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U799 ( .A1(n749), .A2(n748), .ZN(G66) );
  NAND2_X1 U800 ( .A1(n750), .A2(n762), .ZN(n754) );
  NAND2_X1 U801 ( .A1(G953), .A2(G224), .ZN(n751) );
  XNOR2_X1 U802 ( .A(KEYINPUT61), .B(n751), .ZN(n752) );
  NAND2_X1 U803 ( .A1(n752), .A2(G898), .ZN(n753) );
  NAND2_X1 U804 ( .A1(n754), .A2(n753), .ZN(n758) );
  NOR2_X1 U805 ( .A1(n762), .A2(G898), .ZN(n755) );
  NOR2_X1 U806 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U807 ( .A(n758), .B(n757), .ZN(G69) );
  XNOR2_X1 U808 ( .A(n759), .B(KEYINPUT126), .ZN(n761) );
  XNOR2_X1 U809 ( .A(n760), .B(n761), .ZN(n764) );
  XNOR2_X1 U810 ( .A(n683), .B(n764), .ZN(n763) );
  NAND2_X1 U811 ( .A1(n763), .A2(n762), .ZN(n769) );
  XNOR2_X1 U812 ( .A(n764), .B(G227), .ZN(n765) );
  NAND2_X1 U813 ( .A1(n765), .A2(G900), .ZN(n766) );
  NAND2_X1 U814 ( .A1(G953), .A2(n766), .ZN(n767) );
  XOR2_X1 U815 ( .A(KEYINPUT127), .B(n767), .Z(n768) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(G72) );
  XOR2_X1 U817 ( .A(G140), .B(n770), .Z(G42) );
  XOR2_X1 U818 ( .A(G125), .B(KEYINPUT37), .Z(n771) );
  XNOR2_X1 U819 ( .A(n772), .B(n771), .ZN(G27) );
  XNOR2_X1 U820 ( .A(G119), .B(n773), .ZN(G21) );
  XOR2_X1 U821 ( .A(n774), .B(G131), .Z(G33) );
  XOR2_X1 U822 ( .A(n775), .B(G137), .Z(G39) );
endmodule

