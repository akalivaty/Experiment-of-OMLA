//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G13), .ZN(new_n206));
  INV_X1    g0006(.A(KEYINPUT65), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g0008(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G20), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT66), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n202), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT67), .Z(new_n216));
  AND2_X1   g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT0), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT68), .B(G68), .ZN(new_n225));
  INV_X1    g0025(.A(G238), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G58), .A2(G232), .ZN(new_n231));
  NAND4_X1  g0031(.A1(new_n228), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n221), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n224), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n217), .B(new_n234), .C1(KEYINPUT1), .C2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT69), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n240), .B(new_n243), .Z(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XOR2_X1   g0045(.A(G50), .B(G58), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G179), .ZN(new_n252));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT71), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G33), .A3(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n206), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT70), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n218), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n258), .A2(G274), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g0073(.A1(new_n270), .A2(G223), .B1(new_n273), .B2(G77), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1698), .B1(new_n268), .B2(new_n269), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n210), .A2(new_n253), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n264), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n258), .A2(new_n281), .A3(new_n259), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n258), .B2(new_n259), .ZN(new_n283));
  OAI21_X1  g0083(.A(G226), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n279), .A2(new_n280), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n280), .B1(new_n279), .B2(new_n284), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n252), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n287), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n289), .A2(new_n290), .A3(new_n285), .ZN(new_n291));
  INV_X1    g0091(.A(G58), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(KEYINPUT8), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(KEYINPUT8), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(KEYINPUT74), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n294), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n219), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g0103(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n208), .A2(new_n209), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n208), .A2(new_n307), .A3(new_n209), .A4(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n218), .A2(G20), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G50), .ZN(new_n310));
  OAI22_X1  g0110(.A1(new_n308), .A2(new_n310), .B1(G50), .B2(new_n307), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n288), .A2(new_n291), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(G190), .B1(new_n286), .B2(new_n287), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n289), .A2(G200), .A3(new_n285), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n306), .A2(KEYINPUT9), .A3(new_n312), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT9), .ZN(new_n319));
  INV_X1    g0119(.A(new_n305), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n320), .B1(new_n300), .B2(new_n302), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n319), .B1(new_n321), .B2(new_n311), .ZN(new_n322));
  AND2_X1   g0122(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n316), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT10), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT10), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n316), .A2(new_n317), .A3(new_n323), .A4(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n315), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT75), .ZN(new_n329));
  INV_X1    g0129(.A(G244), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n258), .A2(new_n259), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT72), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n258), .A2(new_n281), .A3(new_n259), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n329), .B1(new_n334), .B2(new_n264), .ZN(new_n335));
  OAI21_X1  g0135(.A(G244), .B1(new_n282), .B2(new_n283), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT75), .A3(new_n263), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n275), .A2(G232), .B1(new_n273), .B2(G107), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n270), .A2(G238), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n278), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n335), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(G179), .ZN(new_n343));
  INV_X1    g0143(.A(new_n308), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(G77), .A3(new_n309), .ZN(new_n345));
  NAND2_X1  g0145(.A1(G20), .A2(G77), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  INV_X1    g0147(.A(new_n295), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n293), .ZN(new_n349));
  INV_X1    g0149(.A(new_n301), .ZN(new_n350));
  OAI221_X1 g0150(.A(new_n346), .B1(new_n347), .B2(new_n298), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  INV_X1    g0152(.A(new_n307), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n351), .A2(new_n305), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n342), .A2(new_n290), .B1(new_n345), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n343), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(G200), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n210), .A2(new_n253), .ZN(new_n359));
  INV_X1    g0159(.A(G87), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n267), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n270), .B2(G226), .ZN(new_n362));
  OAI211_X1 g0162(.A(G223), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n258), .A2(G232), .A3(new_n259), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n263), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n358), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(G226), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n363), .B(new_n368), .C1(new_n267), .C2(new_n360), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n278), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n370), .A2(new_n371), .A3(new_n263), .A4(new_n365), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT16), .ZN(new_n374));
  INV_X1    g0174(.A(G159), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n350), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G68), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT68), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT68), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n202), .B1(new_n382), .B2(G58), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n377), .B1(new_n383), .B2(new_n219), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n268), .A2(new_n219), .A3(new_n269), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n269), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n225), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n374), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n273), .B2(new_n219), .ZN(new_n391));
  INV_X1    g0191(.A(new_n388), .ZN(new_n392));
  OAI21_X1  g0192(.A(G68), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n214), .B1(new_n225), .B2(new_n292), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n376), .B1(new_n394), .B2(G20), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n390), .A2(new_n396), .A3(new_n305), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n297), .A2(new_n309), .ZN(new_n398));
  INV_X1    g0198(.A(new_n297), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n398), .A2(new_n344), .B1(new_n353), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n373), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  XOR2_X1   g0201(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT17), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n373), .A2(new_n397), .A3(new_n400), .A4(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n397), .A2(new_n400), .ZN(new_n409));
  OAI21_X1  g0209(.A(G169), .B1(new_n364), .B2(new_n366), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n370), .A2(G179), .A3(new_n263), .A4(new_n365), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT18), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n357), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n299), .A2(G77), .B1(new_n301), .B2(G50), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n225), .A2(G20), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n305), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT11), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n307), .A2(G68), .ZN(new_n425));
  INV_X1    g0225(.A(G13), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n426), .A2(G1), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT12), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n424), .B1(KEYINPUT12), .B2(new_n425), .C1(new_n420), .C2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n344), .A2(G68), .A3(new_n309), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n422), .B2(new_n423), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n226), .B1(new_n332), .B2(new_n333), .ZN(new_n433));
  NOR2_X1   g0233(.A1(G226), .A2(G1698), .ZN(new_n434));
  INV_X1    g0234(.A(G232), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n268), .A2(new_n269), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n436), .A2(new_n437), .B1(G33), .B2(G97), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n263), .B1(new_n438), .B2(new_n359), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT13), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n441));
  INV_X1    g0241(.A(G274), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n261), .A2(new_n262), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G97), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n435), .A2(G1698), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(G226), .B2(G1698), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n447), .B2(new_n273), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n443), .A2(new_n444), .B1(new_n278), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(G238), .B1(new_n282), .B2(new_n283), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT13), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n440), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G200), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n440), .A2(G190), .A3(new_n452), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n432), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n440), .A2(G179), .A3(new_n452), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT78), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT14), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n433), .A2(KEYINPUT13), .A3(new_n439), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n451), .B1(new_n449), .B2(new_n450), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n460), .B(G169), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n290), .B1(new_n440), .B2(new_n452), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(KEYINPUT78), .A3(new_n460), .ZN(new_n466));
  OAI21_X1  g0266(.A(KEYINPUT14), .B1(new_n465), .B2(KEYINPUT77), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n453), .A2(KEYINPUT77), .A3(G169), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n464), .B(new_n466), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n432), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n457), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n342), .A2(new_n371), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n354), .A2(new_n345), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n342), .B2(G200), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n472), .B1(new_n475), .B2(KEYINPUT76), .ZN(new_n476));
  AOI211_X1 g0276(.A(KEYINPUT76), .B(new_n473), .C1(new_n342), .C2(G200), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n328), .A2(new_n418), .A3(new_n471), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n258), .A2(G274), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n482), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n258), .A2(new_n488), .A3(G257), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT81), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n484), .A2(new_n489), .A3(KEYINPUT81), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT4), .A2(G244), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n265), .B(new_n495), .C1(new_n271), .C2(new_n272), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n330), .B1(new_n268), .B2(new_n269), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g0299(.A(G250), .B1(new_n271), .B2(new_n272), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n265), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n278), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT80), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n504), .B(new_n278), .C1(new_n499), .C2(new_n501), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n494), .A2(new_n503), .A3(new_n252), .A4(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n484), .A3(new_n489), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n290), .ZN(new_n508));
  AND2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT6), .ZN(new_n510));
  AND2_X1   g0310(.A1(G97), .A2(G107), .ZN(new_n511));
  NOR2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n514), .A2(KEYINPUT6), .A3(G97), .ZN(new_n515));
  AND2_X1   g0315(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n516), .A2(new_n219), .B1(new_n352), .B2(new_n350), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n387), .B2(new_n388), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n305), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(G97), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n353), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n267), .A2(G1), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n320), .A2(new_n307), .A3(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n520), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n519), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT82), .ZN(new_n528));
  OAI21_X1  g0328(.A(G107), .B1(new_n391), .B2(new_n392), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n513), .A2(new_n515), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n530), .A2(G20), .B1(G77), .B2(new_n301), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n320), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n532), .A2(new_n525), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT82), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n528), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n494), .A2(new_n503), .A3(new_n505), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G200), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G1698), .ZN(new_n540));
  OR2_X1    g0340(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n496), .A2(new_n497), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n490), .B1(new_n543), .B2(new_n278), .ZN(new_n544));
  AOI211_X1 g0344(.A(new_n525), .B(new_n532), .C1(new_n544), .C2(G190), .ZN(new_n545));
  AOI22_X1  g0345(.A1(new_n509), .A2(new_n536), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n320), .A2(G116), .A3(new_n307), .A4(new_n523), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n353), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(G20), .B1(G33), .B2(G283), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n267), .A2(G97), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(G20), .B2(new_n548), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n552), .A2(new_n305), .A3(KEYINPUT20), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT20), .B1(new_n552), .B2(new_n305), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n547), .B(new_n549), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G264), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n556));
  OAI211_X1 g0356(.A(G257), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n268), .A2(G303), .A3(new_n269), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n278), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n258), .A2(new_n488), .A3(G270), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n484), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(G200), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n563), .A2(KEYINPUT85), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n562), .A2(new_n371), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n563), .B2(KEYINPUT85), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G33), .A2(G116), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n567), .A2(G20), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT87), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n219), .B2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT23), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT23), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n569), .B(new_n572), .C1(new_n219), .C2(G107), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n568), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g0374(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n437), .A2(new_n575), .A3(new_n219), .A4(G87), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n219), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n577));
  XOR2_X1   g0377(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT24), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n320), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n574), .A2(new_n576), .A3(new_n579), .A4(KEYINPUT24), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(G257), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n585));
  OAI211_X1 g0385(.A(G250), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n586));
  NAND2_X1  g0386(.A1(G33), .A2(G294), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n278), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n258), .A2(new_n488), .A3(G264), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n484), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT89), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n358), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n218), .A2(new_n514), .A3(G13), .A4(G20), .ZN(new_n594));
  XOR2_X1   g0394(.A(new_n594), .B(KEYINPUT25), .Z(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(KEYINPUT88), .C1(new_n524), .C2(new_n514), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT88), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n308), .A2(new_n514), .A3(new_n522), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n594), .B(KEYINPUT25), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n584), .A2(new_n593), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n592), .B1(new_n591), .B2(new_n358), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(G190), .B2(new_n591), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n564), .A2(new_n566), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT19), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n219), .B1(new_n445), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n512), .A2(new_n360), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n219), .B(G68), .C1(new_n271), .C2(new_n272), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n606), .B1(new_n298), .B2(new_n520), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n305), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n344), .A2(G87), .A3(new_n523), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n347), .A2(new_n353), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(G244), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n617));
  OAI211_X1 g0417(.A(G238), .B(new_n265), .C1(new_n271), .C2(new_n272), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n618), .A3(new_n567), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n278), .ZN(new_n620));
  INV_X1    g0420(.A(G250), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n481), .B2(G1), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n218), .A2(new_n442), .A3(G45), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n441), .A2(KEYINPUT83), .A3(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT83), .ZN(new_n626));
  INV_X1    g0426(.A(new_n624), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n626), .B1(new_n627), .B2(new_n258), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n620), .B(G190), .C1(new_n625), .C2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT83), .B1(new_n441), .B2(new_n624), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n626), .A3(new_n258), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n630), .A2(new_n631), .B1(new_n278), .B2(new_n619), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n616), .B(new_n629), .C1(new_n358), .C2(new_n632), .ZN(new_n633));
  OAI211_X1 g0433(.A(new_n620), .B(new_n252), .C1(new_n625), .C2(new_n628), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT84), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n347), .B(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n613), .B(new_n615), .C1(new_n524), .C2(new_n636), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n634), .B(new_n637), .C1(G169), .C2(new_n632), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n555), .A2(new_n562), .A3(G169), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT21), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n484), .A2(new_n561), .ZN(new_n643));
  NAND4_X1  g0443(.A1(new_n555), .A2(G179), .A3(new_n560), .A4(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n555), .A2(new_n562), .A3(KEYINPUT21), .A4(G169), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n591), .A2(new_n290), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(G179), .B2(new_n591), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n582), .A2(new_n583), .B1(new_n596), .B2(new_n600), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n546), .A2(new_n605), .A3(new_n639), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n480), .A2(new_n652), .ZN(G372));
  NAND2_X1  g0453(.A1(new_n469), .A2(new_n470), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n457), .B2(new_n356), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n417), .B1(new_n655), .B2(new_n407), .ZN(new_n656));
  INV_X1    g0456(.A(new_n325), .ZN(new_n657));
  INV_X1    g0457(.A(new_n327), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n314), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT91), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(KEYINPUT91), .B(new_n314), .C1(new_n656), .C2(new_n659), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n480), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n509), .A2(new_n639), .A3(new_n666), .A4(new_n527), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n638), .B(KEYINPUT90), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n506), .A2(new_n633), .A3(new_n638), .A4(new_n508), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n534), .B1(new_n519), .B2(new_n526), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n532), .A2(KEYINPUT82), .A3(new_n525), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n667), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n648), .A2(new_n649), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n645), .A2(new_n644), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n290), .B1(new_n643), .B2(new_n560), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT21), .B1(new_n678), .B2(new_n555), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n602), .A2(new_n604), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n546), .A2(new_n639), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n665), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n664), .A2(new_n685), .ZN(G369));
  NAND2_X1  g0486(.A1(new_n427), .A2(new_n219), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(KEYINPUT27), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(new_n689), .A3(G213), .ZN(new_n690));
  INV_X1    g0490(.A(G343), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n646), .A2(new_n555), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n564), .A2(new_n566), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n555), .A2(new_n692), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n680), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT92), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n676), .A2(new_n692), .ZN(new_n700));
  INV_X1    g0500(.A(new_n692), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n649), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n702), .B1(new_n604), .B2(new_n602), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n700), .B1(new_n704), .B2(new_n676), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n646), .A2(new_n701), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT93), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n700), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(G399));
  INV_X1    g0510(.A(new_n222), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(G41), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n608), .A2(G116), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(G1), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n215), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT28), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n681), .A2(new_n682), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n545), .A2(new_n538), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n508), .B(new_n506), .C1(new_n671), .C2(new_n672), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(new_n639), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n667), .A2(new_n669), .A3(new_n674), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n701), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n724), .A2(KEYINPUT29), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n509), .A2(new_n639), .A3(new_n536), .A4(new_n666), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT26), .B1(new_n670), .B2(new_n533), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n669), .A3(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n701), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT29), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n643), .A2(G179), .A3(new_n560), .ZN(new_n731));
  AND2_X1   g0531(.A1(new_n589), .A2(new_n590), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n544), .A3(new_n632), .A4(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT30), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n732), .A2(new_n632), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(KEYINPUT30), .A3(new_n544), .A4(new_n731), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n620), .B1(new_n625), .B2(new_n628), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n738), .A2(new_n562), .A3(new_n252), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n537), .A2(new_n739), .A3(new_n591), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n741), .A2(new_n742), .A3(new_n692), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n742), .B1(new_n741), .B2(new_n692), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n652), .A2(new_n692), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G330), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n725), .A2(new_n730), .A3(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n717), .B1(new_n748), .B2(G1), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT94), .ZN(G364));
  XOR2_X1   g0550(.A(new_n698), .B(KEYINPUT92), .Z(new_n751));
  NOR2_X1   g0551(.A1(new_n426), .A2(G20), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n218), .B1(new_n752), .B2(G45), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n712), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n751), .B(new_n756), .C1(G330), .C2(new_n697), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n711), .A2(new_n273), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G355), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G116), .B2(new_n222), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n222), .A2(new_n273), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT95), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n763), .B1(new_n481), .B2(new_n216), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n247), .A2(G45), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n760), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G13), .A2(G33), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(G20), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n210), .B1(new_n219), .B2(G169), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n755), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n219), .A2(new_n252), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT33), .B(G317), .Z(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(G190), .A3(new_n358), .ZN(new_n780));
  INV_X1    g0580(.A(G322), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT100), .Z(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n775), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n219), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G311), .A2(new_n786), .B1(new_n789), .B2(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(new_n371), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(G294), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n371), .A2(G179), .A3(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n219), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n790), .B1(new_n791), .B2(new_n792), .C1(new_n793), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT98), .B(G326), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n796), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n273), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT99), .Z(new_n805));
  NAND3_X1  g0605(.A1(new_n783), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n802), .A2(new_n360), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n789), .A2(G159), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(KEYINPUT32), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n807), .B(new_n809), .C1(G68), .C2(new_n777), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n437), .B1(new_n785), .B2(new_n352), .ZN(new_n811));
  INV_X1    g0611(.A(new_n780), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n811), .B1(G58), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n792), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n808), .A2(KEYINPUT32), .B1(G107), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n795), .ZN(new_n816));
  INV_X1    g0616(.A(new_n797), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G97), .A2(new_n816), .B1(new_n817), .B2(G50), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n810), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n770), .B1(new_n806), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n774), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n769), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n697), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n757), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NAND2_X1  g0625(.A1(new_n473), .A2(new_n692), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT76), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n474), .A2(new_n827), .B1(new_n371), .B2(new_n342), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n826), .B1(new_n828), .B2(new_n477), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n829), .A2(new_n356), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n356), .A2(new_n692), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n724), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n692), .B1(new_n675), .B2(new_n683), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(new_n829), .B2(new_n356), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n755), .B1(new_n836), .B2(new_n746), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n837), .B1(new_n746), .B2(new_n836), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n797), .A2(new_n803), .B1(new_n792), .B2(new_n360), .ZN(new_n839));
  INV_X1    g0639(.A(new_n802), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(G107), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n437), .B1(new_n786), .B2(G116), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n812), .A2(G294), .B1(new_n789), .B2(G311), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G97), .A2(new_n816), .B1(new_n777), .B2(G283), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n792), .A2(new_n378), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n273), .B(new_n846), .C1(G132), .C2(new_n789), .ZN(new_n847));
  INV_X1    g0647(.A(G50), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n848), .B2(new_n802), .C1(new_n292), .C2(new_n795), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT102), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n812), .A2(G143), .B1(new_n786), .B2(G159), .ZN(new_n851));
  INV_X1    g0651(.A(G150), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n852), .B2(new_n778), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G137), .B2(new_n817), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT34), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n845), .B1(new_n850), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n771), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n770), .A2(new_n768), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT101), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n756), .B1(new_n860), .B2(new_n352), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n857), .B(new_n861), .C1(new_n834), .C2(new_n768), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n838), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n530), .B(KEYINPUT103), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n213), .B(G116), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n868), .B(KEYINPUT36), .ZN(new_n869));
  INV_X1    g0669(.A(new_n215), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n870), .B(G77), .C1(new_n292), .C2(new_n225), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n201), .A2(G68), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n218), .B(G13), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g0674(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n875));
  NAND2_X1  g0675(.A1(new_n396), .A2(new_n305), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT16), .B1(new_n393), .B2(new_n395), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n400), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n690), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n408), .B2(new_n417), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n410), .A2(new_n411), .A3(new_n690), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n409), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  AND3_X1   g0685(.A1(new_n884), .A2(new_n885), .A3(new_n401), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n883), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n885), .B1(new_n887), .B2(new_n401), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n882), .A2(new_n889), .A3(KEYINPUT38), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT38), .ZN(new_n891));
  AOI221_X4 g0691(.A(KEYINPUT18), .B1(new_n410), .B2(new_n411), .C1(new_n397), .C2(new_n400), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n415), .B1(new_n409), .B2(new_n412), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n880), .B1(new_n894), .B2(new_n407), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n886), .A2(new_n888), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT105), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(KEYINPUT105), .B(new_n891), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n470), .B(new_n692), .C1(new_n469), .C2(new_n457), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n432), .A2(new_n701), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n457), .B(new_n904), .C1(new_n469), .C2(new_n470), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n745), .A2(new_n834), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n875), .B1(new_n901), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n409), .A2(new_n879), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n894), .B2(new_n407), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n884), .A2(new_n401), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT106), .B1(new_n409), .B2(new_n883), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n885), .B2(new_n914), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n884), .A2(new_n401), .A3(KEYINPUT106), .A4(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n891), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n910), .B1(new_n918), .B2(new_n890), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n909), .B1(new_n908), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n665), .A2(new_n745), .ZN(new_n921));
  OAI21_X1  g0721(.A(G330), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT108), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n920), .A2(new_n921), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT39), .B1(new_n918), .B2(new_n890), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n899), .A2(new_n900), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(KEYINPUT39), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n654), .A2(new_n692), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n933));
  OAI21_X1  g0733(.A(KEYINPUT104), .B1(new_n933), .B2(new_n906), .ZN(new_n934));
  INV_X1    g0734(.A(new_n831), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n724), .B2(new_n830), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  INV_X1    g0737(.A(new_n904), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n471), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n902), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n941), .A3(new_n901), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n417), .A2(new_n690), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n932), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n725), .A2(new_n730), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n662), .A2(new_n663), .B1(new_n665), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n927), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n218), .B2(new_n752), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n927), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n874), .B1(new_n949), .B2(new_n950), .ZN(G367));
  NOR2_X1   g0751(.A1(new_n533), .A2(new_n701), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  MUX2_X1   g0753(.A(new_n509), .B(new_n546), .S(new_n953), .Z(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n705), .A3(new_n708), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT42), .Z(new_n956));
  AND2_X1   g0756(.A1(new_n954), .A2(new_n650), .ZN(new_n957));
  INV_X1    g0757(.A(new_n720), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n701), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n701), .A2(new_n616), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n669), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n963), .B1(new_n639), .B2(new_n962), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n960), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n961), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT109), .Z(new_n967));
  AND2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n967), .ZN(new_n969));
  INV_X1    g0769(.A(new_n706), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n954), .ZN(new_n971));
  OR3_X1    g0771(.A1(new_n968), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n971), .B1(new_n968), .B2(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n709), .A2(new_n954), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT110), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT110), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n709), .A2(new_n977), .A3(new_n954), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n709), .A2(new_n954), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT44), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n976), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n970), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n705), .B(new_n708), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n699), .B(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n981), .A2(new_n983), .A3(new_n706), .A4(new_n984), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n986), .A2(new_n748), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n748), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n712), .B(KEYINPUT41), .Z(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n754), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n964), .A2(new_n769), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n762), .A2(new_n243), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n996), .B(new_n772), .C1(new_n222), .C2(new_n347), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n795), .A2(new_n378), .B1(new_n792), .B2(new_n352), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n437), .B1(new_n201), .B2(new_n785), .C1(new_n852), .C2(new_n780), .ZN(new_n999));
  AOI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(G159), .C2(new_n777), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n840), .A2(G58), .B1(new_n789), .B2(G137), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n799), .A2(G143), .B1(KEYINPUT112), .B2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(KEYINPUT112), .C2(new_n1001), .ZN(new_n1003));
  INV_X1    g0803(.A(G317), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n273), .B1(new_n788), .B2(new_n1004), .C1(new_n791), .C2(new_n785), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n778), .A2(new_n793), .B1(new_n792), .B2(new_n520), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(G107), .C2(new_n816), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n840), .A2(G116), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT111), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n799), .A2(G311), .B1(G303), .B2(new_n812), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1007), .B(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1011), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(KEYINPUT111), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1003), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  OAI211_X1 g0816(.A(new_n755), .B(new_n997), .C1(new_n1016), .C2(new_n770), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n974), .A2(new_n994), .B1(new_n995), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(KEYINPUT113), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1018), .B(new_n1019), .ZN(G387));
  AOI21_X1  g0820(.A(new_n713), .B1(new_n988), .B2(new_n748), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n748), .B2(new_n988), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n988), .A2(new_n754), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n714), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n758), .A2(new_n1024), .B1(new_n514), .B2(new_n711), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n240), .A2(new_n481), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n349), .A2(G50), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT50), .Z(new_n1028));
  OAI211_X1 g0828(.A(new_n714), .B(new_n481), .C1(new_n378), .C2(new_n352), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n762), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1025), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n756), .B1(new_n1031), .B2(new_n772), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n797), .A2(new_n375), .B1(new_n792), .B2(new_n520), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n780), .A2(new_n848), .B1(new_n788), .B2(new_n852), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n273), .B(new_n1034), .C1(G68), .C2(new_n786), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n636), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n816), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n399), .C2(new_n778), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1033), .B(new_n1038), .C1(G77), .C2(new_n840), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n812), .A2(G317), .B1(new_n786), .B2(G303), .ZN(new_n1040));
  INV_X1    g0840(.A(G311), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1040), .B1(new_n1041), .B2(new_n778), .C1(new_n798), .C2(new_n781), .ZN(new_n1042));
  INV_X1    g0842(.A(KEYINPUT48), .ZN(new_n1043));
  OR2_X1    g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n816), .A2(G283), .B1(new_n840), .B2(G294), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n789), .A2(new_n800), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1050), .B(new_n273), .C1(new_n548), .C2(new_n792), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1039), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1032), .B1(new_n705), .B2(new_n822), .C1(new_n1054), .C2(new_n770), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1023), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1022), .A2(new_n1056), .ZN(G393));
  NAND2_X1  g0857(.A1(new_n986), .A2(new_n989), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n988), .A2(new_n748), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n712), .A3(new_n990), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n986), .A2(new_n754), .A3(new_n989), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n772), .B1(new_n520), .B2(new_n222), .C1(new_n763), .C2(new_n250), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n755), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n778), .A2(new_n201), .B1(new_n792), .B2(new_n360), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n273), .B1(new_n789), .B2(G143), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n349), .B2(new_n785), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n795), .A2(new_n352), .B1(new_n802), .B2(new_n225), .ZN(new_n1068));
  OR3_X1    g0868(.A1(new_n1065), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n852), .A2(new_n797), .B1(new_n780), .B2(new_n375), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  OAI22_X1  g0871(.A1(new_n778), .A2(new_n803), .B1(new_n548), .B2(new_n795), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n273), .B1(new_n788), .B2(new_n781), .C1(new_n793), .C2(new_n785), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n514), .A2(new_n792), .B1(new_n802), .B2(new_n791), .ZN(new_n1074));
  OR3_X1    g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n1041), .A2(new_n780), .B1(new_n797), .B2(new_n1004), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1076), .B(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1069), .A2(new_n1071), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1064), .B1(new_n1079), .B2(new_n771), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n954), .B2(new_n822), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1062), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1061), .A2(new_n1082), .ZN(G390));
  NAND4_X1  g0883(.A1(new_n940), .A2(G330), .A3(new_n745), .A4(new_n834), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n931), .B1(new_n918), .B2(new_n890), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n728), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n692), .B1(new_n1086), .B2(new_n683), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n829), .A2(new_n356), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n831), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1089), .B2(new_n906), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n931), .B1(new_n936), .B2(new_n940), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1084), .B(new_n1090), .C1(new_n930), .C2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n933), .A2(new_n906), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT39), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n899), .B2(new_n900), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n1094), .A2(new_n931), .B1(new_n1096), .B2(new_n928), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1084), .B1(new_n1097), .B2(new_n1090), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n754), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n756), .B1(new_n860), .B2(new_n399), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(G159), .A2(new_n816), .B1(new_n777), .B2(G137), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n817), .A2(G128), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n201), .C2(new_n792), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(KEYINPUT54), .B(G143), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n437), .B1(new_n785), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(G132), .ZN(new_n1107));
  INV_X1    g0907(.A(G125), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n780), .A2(new_n1107), .B1(new_n788), .B2(new_n1108), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1104), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n802), .A2(new_n852), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G97), .A2(new_n786), .B1(new_n789), .B2(G294), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1113), .B1(new_n548), .B2(new_n780), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n778), .A2(new_n514), .B1(new_n791), .B2(new_n797), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n795), .A2(new_n352), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1114), .A2(new_n1115), .A3(new_n846), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n807), .A2(new_n437), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT116), .Z(new_n1119));
  AOI22_X1  g0919(.A1(new_n1110), .A2(new_n1112), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1101), .B1(new_n770), .B2(new_n1120), .C1(new_n930), .C2(new_n768), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1100), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1090), .B1(new_n930), .B2(new_n1091), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1084), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1092), .ZN(new_n1127));
  INV_X1    g0927(.A(G330), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n906), .B1(new_n907), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1084), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n936), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1129), .A2(new_n1084), .A3(new_n1089), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n746), .A2(new_n480), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n946), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n713), .B1(new_n1127), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g0937(.A1(new_n946), .A2(new_n1135), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1138), .A2(new_n1126), .A3(new_n1092), .A4(new_n1133), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1137), .A2(new_n1139), .A3(KEYINPUT115), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT115), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1123), .B1(new_n1140), .B2(new_n1141), .ZN(G378));
  AOI211_X1 g0942(.A(G41), .B(new_n437), .C1(new_n789), .C2(G283), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n292), .B2(new_n792), .C1(new_n352), .C2(new_n802), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT117), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n795), .A2(new_n378), .B1(new_n780), .B2(new_n514), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n778), .A2(new_n520), .B1(new_n548), .B2(new_n797), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n1036), .C2(new_n786), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT58), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(G33), .A2(G41), .ZN(new_n1151));
  INV_X1    g0951(.A(G41), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1151), .C1(new_n273), .C2(new_n1152), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n778), .A2(new_n1107), .B1(new_n1108), .B2(new_n797), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G150), .B2(new_n816), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n812), .A2(G128), .B1(new_n786), .B2(G137), .ZN(new_n1156));
  OAI211_X1 g0956(.A(new_n1155), .B(new_n1156), .C1(new_n802), .C2(new_n1105), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  INV_X1    g0958(.A(G124), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1151), .B1(new_n788), .B2(new_n1159), .C1(new_n375), .C2(new_n792), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1157), .B2(KEYINPUT59), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n770), .B1(new_n1150), .B2(new_n1162), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n756), .B(new_n1163), .C1(new_n201), .C2(new_n860), .ZN(new_n1164));
  XOR2_X1   g0964(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n328), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n313), .A2(new_n879), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT118), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n328), .A2(new_n1166), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1169), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n328), .A2(new_n1166), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1165), .B(new_n315), .C1(new_n325), .C2(new_n327), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1164), .B1(new_n1176), .B2(new_n768), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT119), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n919), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n745), .B(new_n834), .C1(new_n903), .C2(new_n905), .ZN(new_n1181));
  OAI21_X1  g0981(.A(G330), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1179), .B1(new_n909), .B2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1128), .B1(new_n908), .B2(new_n919), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n875), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1185), .B1(new_n929), .B2(new_n1181), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1186), .A3(new_n1176), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n930), .A2(new_n931), .B1(new_n417), .B2(new_n690), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1183), .A2(new_n1187), .A3(new_n942), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT121), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n944), .A2(KEYINPUT121), .A3(new_n1187), .A4(new_n1183), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT120), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1183), .A2(new_n1187), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n932), .A2(new_n942), .A3(new_n943), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n909), .A2(new_n1182), .A3(new_n1179), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1176), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1194), .B(new_n1196), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1178), .B1(new_n1202), .B2(new_n754), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n946), .A2(new_n1135), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n1099), .B2(new_n1133), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1189), .ZN(new_n1210));
  OAI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n712), .B1(new_n1211), .B2(new_n1205), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1203), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(KEYINPUT122), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT122), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1215), .B(new_n1203), .C1(new_n1207), .C2(new_n1212), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1214), .A2(new_n1216), .ZN(G375));
  OR2_X1    g1017(.A1(new_n940), .A2(new_n768), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1218), .A2(KEYINPUT123), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n792), .A2(new_n352), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n797), .A2(new_n793), .B1(new_n802), .B2(new_n520), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(G116), .C2(new_n777), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n780), .A2(new_n791), .B1(new_n785), .B2(new_n514), .ZN(new_n1224));
  AOI211_X1 g1024(.A(new_n437), .B(new_n1224), .C1(G303), .C2(new_n789), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1223), .A2(new_n1225), .A3(new_n1037), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n795), .A2(new_n848), .B1(new_n797), .B2(new_n1107), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(G159), .B2(new_n840), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n273), .B1(new_n812), .B2(G137), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G150), .A2(new_n786), .B1(new_n789), .B2(G128), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1105), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n777), .A2(new_n1231), .B1(new_n814), .B2(G58), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n770), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n756), .B(new_n1234), .C1(new_n378), .C2(new_n860), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n1235), .B(KEYINPUT124), .Z(new_n1236));
  NOR3_X1   g1036(.A1(new_n1219), .A2(new_n1220), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n754), .B2(new_n1133), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1136), .A2(new_n993), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1133), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1204), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1239), .B1(new_n1240), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G381));
  NOR4_X1   g1044(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1122), .B1(new_n1139), .B2(new_n1137), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(G375), .A2(G387), .A3(new_n1247), .ZN(G407));
  NAND2_X1  g1048(.A1(new_n691), .A2(G213), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT125), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1246), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(G407), .B(G213), .C1(G375), .C2(new_n1251), .ZN(G409));
  NAND2_X1  g1052(.A1(new_n1136), .A2(KEYINPUT60), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(new_n1242), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1204), .A2(new_n1241), .A3(KEYINPUT60), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1254), .A2(new_n712), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(G384), .A3(new_n1238), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(G384), .B1(new_n1256), .B2(new_n1238), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1249), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(G2897), .A3(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1250), .A2(G2897), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1260), .B2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G378), .B(new_n1203), .C1(new_n1207), .C2(new_n1212), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1201), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(new_n1197), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n992), .B(new_n1205), .C1(new_n1267), .C2(new_n1193), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n754), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1177), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1246), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1265), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT126), .B1(new_n1272), .B2(new_n1249), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT126), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n1274), .B(new_n1261), .C1(new_n1265), .C2(new_n1271), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1264), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(KEYINPUT127), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1278), .B(new_n1264), .C1(new_n1273), .C2(new_n1275), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1250), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1280), .A4(new_n1260), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G393), .A2(G396), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n824), .B1(new_n1022), .B2(new_n1056), .ZN(new_n1283));
  OAI21_X1  g1083(.A(G390), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1019), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1285), .A2(new_n1061), .A3(new_n1082), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1284), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1018), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT61), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1018), .A2(new_n1286), .A3(new_n1284), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1289), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1281), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1261), .B1(new_n1265), .B2(new_n1271), .ZN(new_n1294));
  AOI21_X1  g1094(.A(KEYINPUT63), .B1(new_n1294), .B2(new_n1260), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1277), .A2(new_n1279), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1272), .A2(new_n1280), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1260), .ZN(new_n1300));
  OAI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1298), .B2(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT62), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1294), .A2(new_n1302), .A3(new_n1260), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1299), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1297), .A2(new_n1306), .ZN(G405));
  NAND3_X1  g1107(.A1(new_n1214), .A2(new_n1216), .A3(new_n1246), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(new_n1265), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1309), .A2(new_n1260), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1308), .A2(new_n1300), .A3(new_n1265), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1312), .A2(new_n1305), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1310), .A2(new_n1289), .A3(new_n1291), .A4(new_n1311), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(G402));
endmodule


