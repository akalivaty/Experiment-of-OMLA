//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:45 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n240,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1277, new_n1278, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n206), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n209), .B1(new_n213), .B2(new_n214), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XOR2_X1   g0023(.A(G250), .B(G257), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT65), .ZN(new_n225));
  XNOR2_X1  g0025(.A(G264), .B(G270), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n227), .B(new_n231), .ZN(G358));
  XOR2_X1   g0032(.A(G87), .B(G97), .Z(new_n233));
  XNOR2_X1  g0033(.A(G107), .B(G116), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G68), .B(G77), .Z(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G351));
  INV_X1    g0039(.A(G1), .ZN(new_n240));
  NAND3_X1  g0040(.A1(new_n240), .A2(G13), .A3(G20), .ZN(new_n241));
  INV_X1    g0041(.A(KEYINPUT68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g0043(.A1(new_n240), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n210), .B1(new_n206), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n245), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n251), .B1(new_n240), .B2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(new_n245), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n250), .A2(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT8), .B(G58), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n211), .A2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G20), .A2(G33), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n256), .A2(new_n258), .B1(G150), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n203), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT67), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT67), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n203), .A2(new_n264), .A3(G20), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g0066(.A(KEYINPUT9), .B(new_n254), .C1(new_n266), .C2(new_n248), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G223), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n270), .B1(new_n271), .B2(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n240), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(new_n276), .A3(G274), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n279), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n276), .A2(KEYINPUT66), .A3(new_n279), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(G226), .ZN(new_n287));
  NAND4_X1  g0087(.A1(new_n278), .A2(G190), .A3(new_n281), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n267), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n265), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n264), .B1(new_n203), .B2(G20), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n260), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n247), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT9), .B1(new_n293), .B2(new_n254), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n278), .A2(new_n281), .A3(new_n287), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT70), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n295), .B(new_n297), .C1(new_n298), .C2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(G238), .ZN(new_n300));
  INV_X1    g0100(.A(G107), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n272), .A2(new_n300), .B1(new_n301), .B2(new_n268), .ZN(new_n302));
  AND3_X1   g0102(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n277), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n281), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n305), .B1(new_n286), .B2(G244), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT69), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n245), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n243), .A2(KEYINPUT69), .A3(new_n244), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n240), .A2(G20), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(G77), .A3(new_n248), .A4(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n259), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n255), .A2(new_n316), .B1(new_n211), .B2(new_n271), .ZN(new_n317));
  XNOR2_X1  g0117(.A(KEYINPUT15), .B(G87), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n318), .A2(new_n257), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n247), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n315), .B(new_n320), .C1(G77), .C2(new_n313), .ZN(new_n321));
  INV_X1    g0121(.A(G200), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n304), .B2(new_n306), .ZN(new_n323));
  OR3_X1    g0123(.A1(new_n309), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n307), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n321), .B(new_n326), .C1(G179), .C2(new_n307), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n254), .B1(new_n266), .B2(new_n248), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT9), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n331), .A2(new_n297), .A3(new_n288), .A4(new_n267), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n331), .A2(new_n298), .A3(new_n288), .A4(new_n267), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT10), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  OR2_X1    g0135(.A1(new_n296), .A2(G179), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n296), .A2(new_n325), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n329), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n299), .A2(new_n328), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT71), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT79), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n255), .B1(new_n240), .B2(G20), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n250), .A2(new_n343), .B1(new_n255), .B2(new_n253), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n268), .A2(new_n346), .A3(G20), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(G33), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(KEYINPUT7), .B1(new_n351), .B2(new_n211), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT74), .ZN(new_n354));
  AND2_X1   g0154(.A1(G58), .A2(G68), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT73), .B(G20), .C1(new_n355), .C2(new_n202), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n259), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(G58), .B(G68), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT73), .B1(new_n359), .B2(G20), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n354), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(G20), .B1(new_n355), .B2(new_n202), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT74), .A3(new_n357), .A4(new_n356), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n353), .A2(new_n361), .A3(KEYINPUT16), .A4(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT75), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G68), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n346), .B1(new_n268), .B2(G20), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n351), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(KEYINPUT75), .A3(new_n361), .A4(new_n365), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n357), .A3(new_n356), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n373), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n247), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n345), .B1(new_n376), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n276), .A2(G232), .A3(new_n279), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n281), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n348), .A2(new_n350), .A3(G226), .A4(G1698), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n348), .A2(new_n350), .A3(G223), .A4(new_n269), .ZN(new_n385));
  NAND2_X1  g0185(.A1(G33), .A2(G87), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n383), .B1(new_n277), .B2(new_n387), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n388), .A2(new_n308), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(G200), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n342), .B1(new_n381), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n379), .B1(new_n368), .B2(new_n375), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n396));
  NOR4_X1   g0196(.A1(new_n394), .A2(new_n391), .A3(new_n345), .A4(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  INV_X1    g0199(.A(new_n383), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n387), .A2(new_n277), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n400), .A2(new_n401), .A3(G179), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n325), .B1(new_n400), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n399), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n401), .A3(G179), .ZN(new_n405));
  OAI211_X1 g0205(.A(new_n405), .B(KEYINPUT76), .C1(new_n388), .C2(new_n325), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT18), .B1(new_n381), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n404), .A2(new_n406), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n409), .B(new_n410), .C1(new_n394), .C2(new_n345), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(KEYINPUT78), .B1(new_n398), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n316), .A2(new_n251), .ZN(new_n414));
  OAI22_X1  g0214(.A1(new_n257), .A2(new_n271), .B1(new_n211), .B2(G68), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n247), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT11), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n313), .A2(G68), .A3(new_n248), .A4(new_n314), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n311), .A2(KEYINPUT12), .A3(new_n369), .A4(new_n312), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT12), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n245), .B2(G68), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n417), .A2(new_n418), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT13), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n305), .B1(new_n286), .B2(G238), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n348), .A2(new_n350), .A3(G232), .A4(G1698), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n348), .A2(new_n350), .A3(G226), .A4(new_n269), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G97), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n277), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n425), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n276), .A2(KEYINPUT66), .A3(new_n279), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT66), .B1(new_n276), .B2(new_n279), .ZN(new_n434));
  OAI21_X1  g0234(.A(G238), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AND4_X1   g0235(.A1(new_n425), .A2(new_n431), .A3(new_n435), .A4(new_n281), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n424), .B(G169), .C1(new_n432), .C2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n426), .A2(new_n425), .A3(new_n431), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n431), .A2(new_n435), .A3(new_n281), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT13), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n440), .A3(G179), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n437), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n440), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n424), .B1(new_n443), .B2(G169), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT72), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n432), .B2(new_n436), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT14), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT72), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n441), .A4(new_n437), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n423), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n423), .B1(new_n308), .B2(new_n443), .ZN(new_n451));
  INV_X1    g0251(.A(new_n443), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n452), .A2(new_n322), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n396), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n381), .A2(new_n392), .A3(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n394), .A2(new_n345), .A3(new_n391), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n457), .B1(new_n458), .B2(new_n342), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT78), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n408), .A4(new_n411), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n413), .A2(new_n455), .A3(new_n461), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n340), .A2(new_n341), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n341), .B1(new_n340), .B2(new_n462), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT87), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n348), .A2(new_n350), .A3(G264), .A4(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n348), .A2(new_n350), .A3(G257), .A4(new_n269), .ZN(new_n468));
  INV_X1    g0268(.A(G303), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(new_n268), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n277), .ZN(new_n471));
  INV_X1    g0271(.A(G41), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n240), .B(G45), .C1(new_n472), .C2(KEYINPUT5), .ZN(new_n475));
  OAI211_X1 g0275(.A(G270), .B(new_n276), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n276), .A2(G274), .A3(new_n473), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OR2_X1    g0278(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(KEYINPUT80), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n471), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT84), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT84), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n471), .A2(new_n484), .A3(new_n476), .A4(new_n481), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(G169), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(G33), .A2(G283), .ZN(new_n487));
  INV_X1    g0287(.A(G97), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n211), .C1(G33), .C2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  INV_X1    g0291(.A(G116), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(G20), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n493), .A3(new_n247), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT86), .A2(KEYINPUT20), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n311), .A2(new_n492), .A3(new_n312), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n246), .A2(G1), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n499), .A2(new_n492), .ZN(new_n500));
  INV_X1    g0300(.A(new_n312), .ZN(new_n501));
  AOI21_X1  g0301(.A(KEYINPUT69), .B1(new_n243), .B2(new_n244), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n248), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT85), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT85), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n313), .A2(new_n505), .A3(new_n248), .A4(new_n500), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n498), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n466), .B1(new_n486), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT21), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n466), .B(new_n510), .C1(new_n486), .C2(new_n507), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n471), .A2(G179), .A3(new_n476), .A4(new_n481), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n483), .A2(G200), .A3(new_n485), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n483), .A2(new_n485), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n507), .B(new_n514), .C1(new_n515), .C2(new_n308), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n509), .A2(new_n511), .A3(new_n513), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT24), .ZN(new_n519));
  OAI22_X1  g0319(.A1(new_n518), .A2(G20), .B1(new_n519), .B2(KEYINPUT89), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n211), .B2(G107), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n301), .A2(KEYINPUT23), .A3(G20), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g0324(.A1(KEYINPUT88), .A2(G87), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n348), .A2(new_n350), .A3(new_n525), .A4(new_n211), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n268), .A2(KEYINPUT22), .A3(new_n211), .A4(new_n525), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT89), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n530), .B1(new_n531), .B2(KEYINPUT24), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n531), .A2(KEYINPUT24), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n524), .A2(new_n528), .A3(new_n529), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n248), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n249), .A2(new_n499), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n253), .A2(KEYINPUT25), .A3(new_n301), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT25), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n245), .B2(G107), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n537), .A2(G107), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n348), .A2(new_n350), .A3(G250), .A4(new_n269), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT80), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n475), .B(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n277), .A2(new_n545), .B1(new_n547), .B2(new_n478), .ZN(new_n548));
  OAI211_X1 g0348(.A(G264), .B(new_n276), .C1(new_n474), .C2(new_n475), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n548), .A2(new_n308), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT90), .ZN(new_n551));
  XNOR2_X1  g0351(.A(new_n549), .B(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(G200), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n536), .B(new_n541), .C1(new_n550), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n548), .A2(new_n552), .ZN(new_n555));
  INV_X1    g0355(.A(G179), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n325), .B1(new_n548), .B2(new_n549), .ZN(new_n558));
  INV_X1    g0358(.A(new_n541), .ZN(new_n559));
  OAI22_X1  g0359(.A1(new_n557), .A2(new_n558), .B1(new_n535), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n211), .B1(new_n429), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G87), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n488), .A3(new_n301), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n348), .A2(new_n350), .A3(new_n211), .A4(G68), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n563), .B1(new_n257), .B2(new_n488), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n247), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT83), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT83), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n562), .A2(new_n574), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n348), .A2(new_n350), .A3(G244), .A4(G1698), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT81), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n268), .A2(new_n579), .A3(G244), .A4(G1698), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n348), .A2(new_n350), .A3(G238), .A4(new_n269), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(new_n518), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(G45), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(G1), .ZN(new_n587));
  INV_X1    g0387(.A(G274), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n587), .A2(G250), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n590), .A2(new_n277), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n585), .A2(new_n277), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n537), .A2(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n589), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n583), .B1(new_n580), .B2(new_n578), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n595), .B1(new_n596), .B2(new_n276), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n576), .A2(new_n593), .A3(new_n594), .A4(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n245), .A2(G97), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n537), .B2(G97), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT6), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n602), .A2(new_n488), .A3(G107), .ZN(new_n603));
  XNOR2_X1  g0403(.A(G97), .B(G107), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  OAI22_X1  g0405(.A1(new_n605), .A2(new_n211), .B1(new_n271), .B2(new_n316), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n301), .B1(new_n370), .B2(new_n371), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n247), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n601), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n348), .A2(new_n350), .A3(G250), .A4(G1698), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n348), .A2(new_n350), .A3(G244), .A4(new_n269), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT4), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n487), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n277), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G257), .B(new_n276), .C1(new_n474), .C2(new_n475), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n481), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n609), .B1(G200), .B2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n617), .A2(new_n308), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n615), .A2(new_n556), .A3(new_n481), .A4(new_n616), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n325), .A2(new_n617), .B1(new_n601), .B2(new_n608), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(G179), .B(new_n595), .C1(new_n596), .C2(new_n276), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n592), .B2(new_n325), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT82), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n623), .B(KEYINPUT82), .C1(new_n592), .C2(new_n325), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n562), .A2(new_n574), .A3(new_n571), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n574), .B1(new_n562), .B2(new_n571), .ZN(new_n629));
  INV_X1    g0429(.A(new_n537), .ZN(new_n630));
  OAI22_X1  g0430(.A1(new_n628), .A2(new_n629), .B1(new_n318), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n561), .A2(new_n599), .A3(new_n622), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n465), .A2(new_n517), .A3(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n617), .A2(new_n325), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n635), .A2(new_n620), .A3(new_n609), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n631), .A2(new_n624), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(new_n599), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n632), .A2(KEYINPUT26), .A3(new_n599), .A4(new_n636), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n638), .A2(KEYINPUT91), .A3(new_n639), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n637), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n509), .A2(new_n511), .A3(new_n513), .A4(new_n560), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n554), .A2(new_n599), .A3(new_n637), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n617), .A2(G200), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n619), .A2(new_n608), .A3(new_n601), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n621), .A2(new_n620), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n646), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n655), .B1(new_n463), .B2(new_n464), .ZN(new_n656));
  INV_X1    g0456(.A(new_n338), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n454), .A2(new_n327), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n459), .B1(new_n450), .B2(new_n658), .ZN(new_n659));
  OAI22_X1  g0459(.A1(new_n394), .A2(new_n345), .B1(new_n403), .B2(new_n402), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(new_n410), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n299), .A2(new_n335), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n657), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(G369));
  NAND3_X1  g0465(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n240), .A2(new_n211), .A3(G13), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(KEYINPUT27), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(G213), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(G343), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n507), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(KEYINPUT92), .ZN(new_n676));
  AND2_X1   g0476(.A1(new_n675), .A2(KEYINPUT92), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n517), .A2(new_n674), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n676), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(G330), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n672), .B1(new_n559), .B2(new_n535), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n561), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT93), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n561), .A2(KEYINPUT93), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n560), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n672), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n680), .A2(new_n690), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n666), .A2(KEYINPUT94), .A3(new_n673), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT94), .B1(new_n666), .B2(new_n673), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n689), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  XNOR2_X1  g0494(.A(new_n672), .B(KEYINPUT95), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n687), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n691), .A2(new_n698), .ZN(G399));
  INV_X1    g0499(.A(new_n207), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G41), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n566), .A2(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(new_n214), .B2(new_n702), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT28), .ZN(new_n706));
  INV_X1    g0506(.A(new_n653), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n647), .A2(KEYINPUT96), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n647), .A2(KEYINPUT96), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n646), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n632), .A2(new_n599), .A3(new_n636), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(KEYINPUT26), .B2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n673), .C1(new_n710), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n655), .A2(new_n696), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  AND3_X1   g0518(.A1(new_n483), .A2(new_n485), .A3(new_n617), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n555), .A2(new_n597), .A3(new_n556), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n548), .A2(new_n552), .A3(new_n616), .A4(new_n615), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n597), .A2(new_n512), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR4_X1   g0526(.A1(new_n723), .A2(new_n597), .A3(KEYINPUT30), .A4(new_n512), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT31), .B1(new_n728), .B2(new_n672), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n696), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n517), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n650), .A2(new_n554), .A3(new_n560), .A4(new_n651), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n632), .A2(new_n599), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n733), .A2(new_n736), .A3(new_n696), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n732), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G330), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n718), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n706), .B1(new_n741), .B2(G1), .ZN(G364));
  AND2_X1   g0542(.A1(new_n211), .A2(G13), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n240), .B1(new_n743), .B2(G45), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n701), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n746), .B1(new_n679), .B2(G330), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n679), .A2(G330), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  XOR2_X1   g0552(.A(new_n752), .B(KEYINPUT99), .Z(new_n753));
  NOR2_X1   g0553(.A1(new_n679), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n746), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n700), .A2(new_n268), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n214), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(new_n586), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n760), .B1(new_n238), .B2(new_n586), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G355), .A2(KEYINPUT97), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n700), .A2(new_n351), .ZN(new_n763));
  NAND2_X1  g0563(.A1(G355), .A2(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n761), .B1(G116), .B2(new_n207), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n210), .B1(G20), .B2(new_n325), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n752), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n756), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n211), .A2(new_n556), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G200), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n308), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n211), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n308), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n772), .A2(G50), .B1(new_n775), .B2(G107), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n771), .A2(G190), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n211), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n776), .B1(new_n369), .B2(new_n778), .C1(new_n488), .C2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G190), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n773), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n783), .A2(KEYINPUT32), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G87), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT32), .B1(new_n783), .B2(new_n784), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n770), .A2(new_n782), .ZN(new_n791));
  INV_X1    g0591(.A(G58), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n770), .A2(G190), .A3(new_n322), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n268), .B1(new_n791), .B2(new_n271), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n781), .A2(new_n785), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n793), .ZN(new_n796));
  INV_X1    g0596(.A(new_n783), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n796), .A2(G322), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G311), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n351), .C1(new_n799), .C2(new_n791), .ZN(new_n800));
  INV_X1    g0600(.A(G317), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n777), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n772), .A2(G326), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n804), .B(new_n805), .C1(new_n469), .C2(new_n786), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n780), .A2(new_n807), .B1(new_n774), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n800), .A2(new_n806), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n767), .B1(new_n795), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n769), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT98), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n747), .A2(new_n749), .B1(new_n755), .B2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n321), .A2(new_n672), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n324), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n327), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n327), .A2(new_n672), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n715), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n820), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n655), .A2(new_n696), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n746), .B1(new_n824), .B2(new_n739), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n825), .B1(new_n739), .B2(new_n824), .ZN(new_n826));
  INV_X1    g0626(.A(new_n791), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n796), .A2(G143), .B1(new_n827), .B2(G159), .ZN(new_n828));
  INV_X1    g0628(.A(new_n772), .ZN(new_n829));
  INV_X1    g0629(.A(G137), .ZN(new_n830));
  INV_X1    g0630(.A(G150), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n828), .B1(new_n829), .B2(new_n830), .C1(new_n831), .C2(new_n778), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(new_n833), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n775), .A2(G68), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n268), .C1(new_n837), .C2(new_n783), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n780), .A2(new_n792), .B1(new_n786), .B2(new_n251), .ZN(new_n839));
  NOR4_X1   g0639(.A1(new_n834), .A2(new_n835), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n772), .A2(G303), .B1(new_n827), .B2(G116), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n808), .B2(new_n778), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT100), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n780), .A2(new_n488), .B1(new_n793), .B2(new_n807), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT101), .Z(new_n845));
  OAI221_X1 g0645(.A(new_n351), .B1(new_n783), .B2(new_n799), .C1(new_n301), .C2(new_n786), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G87), .B2(new_n775), .ZN(new_n847));
  AND3_X1   g0647(.A1(new_n843), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n767), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n767), .A2(new_n750), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n756), .B1(new_n271), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n849), .B(new_n851), .C1(new_n822), .C2(new_n751), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n826), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  INV_X1    g0654(.A(KEYINPUT35), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n605), .A2(new_n855), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n492), .B(new_n213), .C1(new_n605), .C2(new_n855), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n856), .B1(new_n858), .B2(KEYINPUT102), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(KEYINPUT102), .B2(new_n858), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT36), .Z(new_n861));
  NAND2_X1  g0661(.A1(new_n201), .A2(G68), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n759), .B(G77), .C1(new_n792), .C2(new_n369), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n240), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g0665(.A1(new_n633), .A2(new_n517), .A3(new_n695), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n597), .A2(new_n512), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT30), .B1(new_n867), .B2(new_n723), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n724), .A2(new_n725), .A3(new_n722), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n868), .A2(new_n869), .B1(new_n720), .B2(new_n719), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n730), .B1(new_n870), .B2(new_n673), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n672), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(KEYINPUT107), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n870), .A2(new_n730), .A3(new_n673), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n875), .A2(new_n729), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT107), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n737), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n874), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g0679(.A(G330), .B(new_n879), .C1(new_n463), .C2(new_n464), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n409), .B1(new_n394), .B2(new_n345), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n376), .A2(new_n380), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n344), .A3(new_n392), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  INV_X1    g0684(.A(new_n670), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n394), .B2(new_n345), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n881), .A2(new_n883), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n353), .A2(new_n361), .A3(new_n365), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n248), .B1(new_n888), .B2(new_n373), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n361), .A2(new_n365), .ZN(new_n890));
  AOI21_X1  g0690(.A(KEYINPUT75), .B1(new_n890), .B2(new_n374), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n366), .A2(new_n367), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n670), .B1(new_n893), .B2(new_n344), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n402), .A2(new_n403), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n893), .B2(new_n344), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n894), .A2(new_n896), .A3(new_n458), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n887), .B1(new_n897), .B2(new_n884), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n894), .B1(new_n398), .B2(new_n412), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT104), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT104), .A4(KEYINPUT38), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n423), .A2(new_n673), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n445), .A2(new_n449), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n422), .ZN(new_n909));
  INV_X1    g0709(.A(new_n454), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n450), .A2(new_n454), .A3(new_n906), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n822), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n878), .B2(new_n874), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n909), .A2(new_n910), .A3(new_n907), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n906), .B1(new_n450), .B2(new_n454), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n820), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT106), .B1(new_n393), .B2(new_n397), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT106), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n457), .B(new_n919), .C1(new_n458), .C2(new_n342), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n661), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n886), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n883), .A2(new_n660), .A3(new_n886), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT37), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(KEYINPUT105), .A3(KEYINPUT37), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(new_n887), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n923), .B2(new_n929), .ZN(new_n930));
  AND3_X1   g0730(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n879), .B(new_n917), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  AOI22_X1  g0732(.A1(new_n905), .A2(new_n914), .B1(new_n932), .B2(KEYINPUT40), .ZN(new_n933));
  INV_X1    g0733(.A(G330), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n880), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR2_X1    g0735(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n923), .A2(new_n929), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR3_X1   g0739(.A1(new_n866), .A2(KEYINPUT107), .A3(new_n873), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n877), .B1(new_n737), .B2(new_n876), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n917), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(KEYINPUT40), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n902), .A2(new_n901), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n898), .A2(new_n899), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n938), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n904), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT40), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n914), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n879), .C1(new_n463), .C2(new_n464), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n935), .A2(KEYINPUT108), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n936), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n915), .A2(new_n916), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n823), .A2(KEYINPUT103), .A3(new_n819), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT103), .B1(new_n823), .B2(new_n819), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n947), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n661), .A2(new_n885), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n947), .A2(KEYINPUT39), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n937), .A2(new_n938), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT39), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n962), .A2(new_n963), .A3(new_n902), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n909), .A2(new_n672), .ZN(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  OAI211_X1 g0767(.A(new_n958), .B(new_n960), .C1(new_n965), .C2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n717), .B(new_n714), .C1(new_n463), .C2(new_n464), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n664), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n968), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n953), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n240), .B2(new_n743), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n953), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n865), .B1(new_n973), .B2(new_n974), .ZN(G367));
  NOR2_X1   g0775(.A1(new_n227), .A2(new_n758), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n768), .B1(new_n207), .B2(new_n318), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n746), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G283), .A2(new_n827), .B1(new_n797), .B2(G317), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n979), .B(new_n351), .C1(new_n469), .C2(new_n793), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n777), .A2(G294), .B1(new_n775), .B2(G97), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n981), .B1(new_n301), .B2(new_n780), .C1(new_n799), .C2(new_n829), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT46), .B1(new_n786), .B2(new_n492), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n786), .A2(KEYINPUT46), .A3(new_n492), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n980), .B(new_n982), .C1(new_n983), .C2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n777), .A2(G159), .B1(new_n787), .B2(G58), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n369), .B2(new_n780), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n772), .A2(G143), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n271), .B2(new_n774), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n268), .B1(new_n201), .B2(new_n791), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n793), .A2(new_n831), .B1(new_n783), .B2(new_n830), .ZN(new_n991));
  NOR4_X1   g0791(.A1(new_n987), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n985), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  AOI21_X1  g0794(.A(new_n978), .B1(new_n994), .B2(new_n767), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n576), .A2(new_n594), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n672), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n997), .A2(new_n599), .A3(new_n637), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n637), .B2(new_n997), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n999), .A2(new_n753), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT111), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n695), .A2(new_n609), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n622), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n636), .A2(new_n695), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(KEYINPUT44), .B1(new_n698), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT44), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1009), .B(new_n1006), .C1(new_n694), .C2(new_n697), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n691), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n694), .A2(new_n697), .A3(new_n1006), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1017), .A2(new_n1018), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n691), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n692), .A2(new_n693), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n689), .B1(new_n679), .B2(G330), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n691), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1022), .B1(new_n691), .B2(new_n1023), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n740), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1016), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1027), .A2(new_n741), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n701), .B(KEYINPUT41), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n744), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n622), .A2(new_n687), .A3(new_n1003), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n695), .B1(new_n1031), .B2(new_n651), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n689), .B(new_n1006), .C1(new_n692), .C2(new_n693), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1032), .B1(new_n1033), .B2(KEYINPUT42), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT110), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1033), .A2(KEYINPUT42), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1034), .B2(KEYINPUT110), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1035), .A2(new_n1037), .B1(KEYINPUT43), .B2(new_n999), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT109), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1040), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1042), .B(new_n1043), .C1(new_n1035), .C2(new_n1037), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1012), .A2(new_n1007), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1041), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1048), .A2(new_n1044), .B1(new_n1012), .B2(new_n1007), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1002), .B1(new_n1030), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1027), .A2(new_n741), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1029), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n745), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1055), .A2(new_n1050), .A3(KEYINPUT111), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1001), .B1(new_n1052), .B2(new_n1056), .ZN(G387));
  NOR2_X1   g0857(.A1(new_n1026), .A2(new_n702), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n741), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1059), .A2(new_n745), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n268), .B1(new_n797), .B2(G326), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n780), .A2(new_n808), .B1(new_n786), .B2(new_n807), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n796), .A2(G317), .B1(new_n827), .B2(G303), .ZN(new_n1064));
  INV_X1    g0864(.A(G322), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1064), .B1(new_n829), .B2(new_n1065), .C1(new_n799), .C2(new_n778), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT48), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1063), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1068), .B1(new_n1067), .B2(new_n1066), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT49), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1062), .B1(new_n492), .B2(new_n774), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n772), .A2(G159), .ZN(new_n1073));
  XOR2_X1   g0873(.A(new_n1073), .B(KEYINPUT114), .Z(new_n1074));
  XNOR2_X1  g0874(.A(KEYINPUT112), .B(G150), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n786), .A2(new_n271), .B1(new_n783), .B2(new_n1075), .ZN(new_n1076));
  XOR2_X1   g0876(.A(new_n1076), .B(KEYINPUT113), .Z(new_n1077));
  NOR2_X1   g0877(.A1(new_n780), .A2(new_n318), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G97), .B2(new_n775), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n255), .B2(new_n778), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n268), .B1(new_n791), .B2(new_n369), .C1(new_n251), .C2(new_n793), .ZN(new_n1081));
  NOR4_X1   g0881(.A1(new_n1074), .A2(new_n1077), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n767), .B1(new_n1072), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n703), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n763), .A2(new_n1084), .B1(new_n301), .B2(new_n700), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n231), .A2(new_n586), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n256), .A2(new_n251), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(new_n1087), .B(KEYINPUT50), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n703), .B(new_n586), .C1(new_n369), .C2(new_n271), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n757), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n756), .B1(new_n1091), .B2(new_n768), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1083), .B(new_n1092), .C1(new_n689), .C2(new_n753), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1061), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1060), .A2(new_n1094), .ZN(G393));
  INV_X1    g0895(.A(new_n1026), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1012), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1019), .A2(new_n691), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n701), .A3(new_n1027), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT115), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1016), .A2(new_n1020), .A3(KEYINPUT115), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n745), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1007), .A2(new_n752), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n829), .A2(new_n831), .B1(new_n784), .B2(new_n793), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT51), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n780), .A2(new_n271), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(new_n256), .B2(new_n827), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1107), .B(new_n1109), .C1(new_n201), .C2(new_n778), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n351), .B1(new_n797), .B2(G143), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n1111), .B1(new_n369), .B2(new_n786), .C1(new_n565), .C2(new_n774), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT116), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G317), .A2(new_n772), .B1(new_n796), .B2(G311), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT52), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n351), .B1(new_n783), .B2(new_n1065), .C1(new_n807), .C2(new_n791), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n778), .A2(new_n469), .B1(new_n774), .B2(new_n301), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n780), .A2(new_n492), .B1(new_n786), .B2(new_n808), .ZN(new_n1119));
  NOR4_X1   g0919(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n767), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n768), .B1(new_n488), .B2(new_n207), .C1(new_n235), .C2(new_n758), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1105), .A2(new_n746), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1100), .A2(new_n1104), .A3(new_n1123), .ZN(G390));
  OAI211_X1 g0924(.A(new_n673), .B(new_n818), .C1(new_n710), .C2(new_n713), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n819), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n954), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n939), .A2(new_n966), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n820), .A2(new_n934), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n738), .A2(new_n954), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n965), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n823), .A2(new_n819), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT103), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n955), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n966), .B1(new_n1136), .B2(new_n954), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1129), .B(new_n1131), .C1(new_n1132), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n954), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n967), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1140), .A2(new_n965), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n879), .A2(new_n954), .A3(new_n1130), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1138), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n738), .A2(new_n1130), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n954), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1125), .A2(new_n819), .A3(new_n1131), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n879), .A2(new_n1130), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n1145), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1136), .A2(new_n1147), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n969), .A2(new_n880), .A3(new_n664), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1143), .A2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1138), .B(new_n1157), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n701), .A3(new_n1158), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1143), .A2(new_n744), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n850), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n746), .B1(new_n1161), .B2(new_n256), .ZN(new_n1162));
  INV_X1    g0962(.A(G125), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n268), .B1(new_n783), .B2(new_n1163), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n778), .A2(new_n830), .B1(new_n201), .B2(new_n774), .ZN(new_n1165));
  INV_X1    g0965(.A(G128), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n829), .A2(new_n1166), .B1(new_n784), .B2(new_n780), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT54), .B(G143), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n793), .A2(new_n837), .B1(new_n791), .B2(new_n1168), .ZN(new_n1169));
  OR4_X1    g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n786), .A2(new_n1075), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT53), .Z(new_n1172));
  AOI21_X1  g0972(.A(new_n1108), .B1(G283), .B2(new_n772), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n301), .B2(new_n778), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n791), .A2(new_n488), .B1(new_n783), .B2(new_n807), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n268), .B(new_n1175), .C1(G116), .C2(new_n796), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(new_n788), .A3(new_n836), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1170), .A2(new_n1172), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1162), .B1(new_n1178), .B2(new_n767), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1132), .B2(new_n751), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1159), .A2(new_n1160), .A3(new_n1180), .ZN(G378));
  NAND2_X1  g0981(.A1(new_n329), .A2(new_n885), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n663), .A2(new_n338), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n299), .A2(new_n335), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n329), .B(new_n885), .C1(new_n1184), .C2(new_n657), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1186), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n933), .B2(new_n934), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n967), .B1(new_n961), .B2(new_n964), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(new_n959), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1189), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n950), .A2(G330), .A3(new_n1193), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1190), .A2(new_n958), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1193), .B1(new_n950), .B2(G330), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n934), .B(new_n1189), .C1(new_n943), .C2(new_n949), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n968), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1195), .A2(new_n1198), .A3(KEYINPUT119), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT119), .B1(new_n1195), .B2(new_n1198), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1158), .A2(new_n1154), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(KEYINPUT57), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n701), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1203), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n756), .B1(new_n201), .B2(new_n850), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n767), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n1163), .A2(new_n829), .B1(new_n778), .B2(new_n837), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n796), .A2(G128), .B1(new_n827), .B2(G137), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n786), .B2(new_n1168), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n780), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1210), .B(new_n1212), .C1(G150), .C2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n784), .B2(new_n774), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT118), .Z(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1220), .ZN(new_n1221));
  OAI22_X1  g1021(.A1(new_n829), .A2(new_n492), .B1(new_n774), .B2(new_n792), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G97), .B2(new_n777), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n351), .A2(new_n472), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G283), .B2(new_n797), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n791), .A2(new_n318), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(G107), .B2(new_n796), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1213), .A2(G68), .B1(new_n787), .B2(G77), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1223), .A2(new_n1225), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT58), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1224), .B(new_n251), .C1(G33), .C2(G41), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(KEYINPUT117), .ZN(new_n1234));
  AND4_X1   g1034(.A1(new_n1221), .A2(new_n1231), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n1208), .B1(new_n1209), .B2(new_n1235), .C1(new_n1193), .C2(new_n751), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1201), .B2(new_n745), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1207), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(G375));
  AND2_X1   g1041(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT120), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT120), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1245), .A3(new_n1054), .A4(new_n1155), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n756), .B1(new_n369), .B2(new_n850), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n351), .B1(new_n774), .B2(new_n271), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT121), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n791), .A2(new_n301), .B1(new_n783), .B2(new_n469), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(G283), .B2(new_n796), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1078), .B1(G116), .B2(new_n777), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n772), .A2(G294), .B1(new_n787), .B2(G97), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .A4(new_n1253), .ZN(new_n1254));
  OAI22_X1  g1054(.A1(new_n837), .A2(new_n829), .B1(new_n778), .B2(new_n1168), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n268), .B1(new_n791), .B2(new_n831), .C1(new_n830), .C2(new_n793), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n780), .A2(new_n251), .B1(new_n774), .B2(new_n792), .ZN(new_n1257));
  OR3_X1    g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n786), .A2(new_n784), .B1(new_n783), .B2(new_n1166), .ZN(new_n1259));
  XOR2_X1   g1059(.A(new_n1259), .B(KEYINPUT122), .Z(new_n1260));
  OAI21_X1  g1060(.A(new_n1254), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(KEYINPUT123), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n767), .ZN(new_n1264));
  OAI221_X1 g1064(.A(new_n1247), .B1(new_n1262), .B2(new_n1264), .C1(new_n954), .C2(new_n751), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1151), .B2(new_n744), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1246), .A2(new_n1267), .ZN(G381));
  NAND3_X1  g1068(.A1(new_n1030), .A2(new_n1051), .A3(new_n1002), .ZN(new_n1269));
  OAI21_X1  g1069(.A(KEYINPUT111), .B1(new_n1055), .B2(new_n1050), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1060), .A2(new_n814), .A3(new_n1094), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(G390), .A2(G381), .A3(new_n1272), .A4(G384), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1273), .A3(new_n1001), .ZN(new_n1274));
  XOR2_X1   g1074(.A(new_n1274), .B(KEYINPUT124), .Z(new_n1275));
  OR3_X1    g1075(.A1(new_n1275), .A2(G378), .A3(G375), .ZN(G407));
  INV_X1    g1076(.A(G378), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1240), .A2(new_n671), .A3(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(G407), .A2(G213), .A3(new_n1278), .ZN(G409));
  OAI211_X1 g1079(.A(G378), .B(new_n1238), .C1(new_n1203), .C2(new_n1206), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1237), .B1(new_n1204), .B2(new_n745), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT119), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1204), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1195), .A2(new_n1198), .A3(KEYINPUT119), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1202), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1285), .B2(new_n1029), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1277), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1280), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n671), .A2(G213), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1155), .A2(KEYINPUT60), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(new_n1245), .A3(new_n1243), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n702), .B1(new_n1242), .B2(KEYINPUT60), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G384), .B1(new_n1294), .B2(new_n1267), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n853), .B(new_n1266), .C1(new_n1292), .C2(new_n1293), .ZN(new_n1296));
  NOR2_X1   g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n671), .A2(G213), .A3(G2897), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1297), .B(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1100), .A2(new_n1104), .A3(new_n1123), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(G387), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1271), .A2(new_n1001), .A3(G390), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(G393), .A2(G396), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1272), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AND2_X1   g1107(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1303), .B(new_n1304), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(G390), .B1(new_n1271), .B2(new_n1001), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1001), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n1312), .B(new_n1302), .C1(new_n1269), .C2(new_n1270), .ZN(new_n1313));
  OAI22_X1  g1113(.A1(new_n1311), .A2(new_n1313), .B1(KEYINPUT125), .B2(new_n1307), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1310), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1288), .A2(new_n1297), .A3(new_n1289), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT63), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n1280), .A2(new_n1287), .B1(G213), .B2(new_n671), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(KEYINPUT63), .A3(new_n1297), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1301), .A2(new_n1315), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  AND4_X1   g1121(.A1(KEYINPUT62), .A2(new_n1288), .A3(new_n1297), .A4(new_n1289), .ZN(new_n1322));
  AOI21_X1  g1122(.A(KEYINPUT62), .B1(new_n1319), .B2(new_n1297), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1301), .B(KEYINPUT126), .C1(new_n1322), .C2(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(new_n1306), .B(KEYINPUT125), .ZN(new_n1325));
  NOR3_X1   g1125(.A1(new_n1311), .A2(new_n1313), .A3(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1309), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT127), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT127), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1310), .A2(new_n1314), .A3(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1324), .A2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT62), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1316), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1319), .A2(KEYINPUT62), .A3(new_n1297), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT126), .B1(new_n1336), .B2(new_n1301), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1321), .B1(new_n1332), .B2(new_n1337), .ZN(G405));
  NAND2_X1  g1138(.A1(G375), .A2(new_n1277), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(new_n1280), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1297), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1339), .B(new_n1280), .C1(new_n1295), .C2(new_n1296), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(new_n1331), .ZN(new_n1344));
  NAND4_X1  g1144(.A1(new_n1341), .A2(new_n1328), .A3(new_n1342), .A4(new_n1330), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(G402));
endmodule


