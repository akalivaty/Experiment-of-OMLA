//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n774, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n934, new_n935, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  OR2_X1    g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n203), .A2(new_n204), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT14), .ZN(new_n207));
  INV_X1    g006(.A(G29gat), .ZN(new_n208));
  INV_X1    g007(.A(G36gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n210), .A2(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n205), .A2(new_n206), .A3(new_n212), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n212), .A2(new_n204), .A3(new_n203), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n215), .B(KEYINPUT17), .ZN(new_n216));
  XOR2_X1   g015(.A(G15gat), .B(G22gat), .Z(new_n217));
  INV_X1    g016(.A(G1gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT84), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT16), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G1gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n220), .A2(new_n224), .A3(G8gat), .ZN(new_n225));
  INV_X1    g024(.A(G8gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n219), .B(new_n223), .C1(KEYINPUT84), .C2(new_n226), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n215), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n233), .B(KEYINPUT85), .Z(new_n234));
  OAI21_X1  g033(.A(new_n202), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(KEYINPUT11), .B(G169gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(G113gat), .B(G141gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n228), .A2(new_n230), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n234), .B(KEYINPUT86), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n243), .B(KEYINPUT13), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n234), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n229), .A2(KEYINPUT18), .A3(new_n231), .A4(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n235), .A2(new_n240), .A3(new_n245), .A4(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  INV_X1    g051(.A(new_n240), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n245), .A3(new_n247), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n251), .A2(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(G113gat), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G120gat), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT1), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(G134gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G127gat), .ZN(new_n262));
  INV_X1    g061(.A(G127gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G134gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n261), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n270), .B2(new_n260), .ZN(new_n271));
  NAND2_X1  g070(.A1(G183gat), .A2(G190gat), .ZN(new_n272));
  OR2_X1    g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT26), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n276));
  AND2_X1   g075(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT65), .B(G190gat), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT27), .B(G183gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT28), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n275), .B1(new_n281), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n274), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n273), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT64), .B1(new_n294), .B2(KEYINPUT23), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n296), .A3(new_n292), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n293), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n272), .B(KEYINPUT24), .ZN(new_n299));
  INV_X1    g098(.A(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n282), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT25), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n289), .A2(new_n291), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(new_n280), .B2(G183gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n284), .A2(G190gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n282), .A2(KEYINPUT65), .ZN(new_n307));
  OAI211_X1 g106(.A(KEYINPUT66), .B(new_n300), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n305), .A2(new_n299), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(new_n298), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT25), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n271), .B1(new_n303), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n275), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n286), .A2(new_n287), .A3(KEYINPUT28), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT28), .B1(new_n286), .B2(new_n287), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n291), .B(new_n313), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n302), .A2(new_n298), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT25), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(new_n309), .B2(new_n298), .ZN(new_n320));
  INV_X1    g119(.A(new_n271), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G227gat), .ZN(new_n324));
  INV_X1    g123(.A(G233gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT69), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(KEYINPUT34), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n326), .B1(new_n312), .B2(new_n322), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT33), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n321), .B1(new_n318), .B2(new_n320), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n303), .A2(new_n311), .A3(new_n271), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n327), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(KEYINPUT68), .B1(new_n337), .B2(KEYINPUT33), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(KEYINPUT32), .ZN(new_n339));
  XNOR2_X1  g138(.A(G15gat), .B(G43gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(G71gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n341), .B(G99gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n334), .A2(new_n338), .A3(new_n339), .A4(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n331), .B(KEYINPUT32), .C1(new_n333), .C2(new_n342), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n323), .A2(KEYINPUT69), .A3(new_n327), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n346), .B1(new_n344), .B2(new_n345), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n330), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n344), .A2(new_n345), .ZN(new_n350));
  INV_X1    g149(.A(new_n346), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(new_n353), .A3(new_n329), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n349), .A2(new_n354), .A3(KEYINPUT36), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT36), .B1(new_n349), .B2(new_n354), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(G50gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n359), .B(G78gat), .ZN(new_n360));
  INV_X1    g159(.A(G106gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n362), .B(KEYINPUT81), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  INV_X1    g163(.A(G211gat), .ZN(new_n365));
  INV_X1    g164(.A(G218gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n364), .B1(KEYINPUT22), .B2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G211gat), .B(G218gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT2), .ZN(new_n375));
  INV_X1    g174(.A(G141gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(G148gat), .ZN(new_n377));
  INV_X1    g176(.A(G148gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(G141gat), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n375), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n378), .B2(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(G141gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(KEYINPUT73), .A3(G148gat), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G155gat), .ZN(new_n386));
  INV_X1    g185(.A(G162gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n371), .B1(new_n388), .B2(KEYINPUT2), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n374), .A2(new_n380), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT3), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT74), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n385), .A2(new_n389), .ZN(new_n393));
  XNOR2_X1  g192(.A(G141gat), .B(G148gat), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n374), .B1(new_n394), .B2(KEYINPUT2), .ZN(new_n395));
  AND4_X1   g194(.A1(KEYINPUT74), .A2(new_n393), .A3(new_n395), .A4(new_n391), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n370), .B1(new_n397), .B2(KEYINPUT29), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n391), .B1(new_n370), .B2(KEYINPUT29), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n395), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n402), .A2(G22gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT80), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n406), .A2(G228gat), .A3(G233gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n403), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n407), .B1(new_n403), .B2(new_n404), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n363), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n403), .A2(new_n404), .ZN(new_n412));
  INV_X1    g211(.A(new_n407), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n362), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n416), .A3(new_n408), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT29), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n419), .B1(new_n318), .B2(new_n320), .ZN(new_n420));
  INV_X1    g219(.A(G226gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(new_n325), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT70), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n423), .B1(new_n303), .B2(new_n311), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n423), .B2(new_n420), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n370), .B(new_n425), .C1(new_n427), .C2(KEYINPUT70), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n422), .B1(new_n318), .B2(new_n320), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n370), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G8gat), .B(G36gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G92gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT71), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(G64gat), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(KEYINPUT30), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT70), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n420), .B2(new_n423), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT29), .B1(new_n303), .B2(new_n311), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n429), .B1(new_n441), .B2(new_n422), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(new_n439), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n430), .B1(new_n443), .B2(new_n370), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n436), .ZN(new_n445));
  AND2_X1   g244(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT72), .B1(new_n444), .B2(new_n436), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n432), .A2(new_n449), .A3(new_n437), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n446), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n261), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n265), .B2(KEYINPUT67), .ZN(new_n454));
  INV_X1    g253(.A(new_n260), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n400), .A2(new_n456), .A3(new_n266), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n271), .A2(new_n390), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n271), .A2(new_n462), .A3(new_n390), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT77), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n458), .A2(KEYINPUT4), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n464), .A3(KEYINPUT4), .ZN(new_n468));
  INV_X1    g267(.A(new_n396), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n470), .B1(new_n400), .B2(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n391), .B1(new_n393), .B2(new_n395), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n271), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n467), .A2(new_n468), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT39), .B(new_n461), .C1(new_n475), .C2(new_n460), .ZN(new_n476));
  XOR2_X1   g275(.A(G1gat), .B(G29gat), .Z(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G57gat), .B(G85gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n474), .B1(new_n392), .B2(new_n396), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n462), .B1(new_n271), .B2(new_n390), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n483), .B1(new_n464), .B2(new_n463), .ZN(new_n484));
  INV_X1    g283(.A(new_n468), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT39), .ZN(new_n487));
  INV_X1    g286(.A(new_n460), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n476), .A2(KEYINPUT40), .A3(new_n481), .A4(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT82), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g291(.A1(new_n489), .A2(new_n481), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n493), .A2(KEYINPUT82), .A3(KEYINPUT40), .A4(new_n476), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT75), .B(KEYINPUT5), .C1(new_n459), .C2(new_n460), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n466), .A2(new_n463), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n482), .A3(new_n460), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT75), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n460), .B1(new_n457), .B2(new_n458), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT5), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n482), .B(new_n504), .C1(new_n484), .C2(new_n485), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n481), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n493), .A2(new_n476), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n495), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n452), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n447), .A2(new_n450), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n436), .B1(new_n444), .B2(KEYINPUT37), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT37), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n432), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT38), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT83), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n506), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n503), .A2(new_n505), .A3(new_n481), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n506), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n519), .A2(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n437), .B1(new_n432), .B2(new_n514), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n427), .A2(new_n370), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(KEYINPUT37), .C1(new_n443), .C2(new_n370), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n512), .A2(new_n516), .A3(new_n524), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n418), .B1(new_n511), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT78), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n522), .A2(new_n532), .A3(new_n523), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n503), .A2(new_n505), .ZN(new_n534));
  INV_X1    g333(.A(new_n481), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n503), .A2(new_n505), .A3(new_n481), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n523), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(KEYINPUT78), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n533), .A2(new_n539), .A3(new_n517), .ZN(new_n540));
  AND4_X1   g339(.A1(new_n540), .A2(new_n418), .A3(new_n451), .A4(new_n446), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n357), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n411), .A2(new_n417), .ZN(new_n543));
  NOR3_X1   g342(.A1(new_n347), .A2(new_n348), .A3(new_n330), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n329), .B1(new_n352), .B2(new_n353), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n540), .A2(new_n451), .A3(new_n446), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT35), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n418), .B1(new_n349), .B2(new_n354), .ZN(new_n549));
  AND2_X1   g348(.A1(new_n446), .A2(new_n451), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n524), .A2(KEYINPUT35), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n255), .B1(new_n542), .B2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(G190gat), .B(G218gat), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT91), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g357(.A1(G85gat), .A2(G92gat), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n558), .B(new_n559), .Z(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT93), .B(G92gat), .ZN(new_n561));
  INV_X1    g360(.A(G85gat), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G99gat), .ZN(new_n564));
  OR3_X1    g363(.A1(new_n564), .A2(new_n361), .A3(KEYINPUT92), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT92), .B1(new_n564), .B2(new_n361), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(KEYINPUT8), .A3(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n560), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n560), .A2(new_n569), .A3(new_n563), .A4(new_n567), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n215), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT90), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT94), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n573), .A2(KEYINPUT94), .A3(new_n577), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n571), .A2(new_n572), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n216), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n556), .B1(new_n585), .B2(KEYINPUT95), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n576), .A2(KEYINPUT41), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g388(.A1(new_n580), .A2(new_n581), .B1(new_n216), .B2(new_n583), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT95), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n555), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n592), .A2(new_n587), .ZN(new_n593));
  XOR2_X1   g392(.A(G134gat), .B(G162gat), .Z(new_n594));
  NOR3_X1   g393(.A1(new_n589), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n586), .A2(new_n588), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n592), .A2(new_n587), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n590), .A2(new_n591), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n595), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n594), .B1(new_n589), .B2(new_n593), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n598), .A3(new_n596), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(new_n365), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT9), .ZN(new_n610));
  INV_X1    g409(.A(G71gat), .ZN(new_n611));
  INV_X1    g410(.A(G78gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT88), .ZN(new_n614));
  XOR2_X1   g413(.A(G57gat), .B(G64gat), .Z(new_n615));
  INV_X1    g414(.A(KEYINPUT88), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n616), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(G71gat), .B(G78gat), .Z(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n228), .B1(new_n609), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G183gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT89), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n623), .B(new_n300), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT89), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(G231gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n325), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n625), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n625), .B2(new_n628), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n608), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n625), .A2(new_n628), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n625), .A2(new_n628), .A3(new_n630), .ZN(new_n637));
  INV_X1    g436(.A(new_n608), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n636), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n609), .ZN(new_n640));
  XOR2_X1   g439(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AND3_X1   g441(.A1(new_n633), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n633), .B2(new_n639), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n583), .A2(new_n622), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT10), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n571), .A2(new_n621), .A3(new_n620), .A4(new_n572), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n650), .A2(new_n649), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n647), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n646), .B1(new_n648), .B2(new_n650), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G120gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n378), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT98), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n655), .A2(new_n659), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n660), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n663), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n664), .B1(new_n663), .B2(new_n666), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n606), .A2(new_n645), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n606), .A2(new_n645), .A3(KEYINPUT99), .A4(new_n669), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n554), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n540), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(new_n218), .ZN(G1324gat));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n550), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n222), .A2(new_n226), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n679), .B1(new_n222), .B2(new_n226), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n682), .B(new_n683), .C1(new_n226), .C2(new_n677), .ZN(G1325gat));
  OAI21_X1  g483(.A(KEYINPUT101), .B1(new_n355), .B2(new_n356), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT36), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n544), .B2(new_n545), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n349), .A2(new_n354), .A3(KEYINPUT36), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT102), .ZN(new_n692));
  INV_X1    g491(.A(G15gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n674), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n349), .A2(new_n354), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n674), .B2(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(KEYINPUT100), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n694), .B1(new_n698), .B2(new_n699), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n674), .A2(new_n543), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n511), .A2(new_n530), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n541), .B1(new_n704), .B2(new_n543), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n553), .B1(new_n691), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n600), .B1(new_n595), .B2(new_n599), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n603), .A2(new_n602), .A3(new_n604), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n711), .B(new_n606), .C1(new_n542), .C2(new_n553), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n254), .A2(new_n253), .ZN(new_n714));
  INV_X1    g513(.A(new_n252), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n250), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n645), .A2(KEYINPUT104), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n645), .A2(KEYINPUT104), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n716), .B(new_n669), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT105), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n713), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT106), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G29gat), .B1(new_n723), .B2(new_n540), .ZN(new_n724));
  INV_X1    g523(.A(new_n645), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n669), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n554), .A2(new_n709), .A3(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n728), .A2(G29gat), .A3(new_n540), .ZN(new_n729));
  XNOR2_X1  g528(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n724), .A2(new_n731), .ZN(G1328gat));
  OAI21_X1  g531(.A(G36gat), .B1(new_n723), .B2(new_n550), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n728), .A2(G36gat), .A3(new_n550), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n735), .A2(KEYINPUT107), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n733), .B(new_n738), .C1(new_n736), .C2(new_n734), .ZN(G1329gat));
  INV_X1    g538(.A(new_n691), .ZN(new_n740));
  OAI211_X1 g539(.A(KEYINPUT47), .B(G43gat), .C1(new_n721), .C2(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n728), .A2(G43gat), .A3(new_n696), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n741), .B(new_n743), .C1(KEYINPUT108), .C2(KEYINPUT47), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n745));
  INV_X1    g544(.A(new_n692), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n722), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n745), .B1(new_n747), .B2(G43gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n748), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g548(.A(G50gat), .B1(new_n721), .B2(new_n543), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n728), .A2(G50gat), .A3(new_n543), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n750), .A2(KEYINPUT48), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n722), .A2(new_n418), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n751), .B1(new_n754), .B2(G50gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(KEYINPUT48), .ZN(G1331gat));
  OAI211_X1 g555(.A(new_n685), .B(new_n690), .C1(new_n531), .C2(new_n541), .ZN(new_n757));
  AOI211_X1 g556(.A(new_n725), .B(new_n709), .C1(new_n757), .C2(new_n553), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n669), .A2(new_n716), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  AND3_X1   g560(.A1(new_n533), .A2(new_n539), .A3(new_n517), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n760), .A2(new_n550), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  NAND3_X1  g568(.A1(new_n761), .A2(new_n611), .A3(new_n695), .ZN(new_n770));
  OAI21_X1  g569(.A(G71gat), .B1(new_n760), .B2(new_n692), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g572(.A1(new_n760), .A2(new_n543), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(new_n612), .ZN(G1335gat));
  NAND2_X1  g574(.A1(new_n687), .A2(new_n689), .ZN(new_n776));
  AND4_X1   g575(.A1(new_n512), .A2(new_n516), .A3(new_n524), .A4(new_n529), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n495), .A2(new_n509), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n451), .B2(new_n446), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n543), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(new_n541), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT35), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n762), .A2(new_n452), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n549), .ZN(new_n785));
  AND4_X1   g584(.A1(new_n695), .A2(new_n550), .A3(new_n543), .A4(new_n551), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT44), .B(new_n709), .C1(new_n782), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n255), .B1(new_n643), .B2(new_n644), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(KEYINPUT109), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n669), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n606), .B1(new_n757), .B2(new_n553), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n788), .B(new_n792), .C1(new_n793), .C2(KEYINPUT44), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n794), .A2(new_n562), .A3(new_n540), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n790), .A2(new_n791), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n706), .A2(new_n796), .A3(new_n709), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(KEYINPUT51), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n793), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n669), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n762), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n795), .B1(new_n803), .B2(new_n562), .ZN(G1336gat));
  NOR2_X1   g603(.A1(new_n550), .A2(G92gat), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n798), .A2(new_n802), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n794), .A2(new_n550), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n561), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT110), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n808), .B(new_n809), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(KEYINPUT52), .ZN(G1337gat));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n692), .ZN(new_n812));
  XOR2_X1   g611(.A(new_n812), .B(KEYINPUT111), .Z(new_n813));
  NAND2_X1  g612(.A1(new_n801), .A2(new_n802), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n695), .A2(new_n564), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n813), .A2(new_n564), .B1(new_n814), .B2(new_n815), .ZN(G1338gat));
  XNOR2_X1  g615(.A(KEYINPUT112), .B(G106gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n794), .B2(new_n543), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n543), .A2(G106gat), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n798), .A2(new_n802), .A3(new_n800), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT53), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n713), .A2(KEYINPUT113), .A3(new_n418), .A4(new_n792), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n794), .B2(new_n543), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n817), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n826), .A2(new_n828), .A3(KEYINPUT114), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT114), .B1(new_n826), .B2(new_n828), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n822), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT115), .B(new_n822), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(G1339gat));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n651), .A2(new_n652), .A3(new_n647), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT54), .B1(new_n837), .B2(KEYINPUT116), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n651), .A2(new_n652), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n646), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(new_n837), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n659), .B1(new_n653), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n836), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n837), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n848), .B1(new_n841), .B2(new_n840), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n845), .B(KEYINPUT55), .C1(new_n849), .C2(new_n838), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(new_n660), .A3(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n847), .A2(new_n850), .A3(KEYINPUT117), .A4(new_n660), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n716), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n232), .A2(new_n234), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n242), .A2(new_n244), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n239), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n251), .B2(new_n252), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n667), .B2(new_n668), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n606), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n601), .B2(new_n605), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n853), .A2(new_n854), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT118), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n717), .A2(new_n718), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n709), .B1(new_n855), .B2(new_n860), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n863), .A2(new_n864), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n866), .A2(new_n867), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n670), .A2(new_n716), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n546), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n452), .A2(new_n540), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n255), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(new_n258), .ZN(G1340gat));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n669), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(new_n256), .ZN(G1341gat));
  NOR3_X1   g679(.A1(new_n876), .A2(new_n263), .A3(new_n867), .ZN(new_n881));
  INV_X1    g680(.A(new_n876), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n645), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n263), .B2(new_n883), .ZN(G1342gat));
  NOR2_X1   g683(.A1(new_n876), .A2(new_n606), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n261), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(KEYINPUT56), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n887), .B(new_n888), .C1(new_n261), .C2(new_n885), .ZN(G1343gat));
  INV_X1    g688(.A(new_n851), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n716), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n709), .B1(new_n860), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n870), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n873), .B1(new_n893), .B2(new_n645), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(KEYINPUT57), .A3(new_n418), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n543), .B1(new_n872), .B2(new_n873), .ZN(new_n896));
  XNOR2_X1  g695(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n740), .A2(new_n875), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n898), .A2(G141gat), .A3(new_n716), .A4(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n896), .A2(new_n716), .A3(new_n692), .A4(new_n875), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n376), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(KEYINPUT58), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT58), .B1(new_n901), .B2(new_n903), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT121), .B(KEYINPUT58), .C1(new_n901), .C2(new_n903), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n906), .A2(new_n907), .B1(new_n910), .B2(new_n911), .ZN(G1344gat));
  AND2_X1   g711(.A1(new_n896), .A2(new_n692), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n913), .A2(new_n875), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n378), .A3(new_n802), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n898), .A2(new_n900), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n378), .C1(new_n916), .C2(new_n802), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n672), .A2(new_n255), .A3(new_n673), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n709), .A2(new_n890), .A3(new_n859), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n725), .B1(new_n921), .B2(new_n892), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n543), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  OR3_X1    g722(.A1(new_n923), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n896), .A2(new_n897), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT122), .B1(new_n923), .B2(KEYINPUT57), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n802), .A3(new_n900), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n918), .B1(new_n928), .B2(G148gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n915), .B1(new_n917), .B2(new_n929), .ZN(G1345gat));
  AOI21_X1  g729(.A(G155gat), .B1(new_n914), .B2(new_n645), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n867), .A2(new_n386), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n931), .B1(new_n916), .B2(new_n932), .ZN(G1346gat));
  AOI21_X1  g732(.A(G162gat), .B1(new_n914), .B2(new_n709), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n606), .A2(new_n387), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n916), .B2(new_n935), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n550), .A2(new_n762), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n874), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(G169gat), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n939), .A2(new_n940), .A3(new_n716), .ZN(new_n941));
  XOR2_X1   g740(.A(new_n937), .B(KEYINPUT123), .Z(new_n942));
  OR2_X1    g741(.A1(new_n942), .A2(new_n696), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n872), .A2(new_n873), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n418), .B1(new_n943), .B2(KEYINPUT124), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n947), .A2(new_n716), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n941), .B1(new_n948), .B2(new_n940), .ZN(G1348gat));
  NAND3_X1  g748(.A1(new_n947), .A2(G176gat), .A3(new_n802), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  AOI21_X1  g750(.A(G176gat), .B1(new_n939), .B2(new_n802), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1349gat));
  NOR3_X1   g752(.A1(new_n938), .A2(new_n279), .A3(new_n725), .ZN(new_n954));
  INV_X1    g753(.A(new_n867), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n947), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n954), .B1(G183gat), .B2(new_n956), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g757(.A(new_n282), .B1(new_n947), .B2(new_n709), .ZN(new_n959));
  XOR2_X1   g758(.A(new_n959), .B(KEYINPUT61), .Z(new_n960));
  NAND3_X1  g759(.A1(new_n939), .A2(new_n286), .A3(new_n709), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n927), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n924), .A2(new_n925), .A3(new_n964), .A4(new_n926), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n746), .A2(new_n942), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G197gat), .B1(new_n967), .B2(new_n255), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n913), .A2(new_n937), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n969), .A2(G197gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n255), .B2(new_n970), .ZN(G1352gat));
  OAI21_X1  g770(.A(G204gat), .B1(new_n967), .B2(new_n669), .ZN(new_n972));
  OR3_X1    g771(.A1(new_n969), .A2(G204gat), .A3(new_n669), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT62), .ZN(new_n974));
  OR4_X1    g773(.A1(KEYINPUT62), .A2(new_n969), .A3(G204gat), .A4(new_n669), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n972), .A2(new_n974), .A3(new_n975), .ZN(G1353gat));
  NAND3_X1  g775(.A1(new_n927), .A2(new_n645), .A3(new_n966), .ZN(new_n977));
  NOR2_X1   g776(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n977), .A2(G211gat), .A3(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(new_n969), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n980), .A2(new_n365), .A3(new_n645), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n977), .A2(G211gat), .ZN(new_n982));
  XNOR2_X1  g781(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n979), .B(new_n981), .C1(new_n982), .C2(new_n983), .ZN(G1354gat));
  OAI21_X1  g783(.A(G218gat), .B1(new_n967), .B2(new_n606), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n980), .A2(new_n366), .A3(new_n709), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1355gat));
endmodule


