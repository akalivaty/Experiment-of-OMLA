

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775;

  NOR2_X1 U375 ( .A1(n737), .A2(n736), .ZN(n584) );
  XNOR2_X1 U376 ( .A(n533), .B(n352), .ZN(n563) );
  XNOR2_X1 U377 ( .A(KEYINPUT73), .B(KEYINPUT22), .ZN(n352) );
  XNOR2_X2 U378 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n468) );
  NOR2_X2 U379 ( .A1(n775), .A2(n657), .ZN(n379) );
  NOR2_X1 U380 ( .A1(n723), .A2(n612), .ZN(n416) );
  XNOR2_X2 U381 ( .A(n568), .B(n463), .ZN(n615) );
  XNOR2_X2 U382 ( .A(n364), .B(n365), .ZN(n568) );
  INV_X1 U383 ( .A(n603), .ZN(n627) );
  INV_X1 U384 ( .A(KEYINPUT64), .ZN(n404) );
  OR2_X1 U385 ( .A1(n708), .A2(n707), .ZN(n392) );
  NAND2_X1 U386 ( .A1(n407), .A2(n711), .ZN(n406) );
  BUF_X1 U387 ( .A(n704), .Z(n766) );
  XNOR2_X1 U388 ( .A(n633), .B(KEYINPUT82), .ZN(n704) );
  AND2_X1 U389 ( .A1(n632), .A2(n631), .ZN(n633) );
  AND2_X1 U390 ( .A1(n380), .A2(n378), .ZN(n623) );
  AND2_X1 U391 ( .A1(n590), .A2(n605), .ZN(n595) );
  AND2_X1 U392 ( .A1(n534), .A2(n538), .ZN(n539) );
  INV_X1 U393 ( .A(n363), .ZN(n534) );
  NAND2_X2 U394 ( .A1(n401), .A2(n398), .ZN(n605) );
  XNOR2_X1 U395 ( .A(n450), .B(n449), .ZN(n588) );
  AND2_X1 U396 ( .A1(n403), .A2(n402), .ZN(n401) );
  XNOR2_X1 U397 ( .A(n374), .B(n423), .ZN(n355) );
  NAND2_X1 U398 ( .A1(n353), .A2(n363), .ZN(n465) );
  XNOR2_X2 U399 ( .A(n605), .B(KEYINPUT1), .ZN(n363) );
  NOR2_X1 U400 ( .A1(n615), .A2(n713), .ZN(n353) );
  NAND2_X1 U401 ( .A1(n360), .A2(n361), .ZN(n359) );
  INV_X1 U402 ( .A(n354), .ZN(n752) );
  NAND2_X1 U403 ( .A1(n634), .A2(n354), .ZN(n706) );
  XNOR2_X2 U404 ( .A(n359), .B(n567), .ZN(n354) );
  NAND2_X1 U405 ( .A1(n354), .A2(n704), .ZN(n407) );
  NAND2_X1 U406 ( .A1(n710), .A2(n354), .ZN(n712) );
  NAND2_X1 U407 ( .A1(n355), .A2(n435), .ZN(n403) );
  OR2_X1 U408 ( .A1(n355), .A2(n399), .ZN(n398) );
  XNOR2_X1 U409 ( .A(n355), .B(n682), .ZN(n683) );
  NAND2_X1 U410 ( .A1(n662), .A2(n658), .ZN(n544) );
  NAND2_X1 U411 ( .A1(n563), .A2(n539), .ZN(n658) );
  XNOR2_X2 U412 ( .A(n356), .B(KEYINPUT32), .ZN(n662) );
  NAND2_X1 U413 ( .A1(n563), .A2(n357), .ZN(n356) );
  AND2_X1 U414 ( .A1(n536), .A2(n615), .ZN(n357) );
  AND2_X1 U415 ( .A1(n358), .A2(n545), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n543), .B(KEYINPUT70), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n362), .B(KEYINPUT86), .ZN(n361) );
  NOR2_X2 U418 ( .A1(n566), .A2(n565), .ZN(n362) );
  NOR2_X1 U419 ( .A1(n664), .A2(G902), .ZN(n364) );
  XOR2_X1 U420 ( .A(n462), .B(G472), .Z(n365) );
  NOR2_X2 U421 ( .A1(n663), .A2(KEYINPUT44), .ZN(n542) );
  NOR2_X1 U422 ( .A1(n738), .A2(n397), .ZN(n396) );
  OR2_X1 U423 ( .A1(n588), .A2(n587), .ZN(n612) );
  INV_X1 U424 ( .A(KEYINPUT0), .ZN(n376) );
  XNOR2_X1 U425 ( .A(n505), .B(n419), .ZN(n512) );
  AND2_X1 U426 ( .A1(n388), .A2(n410), .ZN(n386) );
  INV_X1 U427 ( .A(n392), .ZN(n388) );
  XNOR2_X1 U428 ( .A(n395), .B(n394), .ZN(n393) );
  INV_X1 U429 ( .A(KEYINPUT47), .ZN(n394) );
  AND2_X1 U430 ( .A1(n381), .A2(n622), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n382), .B(n611), .ZN(n381) );
  INV_X1 U432 ( .A(G237), .ZN(n483) );
  XNOR2_X1 U433 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n436) );
  NOR2_X1 U434 ( .A1(n618), .A2(n694), .ZN(n624) );
  NAND2_X1 U435 ( .A1(n400), .A2(n524), .ZN(n399) );
  XNOR2_X1 U436 ( .A(n639), .B(n638), .ZN(n640) );
  BUF_X1 U437 ( .A(n671), .Z(n680) );
  XNOR2_X1 U438 ( .A(n646), .B(n645), .ZN(n647) );
  NOR2_X1 U439 ( .A1(n750), .A2(n368), .ZN(n410) );
  NAND2_X1 U440 ( .A1(n390), .A2(n389), .ZN(n384) );
  NAND2_X1 U441 ( .A1(n392), .A2(n391), .ZN(n390) );
  XNOR2_X1 U442 ( .A(n379), .B(KEYINPUT46), .ZN(n378) );
  INV_X1 U443 ( .A(KEYINPUT88), .ZN(n540) );
  XNOR2_X1 U444 ( .A(G146), .B(G125), .ZN(n469) );
  NAND2_X1 U445 ( .A1(G234), .A2(G237), .ZN(n490) );
  XNOR2_X1 U446 ( .A(n506), .B(n420), .ZN(n419) );
  INV_X1 U447 ( .A(KEYINPUT101), .ZN(n420) );
  XNOR2_X1 U448 ( .A(KEYINPUT66), .B(G101), .ZN(n472) );
  XNOR2_X1 U449 ( .A(n484), .B(KEYINPUT78), .ZN(n485) );
  NAND2_X1 U450 ( .A1(n435), .A2(G902), .ZN(n402) );
  XNOR2_X1 U451 ( .A(G119), .B(G116), .ZN(n454) );
  XNOR2_X1 U452 ( .A(G107), .B(G104), .ZN(n430) );
  XNOR2_X1 U453 ( .A(n416), .B(n371), .ZN(n590) );
  XNOR2_X1 U454 ( .A(n514), .B(n513), .ZN(n556) );
  XOR2_X1 U455 ( .A(KEYINPUT62), .B(n665), .Z(n666) );
  XNOR2_X1 U456 ( .A(n444), .B(n765), .ZN(n672) );
  XNOR2_X1 U457 ( .A(n409), .B(n439), .ZN(n444) );
  XNOR2_X1 U458 ( .A(n442), .B(n438), .ZN(n409) );
  NAND2_X1 U459 ( .A1(n642), .A2(G953), .ZN(n675) );
  OR2_X1 U460 ( .A1(n621), .A2(n534), .ZN(n661) );
  XNOR2_X1 U461 ( .A(n549), .B(n422), .ZN(n698) );
  NOR2_X1 U462 ( .A1(n727), .A2(n529), .ZN(n549) );
  XNOR2_X1 U463 ( .A(n677), .B(n411), .ZN(n679) );
  INV_X1 U464 ( .A(n678), .ZN(n411) );
  INV_X1 U465 ( .A(KEYINPUT60), .ZN(n412) );
  INV_X1 U466 ( .A(KEYINPUT56), .ZN(n414) );
  NAND2_X1 U467 ( .A1(n384), .A2(n410), .ZN(n383) );
  NAND2_X1 U468 ( .A1(n386), .A2(n366), .ZN(n385) );
  AND2_X1 U469 ( .A1(n387), .A2(KEYINPUT81), .ZN(n366) );
  XOR2_X1 U470 ( .A(n417), .B(n370), .Z(n367) );
  OR2_X1 U471 ( .A1(G953), .A2(n703), .ZN(n368) );
  OR2_X1 U472 ( .A1(G953), .A2(G237), .ZN(n369) );
  XNOR2_X1 U473 ( .A(KEYINPUT85), .B(KEYINPUT39), .ZN(n370) );
  XOR2_X1 U474 ( .A(n589), .B(KEYINPUT28), .Z(n371) );
  XOR2_X1 U475 ( .A(KEYINPUT71), .B(KEYINPUT34), .Z(n372) );
  AND2_X1 U476 ( .A1(n711), .A2(n391), .ZN(n373) );
  INV_X1 U477 ( .A(KEYINPUT81), .ZN(n391) );
  BUF_X1 U478 ( .A(n568), .Z(n723) );
  INV_X1 U479 ( .A(n375), .ZN(n529) );
  INV_X1 U480 ( .A(n594), .ZN(n397) );
  XNOR2_X1 U481 ( .A(n764), .B(n428), .ZN(n374) );
  XNOR2_X1 U482 ( .A(n764), .B(n428), .ZN(n461) );
  XNOR2_X2 U483 ( .A(n497), .B(n376), .ZN(n375) );
  BUF_X1 U484 ( .A(n475), .Z(n377) );
  XNOR2_X1 U485 ( .A(n476), .B(n377), .ZN(n481) );
  NAND2_X2 U486 ( .A1(n408), .A2(n406), .ZN(n405) );
  NAND2_X1 U487 ( .A1(n610), .A2(n609), .ZN(n382) );
  NAND2_X1 U488 ( .A1(n385), .A2(n383), .ZN(n751) );
  NAND2_X1 U489 ( .A1(n712), .A2(n711), .ZN(n387) );
  NAND2_X1 U490 ( .A1(n712), .A2(n373), .ZN(n389) );
  NAND2_X1 U491 ( .A1(n393), .A2(n596), .ZN(n602) );
  NAND2_X1 U492 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U493 ( .A1(n595), .A2(n396), .ZN(n395) );
  INV_X1 U494 ( .A(n435), .ZN(n400) );
  XNOR2_X2 U495 ( .A(n405), .B(n404), .ZN(n671) );
  AND2_X2 U496 ( .A1(n706), .A2(n635), .ZN(n408) );
  XNOR2_X1 U497 ( .A(n528), .B(KEYINPUT35), .ZN(n546) );
  XNOR2_X1 U498 ( .A(n486), .B(n485), .ZN(n574) );
  BUF_X2 U499 ( .A(n546), .Z(n663) );
  BUF_X1 U500 ( .A(n574), .Z(n603) );
  XNOR2_X2 U501 ( .A(n627), .B(n575), .ZN(n734) );
  XNOR2_X1 U502 ( .A(n413), .B(n412), .ZN(G60) );
  NAND2_X1 U503 ( .A1(n643), .A2(n675), .ZN(n413) );
  XNOR2_X1 U504 ( .A(n415), .B(n414), .ZN(G51) );
  NAND2_X1 U505 ( .A1(n649), .A2(n675), .ZN(n415) );
  NAND2_X1 U506 ( .A1(n576), .A2(n577), .ZN(n417) );
  XNOR2_X1 U507 ( .A(n418), .B(KEYINPUT30), .ZN(n573) );
  NOR2_X1 U508 ( .A1(n568), .A2(n582), .ZN(n418) );
  XNOR2_X1 U509 ( .A(n421), .B(n372), .ZN(n527) );
  NOR2_X2 U510 ( .A1(n700), .A2(n529), .ZN(n421) );
  BUF_X1 U511 ( .A(n644), .Z(n646) );
  XNOR2_X1 U512 ( .A(KEYINPUT31), .B(KEYINPUT100), .ZN(n422) );
  XOR2_X1 U513 ( .A(n443), .B(n433), .Z(n423) );
  AND2_X1 U514 ( .A1(n715), .A2(n586), .ZN(n424) );
  INV_X1 U515 ( .A(KEYINPUT19), .ZN(n488) );
  NAND2_X1 U516 ( .A1(n573), .A2(n424), .ZN(n608) );
  XNOR2_X1 U517 ( .A(n674), .B(n673), .ZN(n676) );
  XNOR2_X2 U518 ( .A(G143), .B(KEYINPUT77), .ZN(n425) );
  XNOR2_X2 U519 ( .A(n425), .B(G128), .ZN(n521) );
  XNOR2_X2 U520 ( .A(n521), .B(KEYINPUT4), .ZN(n475) );
  XNOR2_X1 U521 ( .A(G134), .B(G131), .ZN(n426) );
  XNOR2_X1 U522 ( .A(n426), .B(KEYINPUT68), .ZN(n427) );
  XNOR2_X2 U523 ( .A(n475), .B(n427), .ZN(n764) );
  XNOR2_X1 U524 ( .A(n472), .B(G146), .ZN(n428) );
  XOR2_X1 U525 ( .A(G137), .B(G140), .Z(n443) );
  XNOR2_X1 U526 ( .A(KEYINPUT92), .B(G110), .ZN(n429) );
  XNOR2_X1 U527 ( .A(n430), .B(n429), .ZN(n478) );
  INV_X2 U528 ( .A(G953), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n466), .A2(G227), .ZN(n431) );
  XNOR2_X1 U530 ( .A(n431), .B(KEYINPUT96), .ZN(n432) );
  XNOR2_X1 U531 ( .A(n478), .B(n432), .ZN(n433) );
  INV_X1 U532 ( .A(KEYINPUT69), .ZN(n434) );
  XNOR2_X1 U533 ( .A(n434), .B(G469), .ZN(n435) );
  NAND2_X1 U534 ( .A1(n466), .A2(G234), .ZN(n437) );
  XNOR2_X1 U535 ( .A(n437), .B(n436), .ZN(n518) );
  NAND2_X1 U536 ( .A1(n518), .A2(G221), .ZN(n439) );
  XNOR2_X1 U537 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n438) );
  XOR2_X1 U538 ( .A(KEYINPUT97), .B(G110), .Z(n441) );
  XNOR2_X1 U539 ( .A(G119), .B(G128), .ZN(n440) );
  XNOR2_X1 U540 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U541 ( .A(KEYINPUT10), .B(n469), .ZN(n502) );
  XNOR2_X1 U542 ( .A(n502), .B(n443), .ZN(n765) );
  INV_X1 U543 ( .A(G902), .ZN(n524) );
  NAND2_X1 U544 ( .A1(n672), .A2(n524), .ZN(n450) );
  INV_X1 U545 ( .A(KEYINPUT15), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n445), .B(G902), .ZN(n635) );
  INV_X1 U547 ( .A(n635), .ZN(n482) );
  NAND2_X1 U548 ( .A1(G234), .A2(n482), .ZN(n446) );
  XNOR2_X1 U549 ( .A(KEYINPUT20), .B(n446), .ZN(n451) );
  NAND2_X1 U550 ( .A1(G217), .A2(n451), .ZN(n448) );
  INV_X1 U551 ( .A(KEYINPUT25), .ZN(n447) );
  XNOR2_X1 U552 ( .A(n448), .B(n447), .ZN(n449) );
  NAND2_X1 U553 ( .A1(n451), .A2(G221), .ZN(n452) );
  XNOR2_X1 U554 ( .A(n452), .B(KEYINPUT21), .ZN(n720) );
  INV_X1 U555 ( .A(KEYINPUT98), .ZN(n453) );
  XNOR2_X1 U556 ( .A(n720), .B(n453), .ZN(n530) );
  AND2_X1 U557 ( .A1(n588), .A2(n530), .ZN(n715) );
  INV_X1 U558 ( .A(n715), .ZN(n713) );
  XNOR2_X1 U559 ( .A(n454), .B(KEYINPUT3), .ZN(n456) );
  XNOR2_X1 U560 ( .A(G113), .B(KEYINPUT93), .ZN(n455) );
  XNOR2_X1 U561 ( .A(n456), .B(n455), .ZN(n479) );
  XNOR2_X1 U562 ( .A(KEYINPUT75), .B(n369), .ZN(n507) );
  NAND2_X1 U563 ( .A1(n507), .A2(G210), .ZN(n458) );
  XNOR2_X1 U564 ( .A(KEYINPUT5), .B(G137), .ZN(n457) );
  XNOR2_X1 U565 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U566 ( .A(n479), .B(n459), .ZN(n460) );
  XNOR2_X1 U567 ( .A(n461), .B(n460), .ZN(n664) );
  INV_X1 U568 ( .A(KEYINPUT72), .ZN(n462) );
  XNOR2_X1 U569 ( .A(KEYINPUT103), .B(KEYINPUT6), .ZN(n463) );
  INV_X1 U570 ( .A(KEYINPUT33), .ZN(n464) );
  XNOR2_X1 U571 ( .A(n465), .B(n464), .ZN(n700) );
  NAND2_X1 U572 ( .A1(n466), .A2(G224), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n468), .B(n467), .ZN(n470) );
  XNOR2_X1 U574 ( .A(n470), .B(n469), .ZN(n474) );
  XNOR2_X1 U575 ( .A(KEYINPUT76), .B(KEYINPUT89), .ZN(n471) );
  XNOR2_X1 U576 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U577 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U578 ( .A(KEYINPUT16), .B(G122), .ZN(n477) );
  XNOR2_X1 U579 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U580 ( .A(n480), .B(n479), .ZN(n759) );
  XNOR2_X1 U581 ( .A(n481), .B(n759), .ZN(n644) );
  NAND2_X1 U582 ( .A1(n644), .A2(n482), .ZN(n486) );
  NAND2_X1 U583 ( .A1(n524), .A2(n483), .ZN(n487) );
  NAND2_X1 U584 ( .A1(n487), .A2(G210), .ZN(n484) );
  AND2_X1 U585 ( .A1(n487), .A2(G214), .ZN(n582) );
  NOR2_X2 U586 ( .A1(n574), .A2(n582), .ZN(n489) );
  XNOR2_X1 U587 ( .A(n489), .B(n488), .ZN(n593) );
  XNOR2_X1 U588 ( .A(n490), .B(KEYINPUT14), .ZN(n493) );
  NAND2_X1 U589 ( .A1(G952), .A2(n493), .ZN(n491) );
  XNOR2_X1 U590 ( .A(KEYINPUT94), .B(n491), .ZN(n748) );
  NOR2_X1 U591 ( .A1(n748), .A2(G953), .ZN(n492) );
  XNOR2_X1 U592 ( .A(n492), .B(KEYINPUT95), .ZN(n572) );
  NAND2_X1 U593 ( .A1(G902), .A2(n493), .ZN(n569) );
  INV_X1 U594 ( .A(G898), .ZN(n494) );
  NAND2_X1 U595 ( .A1(n494), .A2(G953), .ZN(n760) );
  OR2_X1 U596 ( .A1(n569), .A2(n760), .ZN(n495) );
  NAND2_X1 U597 ( .A1(n572), .A2(n495), .ZN(n496) );
  NAND2_X1 U598 ( .A1(n593), .A2(n496), .ZN(n497) );
  XOR2_X1 U599 ( .A(KEYINPUT12), .B(G140), .Z(n499) );
  XNOR2_X1 U600 ( .A(G143), .B(G122), .ZN(n498) );
  XNOR2_X1 U601 ( .A(n499), .B(n498), .ZN(n506) );
  INV_X1 U602 ( .A(n502), .ZN(n501) );
  INV_X1 U603 ( .A(KEYINPUT11), .ZN(n500) );
  NAND2_X1 U604 ( .A1(n501), .A2(n500), .ZN(n504) );
  NAND2_X1 U605 ( .A1(n502), .A2(KEYINPUT11), .ZN(n503) );
  NAND2_X1 U606 ( .A1(n504), .A2(n503), .ZN(n505) );
  AND2_X1 U607 ( .A1(n507), .A2(G214), .ZN(n510) );
  XNOR2_X1 U608 ( .A(G113), .B(G131), .ZN(n508) );
  XNOR2_X1 U609 ( .A(G104), .B(n508), .ZN(n509) );
  XNOR2_X1 U610 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U611 ( .A(n512), .B(n511), .ZN(n639) );
  NAND2_X1 U612 ( .A1(n639), .A2(n524), .ZN(n514) );
  XOR2_X1 U613 ( .A(KEYINPUT13), .B(G475), .Z(n513) );
  XOR2_X1 U614 ( .A(G122), .B(G107), .Z(n516) );
  XNOR2_X1 U615 ( .A(G116), .B(G134), .ZN(n515) );
  XNOR2_X1 U616 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U617 ( .A(n517), .B(KEYINPUT7), .Z(n520) );
  NAND2_X1 U618 ( .A1(n518), .A2(G217), .ZN(n519) );
  XNOR2_X1 U619 ( .A(n520), .B(n519), .ZN(n523) );
  XNOR2_X1 U620 ( .A(n521), .B(KEYINPUT9), .ZN(n522) );
  XNOR2_X1 U621 ( .A(n523), .B(n522), .ZN(n678) );
  NAND2_X1 U622 ( .A1(n678), .A2(n524), .ZN(n525) );
  XNOR2_X1 U623 ( .A(n525), .B(G478), .ZN(n554) );
  NAND2_X1 U624 ( .A1(n556), .A2(n554), .ZN(n604) );
  INV_X1 U625 ( .A(n604), .ZN(n526) );
  NAND2_X1 U626 ( .A1(n527), .A2(n526), .ZN(n528) );
  OR2_X1 U627 ( .A1(n556), .A2(n554), .ZN(n736) );
  INV_X1 U628 ( .A(n530), .ZN(n531) );
  NOR2_X1 U629 ( .A1(n736), .A2(n531), .ZN(n532) );
  NAND2_X1 U630 ( .A1(n375), .A2(n532), .ZN(n533) );
  INV_X1 U631 ( .A(KEYINPUT104), .ZN(n535) );
  XNOR2_X1 U632 ( .A(n588), .B(n535), .ZN(n719) );
  INV_X1 U633 ( .A(n719), .ZN(n559) );
  NOR2_X1 U634 ( .A1(n534), .A2(n559), .ZN(n536) );
  INV_X1 U635 ( .A(n588), .ZN(n537) );
  AND2_X1 U636 ( .A1(n723), .A2(n537), .ZN(n538) );
  XNOR2_X1 U637 ( .A(n544), .B(n540), .ZN(n541) );
  NAND2_X1 U638 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U639 ( .A1(n544), .A2(KEYINPUT44), .ZN(n545) );
  NAND2_X1 U640 ( .A1(n546), .A2(KEYINPUT44), .ZN(n547) );
  XNOR2_X1 U641 ( .A(n547), .B(KEYINPUT87), .ZN(n566) );
  NOR2_X1 U642 ( .A1(n723), .A2(n713), .ZN(n548) );
  NAND2_X1 U643 ( .A1(n363), .A2(n548), .ZN(n727) );
  INV_X1 U644 ( .A(n605), .ZN(n550) );
  NOR2_X1 U645 ( .A1(n550), .A2(n713), .ZN(n551) );
  NAND2_X1 U646 ( .A1(n551), .A2(n723), .ZN(n552) );
  NOR2_X1 U647 ( .A1(n529), .A2(n552), .ZN(n553) );
  XNOR2_X1 U648 ( .A(n553), .B(KEYINPUT99), .ZN(n689) );
  NAND2_X1 U649 ( .A1(n698), .A2(n689), .ZN(n557) );
  INV_X1 U650 ( .A(n554), .ZN(n555) );
  OR2_X1 U651 ( .A1(n556), .A2(n555), .ZN(n697) );
  NAND2_X1 U652 ( .A1(n556), .A2(n555), .ZN(n617) );
  NAND2_X1 U653 ( .A1(n697), .A2(n617), .ZN(n599) );
  NAND2_X1 U654 ( .A1(n557), .A2(n599), .ZN(n558) );
  XNOR2_X1 U655 ( .A(n558), .B(KEYINPUT102), .ZN(n564) );
  INV_X1 U656 ( .A(n615), .ZN(n561) );
  NAND2_X1 U657 ( .A1(n534), .A2(n559), .ZN(n560) );
  NOR2_X1 U658 ( .A1(n561), .A2(n560), .ZN(n562) );
  NAND2_X1 U659 ( .A1(n563), .A2(n562), .ZN(n656) );
  NAND2_X1 U660 ( .A1(n564), .A2(n656), .ZN(n565) );
  XOR2_X1 U661 ( .A(KEYINPUT83), .B(KEYINPUT45), .Z(n567) );
  NOR2_X1 U662 ( .A1(G900), .A2(n569), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n570), .A2(G953), .ZN(n571) );
  NAND2_X1 U664 ( .A1(n572), .A2(n571), .ZN(n586) );
  INV_X1 U665 ( .A(n608), .ZN(n577) );
  INV_X1 U666 ( .A(KEYINPUT38), .ZN(n575) );
  AND2_X1 U667 ( .A1(n605), .A2(n734), .ZN(n576) );
  INV_X1 U668 ( .A(n617), .ZN(n578) );
  NAND2_X1 U669 ( .A1(n367), .A2(n578), .ZN(n581) );
  XNOR2_X1 U670 ( .A(KEYINPUT110), .B(KEYINPUT40), .ZN(n579) );
  XNOR2_X1 U671 ( .A(n579), .B(KEYINPUT109), .ZN(n580) );
  XNOR2_X1 U672 ( .A(n581), .B(n580), .ZN(n657) );
  INV_X1 U673 ( .A(n582), .ZN(n733) );
  NAND2_X1 U674 ( .A1(n734), .A2(n733), .ZN(n737) );
  XNOR2_X1 U675 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n583) );
  XNOR2_X1 U676 ( .A(n584), .B(n583), .ZN(n732) );
  INV_X1 U677 ( .A(n720), .ZN(n585) );
  NAND2_X1 U678 ( .A1(n586), .A2(n585), .ZN(n587) );
  INV_X1 U679 ( .A(KEYINPUT108), .ZN(n589) );
  NAND2_X1 U680 ( .A1(n732), .A2(n595), .ZN(n592) );
  INV_X1 U681 ( .A(KEYINPUT42), .ZN(n591) );
  XNOR2_X1 U682 ( .A(n592), .B(n591), .ZN(n775) );
  BUF_X1 U683 ( .A(n593), .Z(n594) );
  INV_X1 U684 ( .A(n599), .ZN(n738) );
  INV_X1 U685 ( .A(KEYINPUT79), .ZN(n596) );
  AND2_X1 U686 ( .A1(KEYINPUT79), .A2(KEYINPUT47), .ZN(n598) );
  AND2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U688 ( .A1(n597), .A2(n600), .ZN(n601) );
  NAND2_X1 U689 ( .A1(n602), .A2(n601), .ZN(n610) );
  NOR2_X1 U690 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U691 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U692 ( .A1(n608), .A2(n607), .ZN(n693) );
  INV_X1 U693 ( .A(n693), .ZN(n609) );
  INV_X1 U694 ( .A(KEYINPUT74), .ZN(n611) );
  INV_X1 U695 ( .A(n612), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n613), .A2(n733), .ZN(n614) );
  OR2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n618) );
  INV_X1 U698 ( .A(KEYINPUT105), .ZN(n616) );
  XNOR2_X1 U699 ( .A(n617), .B(n616), .ZN(n694) );
  NAND2_X1 U700 ( .A1(n624), .A2(n627), .ZN(n620) );
  XNOR2_X1 U701 ( .A(KEYINPUT112), .B(KEYINPUT36), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U703 ( .A(n661), .B(KEYINPUT84), .ZN(n622) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT48), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n624), .A2(n534), .ZN(n626) );
  XOR2_X1 U706 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n625) );
  XNOR2_X1 U707 ( .A(n626), .B(n625), .ZN(n628) );
  OR2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n629), .B(KEYINPUT107), .ZN(n774) );
  INV_X1 U710 ( .A(n697), .ZN(n630) );
  AND2_X1 U711 ( .A1(n367), .A2(n630), .ZN(n655) );
  NOR2_X1 U712 ( .A1(n774), .A2(n655), .ZN(n631) );
  AND2_X1 U713 ( .A1(n633), .A2(KEYINPUT2), .ZN(n634) );
  NAND2_X1 U714 ( .A1(n671), .A2(G475), .ZN(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT90), .B(KEYINPUT124), .ZN(n637) );
  XNOR2_X1 U716 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n636) );
  XNOR2_X1 U717 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U718 ( .A(n641), .B(n640), .ZN(n643) );
  INV_X1 U719 ( .A(G952), .ZN(n642) );
  NAND2_X1 U720 ( .A1(n671), .A2(G210), .ZN(n648) );
  XOR2_X1 U721 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n645) );
  XNOR2_X1 U722 ( .A(n648), .B(n647), .ZN(n649) );
  NOR2_X1 U723 ( .A1(n597), .A2(n697), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n651) );
  XNOR2_X1 U725 ( .A(G128), .B(KEYINPUT29), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U727 ( .A(n653), .B(n652), .ZN(G30) );
  NOR2_X1 U728 ( .A1(n597), .A2(n694), .ZN(n654) );
  XOR2_X1 U729 ( .A(G146), .B(n654), .Z(G48) );
  XOR2_X1 U730 ( .A(G134), .B(n655), .Z(G36) );
  XNOR2_X1 U731 ( .A(n656), .B(G101), .ZN(G3) );
  XOR2_X1 U732 ( .A(n657), .B(G131), .Z(G33) );
  XNOR2_X1 U733 ( .A(n658), .B(G110), .ZN(G12) );
  XOR2_X1 U734 ( .A(KEYINPUT117), .B(KEYINPUT37), .Z(n659) );
  XOR2_X1 U735 ( .A(n659), .B(G125), .Z(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(G27) );
  XNOR2_X1 U737 ( .A(n662), .B(G119), .ZN(G21) );
  XOR2_X1 U738 ( .A(n663), .B(G122), .Z(G24) );
  NAND2_X1 U739 ( .A1(n671), .A2(G472), .ZN(n667) );
  BUF_X1 U740 ( .A(n664), .Z(n665) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U742 ( .A1(n668), .A2(n675), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n669) );
  XNOR2_X1 U744 ( .A(n670), .B(n669), .ZN(G57) );
  NAND2_X1 U745 ( .A1(n680), .A2(G217), .ZN(n674) );
  INV_X1 U746 ( .A(n672), .ZN(n673) );
  INV_X1 U747 ( .A(n675), .ZN(n685) );
  NOR2_X1 U748 ( .A1(n676), .A2(n685), .ZN(G66) );
  NAND2_X1 U749 ( .A1(n680), .A2(G478), .ZN(n677) );
  NOR2_X1 U750 ( .A1(n679), .A2(n685), .ZN(G63) );
  NAND2_X1 U751 ( .A1(n680), .A2(G469), .ZN(n684) );
  XNOR2_X1 U752 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n681) );
  XNOR2_X1 U753 ( .A(n681), .B(KEYINPUT58), .ZN(n682) );
  XNOR2_X1 U754 ( .A(n684), .B(n683), .ZN(n686) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(G54) );
  NOR2_X1 U756 ( .A1(n694), .A2(n689), .ZN(n688) );
  XNOR2_X1 U757 ( .A(G104), .B(KEYINPUT113), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n688), .B(n687), .ZN(G6) );
  NOR2_X1 U759 ( .A1(n697), .A2(n689), .ZN(n691) );
  XNOR2_X1 U760 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n690) );
  XNOR2_X1 U761 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U762 ( .A(G107), .B(n692), .ZN(G9) );
  XOR2_X1 U763 ( .A(G143), .B(n693), .Z(G45) );
  NOR2_X1 U764 ( .A1(n698), .A2(n694), .ZN(n695) );
  XOR2_X1 U765 ( .A(KEYINPUT116), .B(n695), .Z(n696) );
  XNOR2_X1 U766 ( .A(G113), .B(n696), .ZN(G15) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U768 ( .A(G116), .B(n699), .Z(G18) );
  BUF_X1 U769 ( .A(n700), .Z(n701) );
  INV_X1 U770 ( .A(n701), .ZN(n741) );
  NAND2_X1 U771 ( .A1(n732), .A2(n741), .ZN(n702) );
  XOR2_X1 U772 ( .A(n702), .B(KEYINPUT122), .Z(n703) );
  NOR2_X1 U773 ( .A1(n766), .A2(KEYINPUT2), .ZN(n705) );
  NOR2_X1 U774 ( .A1(n705), .A2(KEYINPUT80), .ZN(n708) );
  INV_X1 U775 ( .A(n706), .ZN(n707) );
  INV_X1 U776 ( .A(n766), .ZN(n709) );
  NAND2_X1 U777 ( .A1(n709), .A2(KEYINPUT80), .ZN(n710) );
  INV_X1 U778 ( .A(KEYINPUT2), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n534), .A2(n713), .ZN(n714) );
  NAND2_X1 U780 ( .A1(n714), .A2(KEYINPUT50), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n715), .A2(KEYINPUT50), .ZN(n716) );
  NAND2_X1 U782 ( .A1(n534), .A2(n716), .ZN(n717) );
  NAND2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n726) );
  XOR2_X1 U784 ( .A(KEYINPUT118), .B(KEYINPUT49), .Z(n722) );
  NAND2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U786 ( .A(n722), .B(n721), .ZN(n724) );
  AND2_X1 U787 ( .A1(n723), .A2(n724), .ZN(n725) );
  NAND2_X1 U788 ( .A1(n726), .A2(n725), .ZN(n728) );
  AND2_X1 U789 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U790 ( .A(n729), .B(KEYINPUT119), .Z(n730) );
  XNOR2_X1 U791 ( .A(KEYINPUT51), .B(n730), .ZN(n731) );
  NAND2_X1 U792 ( .A1(n732), .A2(n731), .ZN(n744) );
  NOR2_X1 U793 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U794 ( .A1(n736), .A2(n735), .ZN(n740) );
  NOR2_X1 U795 ( .A1(n738), .A2(n737), .ZN(n739) );
  OR2_X1 U796 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U797 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U798 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U799 ( .A(n745), .B(KEYINPUT120), .Z(n746) );
  XNOR2_X1 U800 ( .A(KEYINPUT52), .B(n746), .ZN(n747) );
  NOR2_X1 U801 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U802 ( .A(KEYINPUT121), .B(n749), .Z(n750) );
  XNOR2_X1 U803 ( .A(KEYINPUT53), .B(n751), .ZN(G75) );
  NOR2_X1 U804 ( .A1(n752), .A2(G953), .ZN(n758) );
  XOR2_X1 U805 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n754) );
  NAND2_X1 U806 ( .A1(G224), .A2(G953), .ZN(n753) );
  XNOR2_X1 U807 ( .A(n754), .B(n753), .ZN(n755) );
  NAND2_X1 U808 ( .A1(G898), .A2(n755), .ZN(n756) );
  XOR2_X1 U809 ( .A(KEYINPUT126), .B(n756), .Z(n757) );
  NOR2_X1 U810 ( .A1(n758), .A2(n757), .ZN(n763) );
  XNOR2_X1 U811 ( .A(n759), .B(G101), .ZN(n761) );
  AND2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U813 ( .A(n763), .B(n762), .Z(G69) );
  XOR2_X1 U814 ( .A(n764), .B(n765), .Z(n769) );
  XNOR2_X1 U815 ( .A(n766), .B(n769), .ZN(n767) );
  NOR2_X1 U816 ( .A1(n767), .A2(G953), .ZN(n768) );
  XNOR2_X1 U817 ( .A(KEYINPUT127), .B(n768), .ZN(n773) );
  XNOR2_X1 U818 ( .A(n769), .B(G227), .ZN(n770) );
  NAND2_X1 U819 ( .A1(n770), .A2(G900), .ZN(n771) );
  NAND2_X1 U820 ( .A1(n771), .A2(G953), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n773), .A2(n772), .ZN(G72) );
  XOR2_X1 U822 ( .A(G140), .B(n774), .Z(G42) );
  XOR2_X1 U823 ( .A(n775), .B(G137), .Z(G39) );
endmodule

