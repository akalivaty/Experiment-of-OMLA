

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761;

  XNOR2_X1 U369 ( .A(n508), .B(n401), .ZN(n410) );
  NOR2_X1 U370 ( .A1(G953), .A2(G237), .ZN(n510) );
  XNOR2_X1 U371 ( .A(n425), .B(n346), .ZN(n375) );
  NAND2_X1 U372 ( .A1(n375), .A2(n372), .ZN(n374) );
  INV_X2 U373 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U374 ( .A(n363), .B(n553), .ZN(n681) );
  XNOR2_X1 U375 ( .A(n434), .B(KEYINPUT35), .ZN(n682) );
  NOR2_X2 U376 ( .A1(n606), .A2(n387), .ZN(n726) );
  XNOR2_X2 U377 ( .A(n384), .B(KEYINPUT33), .ZN(n675) );
  AND2_X1 U378 ( .A1(n357), .A2(n353), .ZN(n352) );
  NAND2_X1 U379 ( .A1(n352), .A2(n350), .ZN(n635) );
  NAND2_X1 U380 ( .A1(n351), .A2(n355), .ZN(n350) );
  NAND2_X1 U381 ( .A1(n446), .A2(n445), .ZN(n631) );
  INV_X1 U382 ( .A(KEYINPUT84), .ZN(n377) );
  INV_X1 U383 ( .A(KEYINPUT87), .ZN(n355) );
  INV_X1 U384 ( .A(KEYINPUT44), .ZN(n372) );
  NOR2_X1 U385 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U386 ( .A1(n349), .A2(n745), .ZN(n348) );
  XNOR2_X1 U387 ( .A(n742), .B(KEYINPUT123), .ZN(n349) );
  AND2_X1 U388 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U389 ( .A1(n637), .A2(KEYINPUT2), .ZN(n638) );
  XNOR2_X1 U390 ( .A(n366), .B(n572), .ZN(n365) );
  NAND2_X1 U391 ( .A1(n368), .A2(n367), .ZN(n366) );
  AND2_X1 U392 ( .A1(n635), .A2(n571), .ZN(n368) );
  NAND2_X1 U393 ( .A1(n373), .A2(n372), .ZN(n371) );
  XNOR2_X1 U394 ( .A(n431), .B(n430), .ZN(n429) );
  NAND2_X1 U395 ( .A1(n364), .A2(n398), .ZN(n363) );
  NAND2_X1 U396 ( .A1(n410), .A2(n358), .ZN(n357) );
  XNOR2_X1 U397 ( .A(n508), .B(n401), .ZN(n364) );
  XNOR2_X1 U398 ( .A(n585), .B(KEYINPUT40), .ZN(n760) );
  AND2_X1 U399 ( .A1(n624), .A2(n725), .ZN(n585) );
  AND2_X1 U400 ( .A1(n354), .A2(n657), .ZN(n353) );
  XNOR2_X1 U401 ( .A(n383), .B(n382), .ZN(n561) );
  NAND2_X1 U402 ( .A1(n356), .A2(n355), .ZN(n354) );
  AND2_X1 U403 ( .A1(n578), .A2(n443), .ZN(n611) );
  INV_X1 U404 ( .A(n663), .ZN(n385) );
  INV_X1 U405 ( .A(n396), .ZN(n356) );
  OR2_X2 U406 ( .A1(n564), .A2(n598), .ZN(n384) );
  XNOR2_X1 U407 ( .A(n584), .B(KEYINPUT38), .ZN(n642) );
  NAND2_X1 U408 ( .A1(n392), .A2(n643), .ZN(n440) );
  NAND2_X1 U409 ( .A1(n631), .A2(n542), .ZN(n519) );
  NOR2_X2 U410 ( .A1(n698), .A2(G902), .ZN(n529) );
  XNOR2_X1 U411 ( .A(n518), .B(n462), .ZN(n739) );
  XNOR2_X1 U412 ( .A(n394), .B(n509), .ZN(n749) );
  INV_X1 U413 ( .A(n615), .ZN(n381) );
  NOR2_X1 U414 ( .A1(n625), .A2(n439), .ZN(n403) );
  XNOR2_X1 U415 ( .A(KEYINPUT48), .B(KEYINPUT86), .ZN(n615) );
  XNOR2_X1 U416 ( .A(G119), .B(G116), .ZN(n416) );
  INV_X1 U417 ( .A(KEYINPUT89), .ZN(n346) );
  XOR2_X1 U418 ( .A(KEYINPUT68), .B(G101), .Z(n514) );
  NAND2_X1 U419 ( .A1(n345), .A2(n371), .ZN(n370) );
  INV_X1 U420 ( .A(n375), .ZN(n345) );
  XNOR2_X1 U421 ( .A(n348), .B(n347), .ZN(G69) );
  XNOR2_X1 U422 ( .A(n746), .B(KEYINPUT124), .ZN(n347) );
  INV_X1 U423 ( .A(n410), .ZN(n351) );
  AND2_X1 U424 ( .A1(n396), .A2(KEYINPUT87), .ZN(n358) );
  NAND2_X1 U425 ( .A1(n359), .A2(n404), .ZN(n414) );
  NAND2_X1 U426 ( .A1(n360), .A2(n417), .ZN(n359) );
  AND2_X1 U427 ( .A1(n376), .A2(n400), .ZN(n361) );
  NAND2_X1 U428 ( .A1(n628), .A2(n439), .ZN(n362) );
  NAND2_X1 U429 ( .A1(n681), .A2(n634), .ZN(n425) );
  NAND2_X2 U430 ( .A1(n369), .A2(n365), .ZN(n574) );
  NAND2_X1 U431 ( .A1(n682), .A2(KEYINPUT44), .ZN(n367) );
  NAND2_X1 U432 ( .A1(n374), .A2(n370), .ZN(n369) );
  INV_X1 U433 ( .A(n682), .ZN(n373) );
  AND2_X1 U434 ( .A1(n376), .A2(n736), .ZN(n395) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n376) );
  NAND2_X1 U436 ( .A1(n637), .A2(n403), .ZN(n417) );
  AND2_X1 U437 ( .A1(n637), .A2(n755), .ZN(n742) );
  AND2_X1 U438 ( .A1(n637), .A2(KEYINPUT2), .ZN(n426) );
  XNOR2_X2 U439 ( .A(n574), .B(KEYINPUT45), .ZN(n637) );
  XNOR2_X2 U440 ( .A(n525), .B(n524), .ZN(n698) );
  XNOR2_X2 U441 ( .A(n749), .B(G146), .ZN(n525) );
  NAND2_X1 U442 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U443 ( .A(n636), .ZN(n379) );
  XNOR2_X1 U444 ( .A(n616), .B(n381), .ZN(n380) );
  NAND2_X1 U445 ( .A1(n675), .A2(n561), .ZN(n436) );
  XNOR2_X1 U446 ( .A(n409), .B(KEYINPUT93), .ZN(n382) );
  NOR2_X1 U447 ( .A1(n605), .A2(n472), .ZN(n383) );
  NAND2_X1 U448 ( .A1(n556), .A2(n555), .ZN(n564) );
  NAND2_X1 U449 ( .A1(n506), .A2(n385), .ZN(n566) );
  XNOR2_X2 U450 ( .A(n386), .B(KEYINPUT0), .ZN(n506) );
  NOR2_X2 U451 ( .A1(n605), .A2(n472), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n436), .B(n557), .ZN(n435) );
  NAND2_X1 U453 ( .A1(n435), .A2(n560), .ZN(n434) );
  BUF_X1 U454 ( .A(n605), .Z(n387) );
  NAND2_X1 U455 ( .A1(n441), .A2(n419), .ZN(n390) );
  NAND2_X1 U456 ( .A1(n388), .A2(n389), .ZN(n391) );
  NAND2_X1 U457 ( .A1(n391), .A2(n390), .ZN(n418) );
  INV_X1 U458 ( .A(n441), .ZN(n388) );
  INV_X1 U459 ( .A(n419), .ZN(n389) );
  XNOR2_X2 U460 ( .A(n433), .B(n596), .ZN(n674) );
  INV_X1 U461 ( .A(n392), .ZN(n584) );
  XNOR2_X2 U462 ( .A(n406), .B(n393), .ZN(n392) );
  AND2_X1 U463 ( .A1(n464), .A2(G210), .ZN(n393) );
  XNOR2_X1 U464 ( .A(n481), .B(KEYINPUT4), .ZN(n394) );
  XNOR2_X1 U465 ( .A(n481), .B(KEYINPUT4), .ZN(n441) );
  NOR2_X2 U466 ( .A1(n694), .A2(n709), .ZN(n696) );
  NOR2_X2 U467 ( .A1(n710), .A2(n709), .ZN(n712) );
  XNOR2_X1 U468 ( .A(n416), .B(KEYINPUT3), .ZN(n415) );
  INV_X1 U469 ( .A(KEYINPUT46), .ZN(n430) );
  OR2_X1 U470 ( .A1(n516), .A2(n518), .ZN(n452) );
  XOR2_X1 U471 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n474) );
  XNOR2_X1 U472 ( .A(G122), .B(KEYINPUT99), .ZN(n473) );
  XOR2_X1 U473 ( .A(G131), .B(G134), .Z(n509) );
  XNOR2_X1 U474 ( .A(G137), .B(G140), .ZN(n532) );
  NAND2_X1 U475 ( .A1(n464), .A2(G214), .ZN(n643) );
  XNOR2_X1 U476 ( .A(KEYINPUT16), .B(G122), .ZN(n461) );
  XNOR2_X1 U477 ( .A(n413), .B(KEYINPUT39), .ZN(n624) );
  XOR2_X1 U478 ( .A(G137), .B(KEYINPUT5), .Z(n512) );
  INV_X1 U479 ( .A(KEYINPUT73), .ZN(n459) );
  NAND2_X1 U480 ( .A1(n625), .A2(n439), .ZN(n438) );
  INV_X1 U481 ( .A(KEYINPUT83), .ZN(n439) );
  AND2_X1 U482 ( .A1(n614), .A2(n733), .ZN(n432) );
  INV_X1 U483 ( .A(G237), .ZN(n463) );
  XNOR2_X1 U484 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  XOR2_X1 U485 ( .A(G122), .B(G104), .Z(n489) );
  XNOR2_X1 U486 ( .A(G113), .B(G143), .ZN(n488) );
  XNOR2_X1 U487 ( .A(G131), .B(G140), .ZN(n490) );
  NAND2_X1 U488 ( .A1(G234), .A2(G237), .ZN(n466) );
  INV_X1 U489 ( .A(G902), .ZN(n542) );
  NAND2_X1 U490 ( .A1(n452), .A2(n451), .ZN(n450) );
  XNOR2_X1 U491 ( .A(G119), .B(G128), .ZN(n537) );
  INV_X1 U492 ( .A(KEYINPUT10), .ZN(n494) );
  XOR2_X1 U493 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n480) );
  XNOR2_X1 U494 ( .A(G116), .B(G107), .ZN(n476) );
  NAND2_X1 U495 ( .A1(n395), .A2(n426), .ZN(n437) );
  INV_X1 U496 ( .A(KEYINPUT34), .ZN(n557) );
  INV_X1 U497 ( .A(KEYINPUT0), .ZN(n409) );
  XNOR2_X1 U498 ( .A(n576), .B(n575), .ZN(n578) );
  INV_X1 U499 ( .A(n587), .ZN(n444) );
  XNOR2_X1 U500 ( .A(n691), .B(KEYINPUT59), .ZN(n692) );
  XNOR2_X1 U501 ( .A(n520), .B(KEYINPUT95), .ZN(n521) );
  XNOR2_X1 U502 ( .A(n704), .B(n706), .ZN(n707) );
  NOR2_X1 U503 ( .A1(n755), .A2(G952), .ZN(n709) );
  XNOR2_X1 U504 ( .A(n415), .B(n460), .ZN(n517) );
  AND2_X1 U505 ( .A1(n531), .A2(n598), .ZN(n396) );
  AND2_X1 U506 ( .A1(n680), .A2(n679), .ZN(n397) );
  NOR2_X1 U507 ( .A1(n550), .A2(n549), .ZN(n398) );
  NOR2_X1 U508 ( .A1(n619), .A2(n554), .ZN(n399) );
  AND2_X1 U509 ( .A1(n736), .A2(n438), .ZN(n400) );
  XOR2_X1 U510 ( .A(n507), .B(KEYINPUT22), .Z(n401) );
  XOR2_X1 U511 ( .A(n631), .B(n630), .Z(n402) );
  XNOR2_X1 U512 ( .A(KEYINPUT66), .B(n627), .ZN(n404) );
  XNOR2_X1 U513 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n405) );
  NAND2_X1 U514 ( .A1(n703), .A2(n625), .ZN(n406) );
  XNOR2_X1 U515 ( .A(n407), .B(n739), .ZN(n703) );
  XNOR2_X1 U516 ( .A(n418), .B(n522), .ZN(n407) );
  BUF_X1 U517 ( .A(n761), .Z(n408) );
  XNOR2_X1 U518 ( .A(n574), .B(n573), .ZN(n628) );
  BUF_X1 U519 ( .A(n681), .Z(n411) );
  BUF_X2 U520 ( .A(n702), .Z(n412) );
  AND2_X2 U521 ( .A1(n414), .A2(n437), .ZN(n702) );
  NAND2_X1 U522 ( .A1(n611), .A2(n642), .ZN(n413) );
  XNOR2_X2 U523 ( .A(n547), .B(n546), .ZN(n657) );
  AND2_X1 U524 ( .A1(n577), .A2(n444), .ZN(n443) );
  XNOR2_X1 U525 ( .A(n495), .B(KEYINPUT77), .ZN(n420) );
  XNOR2_X2 U526 ( .A(G146), .B(G125), .ZN(n495) );
  XNOR2_X1 U527 ( .A(n456), .B(n455), .ZN(n421) );
  XNOR2_X1 U528 ( .A(n421), .B(n420), .ZN(n419) );
  XNOR2_X2 U529 ( .A(n442), .B(n454), .ZN(n481) );
  XNOR2_X1 U530 ( .A(n422), .B(n405), .ZN(G75) );
  NAND2_X1 U531 ( .A1(n423), .A2(n397), .ZN(n422) );
  NAND2_X1 U532 ( .A1(n424), .A2(n437), .ZN(n423) );
  XNOR2_X1 U533 ( .A(n641), .B(KEYINPUT80), .ZN(n424) );
  XNOR2_X1 U534 ( .A(n427), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U535 ( .A1(n428), .A2(n633), .ZN(n427) );
  XNOR2_X1 U536 ( .A(n632), .B(n402), .ZN(n428) );
  NAND2_X1 U537 ( .A1(n432), .A2(n429), .ZN(n616) );
  OR2_X2 U538 ( .A1(n761), .A2(n760), .ZN(n431) );
  NOR2_X1 U539 ( .A1(n674), .A2(n606), .ZN(n597) );
  NAND2_X1 U540 ( .A1(n649), .A2(n646), .ZN(n433) );
  XNOR2_X2 U541 ( .A(n595), .B(KEYINPUT109), .ZN(n649) );
  NAND2_X2 U542 ( .A1(n506), .A2(n505), .ZN(n508) );
  XNOR2_X2 U543 ( .A(n602), .B(KEYINPUT19), .ZN(n605) );
  XNOR2_X2 U544 ( .A(n440), .B(n465), .ZN(n602) );
  NAND2_X1 U545 ( .A1(n410), .A2(n399), .ZN(n634) );
  XNOR2_X2 U546 ( .A(G128), .B(KEYINPUT64), .ZN(n442) );
  NAND2_X1 U547 ( .A1(n447), .A2(n525), .ZN(n445) );
  NAND2_X1 U548 ( .A1(n453), .A2(n450), .ZN(n446) );
  INV_X1 U549 ( .A(n525), .ZN(n453) );
  NAND2_X1 U550 ( .A1(n449), .A2(n448), .ZN(n447) );
  NAND2_X1 U551 ( .A1(n516), .A2(n517), .ZN(n448) );
  OR2_X1 U552 ( .A1(n516), .A2(n517), .ZN(n449) );
  NAND2_X1 U553 ( .A1(n518), .A2(n516), .ZN(n451) );
  XNOR2_X2 U554 ( .A(n519), .B(G472), .ZN(n660) );
  XNOR2_X1 U555 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U556 ( .A(n527), .B(n526), .ZN(n528) );
  INV_X1 U557 ( .A(KEYINPUT30), .ZN(n575) );
  XNOR2_X1 U558 ( .A(n748), .B(n521), .ZN(n523) );
  INV_X1 U559 ( .A(G143), .ZN(n454) );
  XNOR2_X1 U560 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n455) );
  NAND2_X1 U561 ( .A1(n755), .A2(G224), .ZN(n456) );
  XNOR2_X1 U562 ( .A(n514), .B(KEYINPUT74), .ZN(n458) );
  XOR2_X1 U563 ( .A(G104), .B(G110), .Z(n457) );
  XNOR2_X1 U564 ( .A(n457), .B(G107), .ZN(n737) );
  XNOR2_X1 U565 ( .A(n458), .B(n737), .ZN(n522) );
  XNOR2_X1 U566 ( .A(n459), .B(G113), .ZN(n460) );
  INV_X1 U567 ( .A(n517), .ZN(n518) );
  XNOR2_X1 U568 ( .A(n461), .B(KEYINPUT76), .ZN(n462) );
  NAND2_X1 U569 ( .A1(n542), .A2(n463), .ZN(n464) );
  INV_X1 U570 ( .A(KEYINPUT90), .ZN(n465) );
  XNOR2_X1 U571 ( .A(n466), .B(KEYINPUT14), .ZN(n467) );
  AND2_X1 U572 ( .A1(n467), .A2(G952), .ZN(n672) );
  AND2_X1 U573 ( .A1(n672), .A2(n755), .ZN(n583) );
  NAND2_X1 U574 ( .A1(G902), .A2(n467), .ZN(n579) );
  INV_X1 U575 ( .A(n579), .ZN(n468) );
  NOR2_X1 U576 ( .A1(G898), .A2(n755), .ZN(n741) );
  NAND2_X1 U577 ( .A1(n468), .A2(n741), .ZN(n470) );
  INV_X1 U578 ( .A(KEYINPUT92), .ZN(n469) );
  XNOR2_X1 U579 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U580 ( .A1(n583), .A2(n471), .ZN(n472) );
  XNOR2_X1 U581 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U582 ( .A(n475), .B(KEYINPUT9), .Z(n477) );
  XNOR2_X1 U583 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U584 ( .A(n478), .B(KEYINPUT7), .Z(n485) );
  NAND2_X1 U585 ( .A1(G234), .A2(n755), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n480), .B(n479), .ZN(n534) );
  AND2_X1 U587 ( .A1(n534), .A2(G217), .ZN(n483) );
  XNOR2_X1 U588 ( .A(n481), .B(G134), .ZN(n482) );
  XNOR2_X1 U589 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U590 ( .A(n485), .B(n484), .ZN(n687) );
  NAND2_X1 U591 ( .A1(n687), .A2(n542), .ZN(n487) );
  INV_X1 U592 ( .A(G478), .ZN(n486) );
  XNOR2_X1 U593 ( .A(n487), .B(n486), .ZN(n568) );
  XNOR2_X1 U594 ( .A(n489), .B(n488), .ZN(n493) );
  XOR2_X1 U595 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n491) );
  XNOR2_X1 U596 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U597 ( .A(n493), .B(n492), .Z(n498) );
  XNOR2_X1 U598 ( .A(n495), .B(n494), .ZN(n747) );
  NAND2_X1 U599 ( .A1(G214), .A2(n510), .ZN(n496) );
  XNOR2_X1 U600 ( .A(n747), .B(n496), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n498), .B(n497), .ZN(n691) );
  NAND2_X1 U602 ( .A1(n691), .A2(n542), .ZN(n500) );
  XNOR2_X1 U603 ( .A(KEYINPUT13), .B(G475), .ZN(n499) );
  XNOR2_X1 U604 ( .A(n500), .B(n499), .ZN(n558) );
  AND2_X1 U605 ( .A1(n568), .A2(n558), .ZN(n646) );
  XOR2_X1 U606 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n503) );
  NAND2_X1 U607 ( .A1(n625), .A2(G234), .ZN(n501) );
  XNOR2_X1 U608 ( .A(n501), .B(KEYINPUT20), .ZN(n543) );
  NAND2_X1 U609 ( .A1(n543), .A2(G221), .ZN(n502) );
  XNOR2_X1 U610 ( .A(n503), .B(n502), .ZN(n656) );
  NAND2_X1 U611 ( .A1(n646), .A2(n656), .ZN(n504) );
  XNOR2_X1 U612 ( .A(n504), .B(KEYINPUT103), .ZN(n505) );
  INV_X1 U613 ( .A(KEYINPUT75), .ZN(n507) );
  NAND2_X1 U614 ( .A1(n510), .A2(G210), .ZN(n511) );
  XNOR2_X1 U615 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U616 ( .A(n513), .B(KEYINPUT98), .Z(n515) );
  XNOR2_X1 U617 ( .A(n660), .B(KEYINPUT6), .ZN(n598) );
  XNOR2_X1 U618 ( .A(n598), .B(KEYINPUT79), .ZN(n550) );
  XNOR2_X1 U619 ( .A(KEYINPUT94), .B(n532), .ZN(n748) );
  NAND2_X1 U620 ( .A1(G227), .A2(n755), .ZN(n520) );
  XNOR2_X1 U621 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U622 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n527) );
  INV_X1 U623 ( .A(G469), .ZN(n526) );
  XNOR2_X2 U624 ( .A(n529), .B(n528), .ZN(n592) );
  INV_X1 U625 ( .A(KEYINPUT1), .ZN(n530) );
  XNOR2_X1 U626 ( .A(n592), .B(n530), .ZN(n556) );
  INV_X1 U627 ( .A(n556), .ZN(n531) );
  INV_X1 U628 ( .A(n531), .ZN(n619) );
  INV_X1 U629 ( .A(n532), .ZN(n533) );
  XOR2_X1 U630 ( .A(n533), .B(KEYINPUT24), .Z(n536) );
  NAND2_X1 U631 ( .A1(G221), .A2(n534), .ZN(n535) );
  XNOR2_X1 U632 ( .A(n536), .B(n535), .ZN(n541) );
  XOR2_X1 U633 ( .A(KEYINPUT23), .B(G110), .Z(n538) );
  XNOR2_X1 U634 ( .A(n538), .B(n537), .ZN(n539) );
  XOR2_X1 U635 ( .A(n539), .B(n747), .Z(n540) );
  XNOR2_X1 U636 ( .A(n541), .B(n540), .ZN(n684) );
  NAND2_X1 U637 ( .A1(n684), .A2(n542), .ZN(n547) );
  NAND2_X1 U638 ( .A1(G217), .A2(n543), .ZN(n545) );
  INV_X1 U639 ( .A(KEYINPUT25), .ZN(n544) );
  XNOR2_X1 U640 ( .A(n545), .B(n544), .ZN(n546) );
  INV_X1 U641 ( .A(n657), .ZN(n548) );
  NAND2_X1 U642 ( .A1(n619), .A2(n548), .ZN(n549) );
  XNOR2_X1 U643 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n552) );
  INV_X1 U644 ( .A(KEYINPUT65), .ZN(n551) );
  XNOR2_X1 U645 ( .A(n552), .B(n551), .ZN(n553) );
  OR2_X1 U646 ( .A1(n660), .A2(n657), .ZN(n554) );
  NAND2_X1 U647 ( .A1(n656), .A2(n657), .ZN(n654) );
  INV_X1 U648 ( .A(n654), .ZN(n555) );
  INV_X1 U649 ( .A(n568), .ZN(n559) );
  INV_X1 U650 ( .A(n558), .ZN(n567) );
  NAND2_X1 U651 ( .A1(n559), .A2(n567), .ZN(n609) );
  INV_X1 U652 ( .A(n609), .ZN(n560) );
  NOR2_X1 U653 ( .A1(n592), .A2(n654), .ZN(n577) );
  NAND2_X1 U654 ( .A1(n561), .A2(n577), .ZN(n562) );
  XNOR2_X1 U655 ( .A(n562), .B(KEYINPUT97), .ZN(n563) );
  INV_X1 U656 ( .A(n660), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n563), .A2(n589), .ZN(n716) );
  OR2_X1 U658 ( .A1(n564), .A2(n589), .ZN(n663) );
  INV_X1 U659 ( .A(KEYINPUT31), .ZN(n565) );
  XNOR2_X1 U660 ( .A(n566), .B(n565), .ZN(n730) );
  NAND2_X1 U661 ( .A1(n716), .A2(n730), .ZN(n570) );
  NOR2_X1 U662 ( .A1(n568), .A2(n567), .ZN(n719) );
  XNOR2_X1 U663 ( .A(KEYINPUT102), .B(n719), .ZN(n623) );
  INV_X1 U664 ( .A(n623), .ZN(n569) );
  NAND2_X1 U665 ( .A1(n568), .A2(n567), .ZN(n728) );
  NAND2_X1 U666 ( .A1(n569), .A2(n728), .ZN(n648) );
  NAND2_X1 U667 ( .A1(n570), .A2(n648), .ZN(n571) );
  INV_X1 U668 ( .A(KEYINPUT88), .ZN(n572) );
  INV_X1 U669 ( .A(KEYINPUT45), .ZN(n573) );
  NAND2_X1 U670 ( .A1(n660), .A2(n643), .ZN(n576) );
  NOR2_X1 U671 ( .A1(G900), .A2(n579), .ZN(n580) );
  NAND2_X1 U672 ( .A1(G953), .A2(n580), .ZN(n581) );
  XOR2_X1 U673 ( .A(KEYINPUT104), .B(n581), .Z(n582) );
  NOR2_X1 U674 ( .A1(n583), .A2(n582), .ZN(n587) );
  INV_X1 U675 ( .A(n728), .ZN(n725) );
  XOR2_X1 U676 ( .A(KEYINPUT107), .B(KEYINPUT28), .Z(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT108), .B(n586), .ZN(n591) );
  NOR2_X1 U678 ( .A1(n587), .A2(n657), .ZN(n588) );
  NAND2_X1 U679 ( .A1(n656), .A2(n588), .ZN(n599) );
  NOR2_X1 U680 ( .A1(n589), .A2(n599), .ZN(n590) );
  XNOR2_X1 U681 ( .A(n591), .B(n590), .ZN(n594) );
  XOR2_X1 U682 ( .A(n592), .B(KEYINPUT106), .Z(n593) );
  NAND2_X1 U683 ( .A1(n594), .A2(n593), .ZN(n606) );
  XOR2_X1 U684 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n596) );
  NAND2_X1 U685 ( .A1(n642), .A2(n643), .ZN(n595) );
  XNOR2_X1 U686 ( .A(n597), .B(KEYINPUT42), .ZN(n761) );
  NOR2_X1 U687 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U688 ( .A(n600), .B(KEYINPUT105), .ZN(n601) );
  NOR2_X1 U689 ( .A1(n728), .A2(n601), .ZN(n617) );
  NAND2_X1 U690 ( .A1(n617), .A2(n602), .ZN(n603) );
  XOR2_X1 U691 ( .A(KEYINPUT36), .B(n603), .Z(n604) );
  NAND2_X1 U692 ( .A1(n604), .A2(n619), .ZN(n733) );
  NAND2_X1 U693 ( .A1(n726), .A2(n648), .ZN(n607) );
  NOR2_X1 U694 ( .A1(n607), .A2(KEYINPUT69), .ZN(n608) );
  XOR2_X1 U695 ( .A(KEYINPUT47), .B(n608), .Z(n613) );
  NOR2_X1 U696 ( .A1(n584), .A2(n609), .ZN(n610) );
  AND2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n723) );
  XOR2_X1 U698 ( .A(KEYINPUT81), .B(n723), .Z(n612) );
  NOR2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n617), .A2(n643), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U702 ( .A(n620), .B(KEYINPUT43), .ZN(n622) );
  INV_X1 U703 ( .A(n584), .ZN(n621) );
  NOR2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n636) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n736) );
  INV_X1 U706 ( .A(n625), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n702), .A2(G472), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT91), .B(KEYINPUT111), .Z(n629) );
  XNOR2_X1 U710 ( .A(n629), .B(KEYINPUT62), .ZN(n630) );
  INV_X1 U711 ( .A(n709), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n634), .B(G110), .ZN(G12) );
  XNOR2_X1 U713 ( .A(n635), .B(G101), .ZN(G3) );
  XOR2_X1 U714 ( .A(G140), .B(n636), .Z(G42) );
  NOR2_X1 U715 ( .A1(n395), .A2(KEYINPUT2), .ZN(n640) );
  XNOR2_X1 U716 ( .A(n638), .B(KEYINPUT82), .ZN(n639) );
  INV_X1 U717 ( .A(n642), .ZN(n645) );
  INV_X1 U718 ( .A(n643), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U721 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U722 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U723 ( .A1(n675), .A2(n652), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT116), .B(n653), .Z(n668) );
  NAND2_X1 U725 ( .A1(n654), .A2(n531), .ZN(n655) );
  XNOR2_X1 U726 ( .A(n655), .B(KEYINPUT50), .ZN(n662) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U728 ( .A(KEYINPUT49), .B(n658), .Z(n659) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n662), .A2(n661), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U732 ( .A(KEYINPUT51), .B(n665), .ZN(n666) );
  NOR2_X1 U733 ( .A1(n674), .A2(n666), .ZN(n667) );
  NOR2_X1 U734 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U735 ( .A(n669), .B(KEYINPUT52), .Z(n671) );
  INV_X1 U736 ( .A(KEYINPUT117), .ZN(n670) );
  XNOR2_X1 U737 ( .A(n671), .B(n670), .ZN(n673) );
  NAND2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n680) );
  INV_X1 U739 ( .A(n674), .ZN(n676) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U741 ( .A(n677), .B(KEYINPUT118), .ZN(n678) );
  AND2_X1 U742 ( .A1(n678), .A2(n755), .ZN(n679) );
  XNOR2_X1 U743 ( .A(n411), .B(G119), .ZN(G21) );
  XOR2_X1 U744 ( .A(n682), .B(G122), .Z(G24) );
  NAND2_X1 U745 ( .A1(n412), .A2(G217), .ZN(n683) );
  XOR2_X1 U746 ( .A(n683), .B(n684), .Z(n685) );
  NOR2_X1 U747 ( .A1(n685), .A2(n709), .ZN(G66) );
  NAND2_X1 U748 ( .A1(n412), .A2(G478), .ZN(n689) );
  XNOR2_X1 U749 ( .A(KEYINPUT121), .B(KEYINPUT122), .ZN(n686) );
  XNOR2_X1 U750 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U751 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U752 ( .A1(n690), .A2(n709), .ZN(G63) );
  NAND2_X1 U753 ( .A1(n702), .A2(G475), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n693), .B(n692), .ZN(n694) );
  XOR2_X1 U755 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n695) );
  XNOR2_X1 U756 ( .A(n696), .B(n695), .ZN(G60) );
  NAND2_X1 U757 ( .A1(n412), .A2(G469), .ZN(n700) );
  XOR2_X1 U758 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n697) );
  XNOR2_X1 U759 ( .A(n698), .B(n697), .ZN(n699) );
  XNOR2_X1 U760 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U761 ( .A1(n701), .A2(n709), .ZN(G54) );
  NAND2_X1 U762 ( .A1(n702), .A2(G210), .ZN(n708) );
  BUF_X1 U763 ( .A(n703), .Z(n704) );
  XNOR2_X1 U764 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n705) );
  XNOR2_X1 U765 ( .A(n705), .B(KEYINPUT55), .ZN(n706) );
  XNOR2_X1 U766 ( .A(n708), .B(n707), .ZN(n710) );
  XOR2_X1 U767 ( .A(KEYINPUT85), .B(KEYINPUT56), .Z(n711) );
  XNOR2_X1 U768 ( .A(n712), .B(n711), .ZN(G51) );
  NOR2_X1 U769 ( .A1(n728), .A2(n716), .ZN(n713) );
  XOR2_X1 U770 ( .A(G104), .B(n713), .Z(G6) );
  XOR2_X1 U771 ( .A(KEYINPUT26), .B(KEYINPUT112), .Z(n715) );
  XNOR2_X1 U772 ( .A(G107), .B(KEYINPUT27), .ZN(n714) );
  XNOR2_X1 U773 ( .A(n715), .B(n714), .ZN(n718) );
  INV_X1 U774 ( .A(n719), .ZN(n731) );
  NOR2_X1 U775 ( .A1(n731), .A2(n716), .ZN(n717) );
  XOR2_X1 U776 ( .A(n718), .B(n717), .Z(G9) );
  XOR2_X1 U777 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n721) );
  NAND2_X1 U778 ( .A1(n726), .A2(n719), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U780 ( .A(G128), .B(n722), .Z(G30) );
  XOR2_X1 U781 ( .A(G143), .B(n723), .Z(n724) );
  XNOR2_X1 U782 ( .A(KEYINPUT114), .B(n724), .ZN(G45) );
  NAND2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U784 ( .A(G146), .B(n727), .ZN(G48) );
  NOR2_X1 U785 ( .A1(n728), .A2(n730), .ZN(n729) );
  XOR2_X1 U786 ( .A(G113), .B(n729), .Z(G15) );
  NOR2_X1 U787 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U788 ( .A(G116), .B(n732), .Z(G18) );
  XNOR2_X1 U789 ( .A(KEYINPUT115), .B(KEYINPUT37), .ZN(n734) );
  XNOR2_X1 U790 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U791 ( .A(G125), .B(n735), .ZN(G27) );
  XNOR2_X1 U792 ( .A(G134), .B(n736), .ZN(G36) );
  XNOR2_X1 U793 ( .A(n737), .B(G101), .ZN(n738) );
  XNOR2_X1 U794 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U795 ( .A1(n741), .A2(n740), .ZN(n746) );
  NAND2_X1 U796 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U797 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U798 ( .A1(n744), .A2(G898), .ZN(n745) );
  XOR2_X1 U799 ( .A(n747), .B(n748), .Z(n750) );
  XNOR2_X1 U800 ( .A(n750), .B(n749), .ZN(n754) );
  XNOR2_X1 U801 ( .A(KEYINPUT125), .B(n754), .ZN(n751) );
  XNOR2_X1 U802 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U803 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U804 ( .A1(n753), .A2(G953), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n395), .B(n754), .ZN(n756) );
  NAND2_X1 U806 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U807 ( .A1(n758), .A2(n757), .ZN(G72) );
  XOR2_X1 U808 ( .A(G131), .B(KEYINPUT126), .Z(n759) );
  XNOR2_X1 U809 ( .A(n760), .B(n759), .ZN(G33) );
  XOR2_X1 U810 ( .A(n408), .B(G137), .Z(G39) );
endmodule

