//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n189));
  OR2_X1    g003(.A1(KEYINPUT72), .A2(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(KEYINPUT72), .A2(G125), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(G140), .A3(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(G125), .A2(G140), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT72), .B(G125), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n188), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT72), .A2(G125), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT72), .A2(G125), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G140), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n189), .A3(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n193), .B1(new_n201), .B2(G140), .ZN(new_n204));
  OAI211_X1 g018(.A(G146), .B(new_n203), .C1(new_n204), .C2(new_n189), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  INV_X1    g022(.A(G237), .ZN(new_n209));
  NAND2_X1  g023(.A1(KEYINPUT69), .A2(G953), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT69), .A2(G953), .ZN(new_n212));
  OAI211_X1 g026(.A(G214), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G143), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(KEYINPUT69), .A2(G953), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n217), .A2(G143), .A3(G214), .A4(new_n209), .ZN(new_n218));
  AOI211_X1 g032(.A(new_n207), .B(new_n208), .C1(new_n215), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n187), .B1(new_n206), .B2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n215), .A2(new_n218), .A3(new_n208), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT81), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(G237), .B1(new_n216), .B2(new_n210), .ZN(new_n224));
  AOI21_X1  g038(.A(G143), .B1(new_n224), .B2(G214), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n213), .A2(new_n214), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n215), .A2(new_n218), .A3(KEYINPUT81), .A4(new_n208), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n223), .A2(new_n227), .A3(new_n207), .A4(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT17), .B(G131), .C1(new_n225), .C2(new_n226), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n230), .A2(KEYINPUT85), .A3(new_n198), .A4(new_n205), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n220), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n215), .B(new_n218), .C1(new_n233), .C2(new_n208), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n204), .A2(G146), .ZN(new_n235));
  XNOR2_X1  g049(.A(G125), .B(G140), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n188), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n234), .B(new_n238), .C1(new_n227), .C2(new_n233), .ZN(new_n239));
  XOR2_X1   g053(.A(G113), .B(G122), .Z(new_n240));
  XNOR2_X1  g054(.A(new_n240), .B(KEYINPUT84), .ZN(new_n241));
  INV_X1    g055(.A(G104), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n232), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n232), .A2(KEYINPUT86), .A3(new_n239), .A4(new_n243), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n223), .A2(new_n227), .A3(new_n228), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT83), .B(KEYINPUT19), .Z(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n236), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n204), .A2(KEYINPUT19), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(KEYINPUT82), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n205), .B(new_n249), .C1(new_n255), .C2(G146), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n243), .B1(new_n256), .B2(new_n239), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n248), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n260));
  NOR2_X1   g074(.A1(G475), .A2(G902), .ZN(new_n261));
  XNOR2_X1  g075(.A(new_n261), .B(KEYINPUT87), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n257), .B1(new_n246), .B2(new_n247), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT20), .B1(new_n265), .B2(new_n262), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n232), .A2(new_n239), .ZN(new_n267));
  INV_X1    g081(.A(new_n243), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n248), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n264), .A2(new_n266), .B1(new_n272), .B2(G475), .ZN(new_n273));
  XOR2_X1   g087(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G143), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n274), .B(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT66), .B(G128), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n278), .A2(new_n214), .ZN(new_n279));
  OAI21_X1  g093(.A(G134), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT89), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n279), .A2(G134), .A3(new_n276), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n282), .B(KEYINPUT90), .ZN(new_n283));
  INV_X1    g097(.A(G116), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G122), .ZN(new_n285));
  INV_X1    g099(.A(G122), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(G116), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G107), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n288), .B(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n291), .B(G134), .C1(new_n277), .C2(new_n279), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n281), .A2(new_n283), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT14), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n295), .B(KEYINPUT91), .ZN(new_n296));
  INV_X1    g110(.A(new_n285), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n287), .B2(new_n294), .ZN(new_n298));
  OAI21_X1  g112(.A(G107), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n288), .A2(new_n289), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n279), .A2(new_n276), .ZN(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n299), .B(new_n300), .C1(new_n282), .C2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(KEYINPUT9), .B(G234), .Z(new_n305));
  INV_X1    g119(.A(G953), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(G217), .A3(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(new_n307), .B(KEYINPUT92), .Z(new_n308));
  NAND3_X1  g122(.A1(new_n293), .A2(new_n304), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n293), .B2(new_n304), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n271), .ZN(new_n313));
  INV_X1    g127(.A(G478), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT15), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n313), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G952), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n318), .A2(KEYINPUT93), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(KEYINPUT93), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n306), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(G234), .B2(G237), .ZN(new_n322));
  INV_X1    g136(.A(new_n217), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n271), .B1(G234), .B2(G237), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(KEYINPUT94), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT21), .B(G898), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n322), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n273), .A2(new_n317), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n188), .A2(G143), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n214), .A2(G146), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .A4(G128), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G143), .B(G146), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n337), .A2(KEYINPUT77), .A3(new_n333), .A4(G128), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n331), .A2(new_n332), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n333), .B1(G143), .B2(new_n188), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n275), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT3), .B1(new_n242), .B2(G107), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(new_n289), .A3(G104), .ZN(new_n345));
  INV_X1    g159(.A(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n242), .A2(G107), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n345), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n289), .A2(G104), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n242), .A2(G107), .ZN(new_n350));
  OAI21_X1  g164(.A(G101), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT66), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G128), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n339), .B1(new_n358), .B2(new_n340), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n354), .B1(new_n359), .B2(new_n334), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n353), .A2(new_n354), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT11), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n302), .B2(G137), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n302), .A2(G137), .ZN(new_n364));
  INV_X1    g178(.A(G137), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT11), .A3(G134), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G131), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n363), .A2(new_n366), .A3(new_n208), .A4(new_n364), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(KEYINPUT68), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n343), .A2(new_n345), .A3(new_n347), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT76), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT76), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n343), .A2(new_n345), .A3(new_n377), .A4(new_n347), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(G101), .A3(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n348), .A2(KEYINPUT4), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT0), .A2(G128), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n337), .B2(KEYINPUT64), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G128), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT64), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n339), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n376), .A2(new_n388), .A3(G101), .A4(new_n378), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n361), .A2(new_n374), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n361), .A2(new_n390), .A3(new_n374), .A4(KEYINPUT78), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n217), .A2(G227), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G140), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n359), .A2(new_n334), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n353), .B1(new_n400), .B2(new_n352), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n370), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT12), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n401), .B1(KEYINPUT79), .B2(KEYINPUT12), .ZN(new_n404));
  INV_X1    g218(.A(new_n374), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n404), .B(new_n405), .C1(KEYINPUT79), .C2(new_n401), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n395), .A2(new_n399), .A3(new_n403), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n374), .B1(new_n361), .B2(new_n390), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n393), .B2(new_n394), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n407), .B1(new_n409), .B2(new_n399), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G469), .ZN(new_n411));
  INV_X1    g225(.A(G469), .ZN(new_n412));
  AND4_X1   g226(.A1(new_n395), .A2(new_n398), .A3(new_n403), .A4(new_n406), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n409), .A2(new_n398), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n412), .B(new_n271), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(G469), .A2(G902), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n411), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(G214), .B1(G237), .B2(G902), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(G116), .B(G119), .Z(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT2), .B(G113), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n381), .A2(new_n422), .A3(new_n389), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n284), .A2(KEYINPUT5), .A3(G119), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT80), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n425), .B(G113), .C1(new_n426), .C2(new_n420), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n420), .A2(new_n421), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(new_n352), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  XOR2_X1   g244(.A(G110), .B(G122), .Z(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n423), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n400), .A2(new_n196), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n387), .A2(new_n201), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G224), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G953), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n440), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n430), .A2(new_n444), .A3(new_n431), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n435), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n441), .B(new_n442), .C1(KEYINPUT7), .C2(new_n440), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n427), .A2(new_n428), .ZN(new_n448));
  INV_X1    g262(.A(new_n352), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n429), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n431), .B(KEYINPUT8), .Z(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  OR3_X1    g267(.A1(new_n438), .A2(KEYINPUT7), .A3(new_n440), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n447), .A2(new_n453), .A3(new_n434), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n446), .A2(new_n271), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n446), .A2(new_n455), .A3(new_n271), .A4(new_n457), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n419), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G221), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n305), .B2(new_n271), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n417), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  OR3_X1    g279(.A1(new_n330), .A2(KEYINPUT95), .A3(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT29), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n372), .A2(new_n387), .A3(new_n373), .ZN(new_n468));
  INV_X1    g282(.A(new_n422), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n365), .A2(G134), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n208), .B1(new_n364), .B2(new_n470), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n359), .A2(new_n334), .B1(KEYINPUT65), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n369), .A2(KEYINPUT65), .ZN(new_n473));
  INV_X1    g287(.A(new_n471), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(KEYINPUT28), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT71), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n472), .A2(new_n475), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n370), .A2(new_n387), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n422), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(G101), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n224), .A2(G210), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n484), .B(new_n485), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n478), .A2(new_n479), .A3(new_n482), .A4(new_n486), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n478), .A2(new_n482), .A3(new_n486), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n489), .B(new_n490), .C1(new_n480), .C2(new_n481), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n472), .A2(new_n475), .B1(new_n370), .B2(new_n387), .ZN(new_n492));
  OAI21_X1  g306(.A(KEYINPUT67), .B1(new_n492), .B2(KEYINPUT30), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n468), .A2(KEYINPUT30), .A3(new_n476), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n491), .A2(new_n493), .A3(new_n494), .A4(new_n422), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n477), .ZN(new_n496));
  INV_X1    g310(.A(new_n486), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT71), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n467), .B(new_n487), .C1(new_n488), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n468), .A2(new_n476), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n422), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n478), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n497), .A2(new_n467), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G472), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT32), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT31), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n509), .B1(new_n496), .B2(new_n497), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n495), .A2(KEYINPUT31), .A3(new_n477), .A4(new_n486), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n478), .A2(new_n482), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n497), .ZN(new_n513));
  NOR2_X1   g327(.A1(G472), .A2(G902), .ZN(new_n514));
  XOR2_X1   g328(.A(new_n514), .B(KEYINPUT70), .Z(new_n515));
  OAI21_X1  g329(.A(new_n508), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n510), .A2(new_n511), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n497), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n515), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT32), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n507), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n275), .A2(G119), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n278), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G110), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT23), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n526), .B2(G128), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n524), .B1(new_n358), .B2(G119), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(new_n530), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n533), .B2(G110), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n206), .ZN(new_n535));
  INV_X1    g349(.A(G110), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n536), .B(new_n531), .C1(new_n532), .C2(new_n530), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(new_n528), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(KEYINPUT73), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n539), .A2(new_n205), .A3(new_n237), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT73), .B1(new_n537), .B2(new_n538), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT22), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(G137), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n545), .B(new_n365), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(new_n535), .C1(new_n541), .C2(new_n540), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n547), .A2(new_n549), .A3(new_n271), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT25), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT25), .A4(new_n271), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n555), .A3(new_n551), .ZN(new_n556));
  INV_X1    g370(.A(G217), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(G234), .B2(new_n271), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n523), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n552), .A2(KEYINPUT74), .A3(new_n553), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n561), .A2(KEYINPUT75), .A3(new_n556), .A4(new_n558), .ZN(new_n562));
  OR2_X1    g376(.A1(new_n550), .A2(new_n558), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AND2_X1   g378(.A1(new_n522), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT95), .B1(new_n330), .B2(new_n465), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n466), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(G101), .ZN(G3));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n464), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n513), .A2(G902), .ZN(new_n570));
  INV_X1    g384(.A(G472), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n513), .A2(new_n515), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n569), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n417), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT96), .Z(new_n578));
  AOI22_X1  g392(.A1(new_n246), .A2(new_n247), .B1(new_n268), .B2(new_n267), .ZN(new_n579));
  OAI21_X1  g393(.A(G475), .B1(new_n579), .B2(G902), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n260), .B1(new_n259), .B2(new_n263), .ZN(new_n581));
  NOR3_X1   g395(.A1(new_n265), .A2(KEYINPUT20), .A3(new_n262), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n311), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT33), .B1(new_n584), .B2(new_n309), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n310), .A2(new_n586), .A3(new_n311), .ZN(new_n587));
  OAI211_X1 g401(.A(G478), .B(new_n271), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n313), .A2(new_n314), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n461), .A2(new_n329), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n578), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT34), .B(G104), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  OAI21_X1  g409(.A(KEYINPUT97), .B1(new_n581), .B2(new_n582), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n313), .B(new_n315), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT97), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n264), .A2(new_n598), .A3(new_n266), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n596), .A2(new_n597), .A3(new_n580), .A4(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n578), .A2(new_n592), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT35), .B(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  NOR2_X1   g417(.A1(new_n546), .A2(KEYINPUT36), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(new_n542), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n605), .B(new_n271), .C1(new_n557), .C2(G234), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n560), .A2(new_n562), .A3(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n466), .A2(new_n566), .A3(new_n574), .A4(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n608), .B(KEYINPUT37), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n536), .ZN(G12));
  AND3_X1   g424(.A1(new_n417), .A2(new_n461), .A3(new_n464), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n611), .A2(new_n522), .A3(new_n607), .ZN(new_n612));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n322), .B1(new_n326), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n596), .A2(new_n580), .A3(new_n599), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n317), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G128), .ZN(G30));
  XOR2_X1   g433(.A(new_n614), .B(KEYINPUT39), .Z(new_n620));
  NAND3_X1  g434(.A1(new_n417), .A2(new_n464), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT40), .Z(new_n622));
  NAND2_X1  g436(.A1(new_n459), .A2(new_n460), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT38), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n496), .A2(new_n497), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n486), .B1(new_n501), .B2(new_n477), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n271), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(G472), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n521), .A2(new_n516), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n583), .A2(new_n597), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n607), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n622), .A2(new_n418), .A3(new_n624), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G143), .ZN(G45));
  NAND3_X1  g448(.A1(new_n583), .A2(new_n590), .A3(new_n615), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n612), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G146), .ZN(G48));
  NOR2_X1   g452(.A1(new_n591), .A2(new_n592), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n271), .B1(new_n413), .B2(new_n414), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G469), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT98), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n415), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(KEYINPUT98), .A3(G469), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n640), .B1(new_n646), .B2(new_n464), .ZN(new_n647));
  AOI211_X1 g461(.A(KEYINPUT99), .B(new_n463), .C1(new_n644), .C2(new_n645), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n565), .B(new_n639), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT41), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(G113), .ZN(G15));
  NOR2_X1   g465(.A1(new_n600), .A2(new_n592), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n565), .B(new_n652), .C1(new_n647), .C2(new_n648), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G116), .ZN(G18));
  INV_X1    g468(.A(new_n461), .ZN(new_n655));
  AOI211_X1 g469(.A(new_n463), .B(new_n655), .C1(new_n645), .C2(new_n644), .ZN(new_n656));
  INV_X1    g470(.A(new_n330), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n656), .A2(new_n522), .A3(new_n657), .A4(new_n607), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G119), .ZN(G21));
  XOR2_X1   g473(.A(new_n515), .B(KEYINPUT100), .Z(new_n660));
  INV_X1    g474(.A(KEYINPUT101), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n486), .B1(new_n502), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n478), .A2(KEYINPUT101), .A3(new_n501), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n664), .B2(new_n517), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n519), .A2(new_n271), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n665), .B1(G472), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n564), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n560), .A2(new_n562), .A3(new_n563), .ZN(new_n670));
  AOI22_X1  g484(.A1(new_n662), .A2(new_n663), .B1(new_n510), .B2(new_n511), .ZN(new_n671));
  OAI22_X1  g485(.A1(new_n570), .A2(new_n571), .B1(new_n671), .B2(new_n660), .ZN(new_n672));
  OAI21_X1  g486(.A(KEYINPUT102), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n328), .B1(new_n669), .B2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n273), .B2(new_n317), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n583), .A2(new_n597), .A3(KEYINPUT103), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n676), .A2(new_n461), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n674), .B(new_n679), .C1(new_n647), .C2(new_n648), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G122), .ZN(G24));
  NAND2_X1  g495(.A1(new_n635), .A2(KEYINPUT104), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n583), .A2(new_n683), .A3(new_n590), .A4(new_n615), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n560), .A2(new_n562), .A3(new_n606), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n672), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n685), .A2(new_n656), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G125), .ZN(G27));
  NOR2_X1   g503(.A1(new_n623), .A2(new_n419), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n416), .B(KEYINPUT105), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n410), .B2(G469), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n463), .B1(new_n693), .B2(new_n415), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI211_X1 g510(.A(KEYINPUT106), .B(new_n463), .C1(new_n693), .C2(new_n415), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n685), .A2(new_n565), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n685), .A2(new_n702), .A3(new_n565), .A4(new_n698), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(new_n573), .B2(KEYINPUT32), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n706), .A2(new_n507), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n521), .A2(new_n516), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(KEYINPUT108), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n670), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n685), .A3(KEYINPUT42), .A4(new_n698), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G131), .ZN(G33));
  AND3_X1   g527(.A1(new_n565), .A2(new_n698), .A3(new_n617), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(new_n302), .ZN(G36));
  NAND2_X1  g529(.A1(new_n273), .A2(new_n590), .ZN(new_n716));
  XOR2_X1   g530(.A(new_n716), .B(KEYINPUT43), .Z(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n575), .A3(new_n607), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n719));
  OR2_X1    g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n410), .B(KEYINPUT45), .Z(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n691), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n691), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n415), .A3(new_n726), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n727), .A2(new_n464), .A3(new_n620), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n718), .A2(new_n719), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n690), .B(KEYINPUT109), .Z(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n720), .A2(new_n728), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G137), .ZN(G39));
  NAND3_X1  g547(.A1(new_n727), .A2(KEYINPUT47), .A3(new_n464), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(KEYINPUT47), .B1(new_n727), .B2(new_n464), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n636), .B(new_n690), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n522), .A2(new_n564), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G140), .ZN(G42));
  AND2_X1   g555(.A1(new_n717), .A2(new_n322), .ZN(new_n742));
  INV_X1    g556(.A(new_n646), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n463), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n669), .A2(new_n673), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n624), .A2(new_n418), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n742), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  XOR2_X1   g561(.A(new_n747), .B(KEYINPUT50), .Z(new_n748));
  INV_X1    g562(.A(new_n690), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n743), .A2(new_n463), .A3(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n750), .A2(new_n564), .A3(new_n322), .A4(new_n630), .ZN(new_n751));
  OR3_X1    g565(.A1(new_n751), .A2(new_n583), .A3(new_n590), .ZN(new_n752));
  INV_X1    g566(.A(new_n736), .ZN(new_n753));
  OAI211_X1 g567(.A(new_n734), .B(new_n753), .C1(new_n464), .C2(new_n743), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n742), .A2(new_n745), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n730), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n742), .A2(new_n750), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n754), .A2(new_n756), .B1(new_n687), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n748), .A2(new_n752), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n321), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n710), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(KEYINPUT48), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n763), .A2(KEYINPUT116), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(KEYINPUT116), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT115), .B1(new_n762), .B2(KEYINPUT48), .ZN(new_n766));
  OR3_X1    g580(.A1(new_n762), .A2(KEYINPUT115), .A3(KEYINPUT48), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n748), .A2(new_n758), .A3(KEYINPUT51), .A4(new_n752), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n761), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n612), .B1(new_n617), .B2(new_n636), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n693), .A2(new_n415), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n464), .A3(new_n615), .ZN(new_n773));
  NOR3_X1   g587(.A1(new_n630), .A2(new_n773), .A3(new_n607), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n655), .B1(new_n631), .B2(new_n675), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n774), .A2(KEYINPUT112), .A3(new_n677), .A4(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n463), .B(new_n614), .C1(new_n693), .C2(new_n415), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n686), .A2(new_n629), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n678), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n771), .A2(new_n776), .A3(new_n688), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n771), .A2(new_n688), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n776), .A2(new_n780), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT52), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n712), .A2(new_n782), .A3(new_n786), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n677), .B(new_n775), .C1(new_n647), .C2(new_n648), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n668), .B1(new_n564), .B2(new_n667), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n670), .A2(new_n672), .A3(KEYINPUT102), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n329), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n653), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n649), .A2(new_n658), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n685), .A2(new_n687), .A3(new_n698), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n685), .A2(KEYINPUT111), .A3(new_n687), .A4(new_n698), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n714), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n592), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n591), .B1(new_n317), .B2(new_n583), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n576), .A2(new_n417), .A3(new_n800), .A4(new_n801), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n802), .A2(new_n608), .A3(new_n567), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n417), .A2(new_n464), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n616), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n749), .A2(new_n597), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n805), .A2(new_n522), .A3(new_n607), .A4(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n794), .A2(new_n799), .A3(new_n803), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n787), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n787), .B2(new_n808), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT54), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n751), .A2(new_n591), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n811), .A2(new_n815), .ZN(new_n816));
  AND4_X1   g630(.A1(KEYINPUT53), .A2(new_n712), .A3(new_n782), .A4(new_n786), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n649), .A2(new_n658), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n680), .A3(new_n819), .A4(new_n653), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT114), .B1(new_n792), .B2(new_n793), .ZN(new_n821));
  AND4_X1   g635(.A1(new_n807), .A2(new_n820), .A3(new_n821), .A4(new_n799), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n822), .A3(new_n803), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT113), .B(new_n809), .C1(new_n787), .C2(new_n808), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n816), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT54), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n770), .A2(new_n813), .A3(new_n814), .A4(new_n826), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n755), .A2(new_n463), .A3(new_n655), .A4(new_n743), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n827), .A2(new_n828), .B1(G952), .B2(G953), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n569), .A2(new_n419), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT110), .Z(new_n831));
  INV_X1    g645(.A(KEYINPUT49), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n273), .B(new_n590), .C1(new_n646), .C2(new_n832), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n624), .B(new_n833), .C1(new_n832), .C2(new_n646), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n630), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n829), .A2(new_n835), .ZN(G75));
  AND2_X1   g650(.A1(new_n435), .A2(new_n445), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT117), .Z(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n825), .A2(G210), .A3(G902), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n443), .B(KEYINPUT55), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n839), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n840), .A2(new_n841), .ZN(new_n846));
  INV_X1    g660(.A(new_n842), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n838), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n217), .A2(G952), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n845), .A2(new_n850), .A3(new_n852), .ZN(G51));
  XNOR2_X1  g667(.A(new_n825), .B(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n691), .A2(KEYINPUT57), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n691), .A2(KEYINPUT57), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n413), .A2(new_n414), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n825), .A2(G469), .A3(G902), .A4(new_n721), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n851), .B1(new_n859), .B2(new_n860), .ZN(G54));
  NAND4_X1  g675(.A1(new_n825), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT118), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(new_n863), .A3(new_n265), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n852), .B1(new_n862), .B2(new_n265), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n862), .B2(new_n265), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G60));
  OR2_X1    g681(.A1(new_n585), .A2(new_n587), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n854), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(G478), .A2(G902), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT59), .Z(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n826), .B2(new_n813), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n852), .B1(new_n873), .B2(new_n868), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(G63));
  NAND2_X1  g689(.A1(G217), .A2(G902), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT60), .Z(new_n877));
  NAND2_X1  g691(.A1(new_n825), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n547), .A2(new_n549), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n605), .B(KEYINPUT119), .Z(new_n881));
  NAND3_X1  g695(.A1(new_n825), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n880), .A2(new_n852), .A3(new_n882), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g698(.A(G953), .B1(new_n327), .B2(new_n439), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(KEYINPUT120), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n794), .A2(new_n803), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n886), .B1(new_n887), .B2(new_n217), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(KEYINPUT120), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n839), .B1(G898), .B2(new_n217), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(G69));
  NAND2_X1  g706(.A1(G227), .A2(G900), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n728), .A2(new_n679), .A3(new_n710), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n732), .B(new_n894), .C1(new_n737), .C2(new_n739), .ZN(new_n895));
  INV_X1    g709(.A(new_n714), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n712), .A2(new_n896), .A3(new_n783), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n217), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT122), .B1(new_n217), .B2(G900), .ZN(new_n899));
  OR3_X1    g713(.A1(new_n217), .A2(KEYINPUT122), .A3(G900), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(KEYINPUT123), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n255), .B(KEYINPUT121), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n491), .A2(new_n493), .A3(new_n494), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n323), .B(new_n893), .C1(new_n904), .C2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n902), .B2(new_n903), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n323), .A2(new_n893), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n740), .A2(new_n732), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n783), .A2(new_n633), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n565), .A2(new_n801), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n621), .A2(new_n749), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n908), .B1(new_n919), .B2(new_n323), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n910), .A2(new_n911), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n909), .A2(new_n921), .ZN(G72));
  XNOR2_X1  g736(.A(KEYINPUT124), .B(KEYINPUT63), .ZN(new_n923));
  NAND2_X1  g737(.A1(G472), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT125), .Z(new_n926));
  OAI21_X1  g740(.A(new_n926), .B1(new_n918), .B2(new_n887), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n496), .B(KEYINPUT126), .Z(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n927), .A2(new_n486), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n496), .A2(new_n497), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT127), .Z(new_n932));
  OAI211_X1 g746(.A(new_n812), .B(new_n925), .C1(new_n625), .C2(new_n932), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n895), .A2(new_n897), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n926), .B1(new_n934), .B2(new_n887), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n497), .A3(new_n928), .ZN(new_n936));
  AND4_X1   g750(.A1(new_n852), .A2(new_n930), .A3(new_n933), .A4(new_n936), .ZN(G57));
endmodule


