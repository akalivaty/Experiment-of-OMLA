//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:50 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  XOR2_X1   g007(.A(KEYINPUT66), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT68), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n459), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G101), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n467), .B2(new_n468), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT68), .B(G2105), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n477), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(G2105), .ZN(new_n485));
  AOI22_X1  g060(.A1(G124), .A2(new_n484), .B1(new_n485), .B2(G136), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n477), .C2(G112), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT69), .ZN(G162));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n492));
  AND2_X1   g067(.A1(G126), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n481), .B2(new_n482), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(G138), .B1(new_n481), .B2(new_n482), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n463), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n467), .A2(new_n468), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n498), .A2(new_n477), .A3(new_n499), .A4(G138), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n495), .B1(new_n497), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G50), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n506), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT6), .B(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(G166));
  INV_X1    g090(.A(KEYINPUT70), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OR2_X1    g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n518), .A2(KEYINPUT70), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n517), .A2(G543), .A3(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G51), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n506), .A2(new_n514), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n524), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n523), .A2(new_n529), .ZN(G168));
  AND2_X1   g105(.A1(new_n506), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G90), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n517), .A2(G52), .A3(G543), .A4(new_n520), .ZN(new_n533));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n504), .B2(new_n505), .ZN(new_n535));
  AND2_X1   g110(.A1(G77), .A2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(G651), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n532), .A2(new_n533), .A3(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(new_n531), .A2(G81), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT71), .B(G43), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n517), .A2(G543), .A3(new_n520), .A4(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n504), .B2(new_n505), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n540), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(G188));
  AOI22_X1  g128(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(G91), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n554), .A2(new_n508), .B1(new_n555), .B2(new_n527), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n517), .A2(G543), .A3(new_n520), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(KEYINPUT72), .ZN(new_n560));
  AOI211_X1 g135(.A(new_n558), .B(new_n560), .C1(KEYINPUT73), .C2(new_n559), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n558), .A2(KEYINPUT73), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n517), .A2(G543), .A3(new_n520), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(new_n560), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n556), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(KEYINPUT74), .ZN(new_n569));
  NAND2_X1  g144(.A1(G166), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n513), .A2(new_n514), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n571), .B1(new_n508), .B2(new_n507), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(KEYINPUT74), .ZN(new_n573));
  AND2_X1   g148(.A1(new_n570), .A2(new_n573), .ZN(G303));
  NAND2_X1  g149(.A1(new_n531), .A2(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n576));
  INV_X1    g151(.A(G49), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n521), .ZN(G288));
  NAND2_X1  g153(.A1(new_n531), .A2(G86), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n580), .B1(new_n504), .B2(new_n505), .ZN(new_n581));
  AND2_X1   g156(.A1(G73), .A2(G543), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n514), .A2(G48), .A3(G543), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n579), .A2(new_n583), .A3(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n511), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n531), .B2(G85), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n557), .A2(G47), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NOR2_X1   g167(.A1(G301), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G92), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n527), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n511), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n594), .A2(new_n597), .B1(new_n600), .B2(G651), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n521), .A2(KEYINPUT75), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT75), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n517), .A2(new_n603), .A3(G543), .A4(new_n520), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(G54), .A3(new_n604), .ZN(new_n605));
  AND3_X1   g180(.A1(new_n601), .A2(new_n605), .A3(KEYINPUT76), .ZN(new_n606));
  AOI21_X1  g181(.A(KEYINPUT76), .B1(new_n601), .B2(new_n605), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n593), .B1(new_n609), .B2(new_n592), .ZN(G284));
  AOI21_X1  g185(.A(new_n593), .B1(new_n609), .B2(new_n592), .ZN(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n566), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(G868), .B2(new_n566), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n547), .A2(new_n592), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n608), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n592), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g195(.A(new_n472), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n498), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  AOI22_X1  g202(.A1(G123), .A2(new_n484), .B1(new_n485), .B2(G135), .ZN(new_n628));
  OAI221_X1 g203(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n477), .C2(G111), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n626), .A2(new_n627), .A3(new_n631), .ZN(G156));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT15), .B(G2435), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT77), .ZN(new_n646));
  INV_X1    g221(.A(G14), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n647), .B1(new_n643), .B2(new_n644), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2072), .B(G2078), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT78), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  OR3_X1    g230(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n653), .B2(new_n655), .ZN(new_n657));
  INV_X1    g232(.A(new_n651), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n652), .B(KEYINPUT17), .Z(new_n659));
  OAI211_X1 g234(.A(new_n656), .B(new_n657), .C1(new_n658), .C2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n655), .A2(new_n651), .A3(new_n652), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT18), .Z(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(new_n655), .A3(new_n658), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(new_n625), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT79), .B(G2096), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT19), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  AND2_X1   g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n670), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(new_n670), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT80), .Z(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1991), .B(G1996), .Z(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  INV_X1    g260(.A(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  AND3_X1   g264(.A1(new_n684), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n684), .B2(new_n688), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(G229));
  NOR2_X1   g267(.A1(G29), .A2(G35), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n693), .B1(G162), .B2(G29), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT29), .ZN(new_n695));
  INV_X1    g270(.A(G2090), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G33), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n477), .A2(G103), .A3(G2104), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT25), .Z(new_n701));
  NAND2_X1  g276(.A1(G115), .A2(G2104), .ZN(new_n702));
  INV_X1    g277(.A(G127), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n483), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n477), .B1(new_n704), .B2(KEYINPUT90), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(KEYINPUT90), .B2(new_n704), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n485), .A2(G139), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n701), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n699), .B1(new_n708), .B2(G29), .ZN(new_n709));
  INV_X1    g284(.A(G2072), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT91), .Z(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT96), .B(KEYINPUT23), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G20), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n713), .B(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G299), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(G1956), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n697), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n698), .A2(G32), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT92), .B(KEYINPUT26), .ZN(new_n721));
  NAND3_X1  g296(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G105), .B2(new_n621), .ZN(new_n724));
  AOI22_X1  g299(.A1(G129), .A2(new_n484), .B1(new_n485), .B2(G141), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n720), .B1(new_n727), .B2(new_n698), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT27), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1996), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n714), .A2(G5), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G171), .B2(new_n714), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT94), .Z(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G1961), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G1961), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n730), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g311(.A1(G168), .A2(new_n714), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n737), .B1(new_n714), .B2(G21), .ZN(new_n738));
  INV_X1    g313(.A(G1966), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT24), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n698), .B1(new_n741), .B2(G34), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(new_n741), .B2(G34), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G160), .B2(G29), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(G2084), .ZN(new_n745));
  XOR2_X1   g320(.A(KEYINPUT31), .B(G11), .Z(new_n746));
  INV_X1    g321(.A(G28), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(KEYINPUT30), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT93), .ZN(new_n749));
  AOI21_X1  g324(.A(G29), .B1(new_n747), .B2(KEYINPUT30), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n630), .B2(new_n698), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G2084), .B2(new_n744), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n548), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G16), .B2(G19), .ZN(new_n755));
  INV_X1    g330(.A(G1341), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n740), .A2(new_n745), .A3(new_n753), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(G27), .A2(G29), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G164), .B2(G29), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT95), .B(G2078), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  OAI22_X1  g337(.A1(new_n738), .A2(new_n739), .B1(new_n756), .B2(new_n755), .ZN(new_n763));
  NOR3_X1   g338(.A1(new_n758), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n698), .A2(G26), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT88), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT28), .ZN(new_n767));
  AOI22_X1  g342(.A1(G128), .A2(new_n484), .B1(new_n485), .B2(G140), .ZN(new_n768));
  OAI221_X1 g343(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n477), .C2(G116), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n770), .A2(KEYINPUT87), .A3(G29), .ZN(new_n771));
  AOI21_X1  g346(.A(KEYINPUT87), .B1(new_n770), .B2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n767), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT89), .B(G2067), .Z(new_n774));
  AOI22_X1  g349(.A1(new_n773), .A2(new_n774), .B1(new_n709), .B2(new_n710), .ZN(new_n775));
  OAI211_X1 g350(.A(new_n764), .B(new_n775), .C1(new_n774), .C2(new_n773), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n719), .A2(new_n736), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(G4), .A2(G16), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n609), .B2(G16), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1348), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n777), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(G288), .A2(KEYINPUT82), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n557), .A2(G49), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT82), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n784), .A2(new_n785), .A3(new_n576), .A4(new_n575), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n714), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n714), .A2(G23), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT33), .B(G1976), .Z(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n789), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n572), .A2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G22), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(G16), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(KEYINPUT83), .ZN(new_n798));
  INV_X1    g373(.A(KEYINPUT83), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n799), .A3(new_n796), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n798), .A2(G1971), .A3(new_n800), .ZN(new_n801));
  MUX2_X1   g376(.A(G6), .B(G305), .S(G16), .Z(new_n802));
  XOR2_X1   g377(.A(KEYINPUT32), .B(G1981), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G1971), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n799), .B1(new_n793), .B2(new_n796), .ZN(new_n806));
  AOI211_X1 g381(.A(KEYINPUT83), .B(new_n795), .C1(new_n572), .C2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n801), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT84), .B1(new_n792), .B2(new_n809), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n801), .A2(new_n804), .A3(new_n808), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n789), .B(new_n790), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT84), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT34), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n698), .A2(G25), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n485), .A2(G131), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT81), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n484), .A2(G119), .ZN(new_n823));
  OAI221_X1 g398(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n477), .C2(G107), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n820), .B1(new_n827), .B2(new_n698), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT35), .B(G1991), .Z(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n828), .B(new_n830), .ZN(new_n831));
  MUX2_X1   g406(.A(G24), .B(G290), .S(G16), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(G1986), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(KEYINPUT85), .B1(new_n819), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(KEYINPUT34), .B1(new_n810), .B2(new_n814), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT85), .ZN(new_n837));
  INV_X1    g412(.A(new_n834), .ZN(new_n838));
  NOR3_X1   g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n818), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(KEYINPUT86), .A2(KEYINPUT36), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n819), .A2(KEYINPUT85), .A3(new_n834), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n818), .A3(new_n841), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n782), .B1(new_n843), .B2(new_n847), .ZN(G311));
  INV_X1    g423(.A(new_n782), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n841), .B1(new_n846), .B2(new_n818), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n817), .B(new_n842), .C1(new_n844), .C2(new_n845), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(G150));
  NAND4_X1  g427(.A1(new_n517), .A2(G55), .A3(G543), .A4(new_n520), .ZN(new_n853));
  INV_X1    g428(.A(G67), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n504), .B2(new_n505), .ZN(new_n855));
  AND2_X1   g430(.A1(G80), .A2(G543), .ZN(new_n856));
  OAI21_X1  g431(.A(G651), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n506), .A2(new_n514), .A3(G93), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(G860), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT98), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n609), .A2(G559), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT38), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n544), .A2(new_n545), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n865), .A2(G651), .B1(G81), .B2(new_n531), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n857), .A2(new_n858), .ZN(new_n867));
  NAND4_X1  g442(.A1(new_n866), .A2(new_n867), .A3(new_n542), .A4(new_n853), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n547), .A2(new_n859), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OR2_X1    g445(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT39), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT97), .Z(new_n874));
  AOI21_X1  g449(.A(KEYINPUT39), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(G860), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n862), .B1(new_n874), .B2(new_n876), .ZN(G145));
  INV_X1    g452(.A(KEYINPUT100), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n770), .B(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n708), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n826), .B(new_n623), .Z(new_n881));
  XNOR2_X1  g456(.A(new_n880), .B(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n495), .ZN(new_n883));
  NOR3_X1   g458(.A1(new_n496), .A2(new_n463), .A3(KEYINPUT4), .ZN(new_n884));
  INV_X1    g459(.A(G138), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(new_n467), .B2(new_n468), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n499), .B1(new_n886), .B2(new_n477), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n883), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n726), .B(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n485), .A2(G142), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT101), .ZN(new_n891));
  INV_X1    g466(.A(G118), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n463), .A2(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(new_n893), .B2(new_n894), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT102), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n897), .B1(new_n484), .B2(G130), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n484), .A2(new_n897), .A3(G130), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n891), .B(new_n896), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n889), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n882), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n882), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n479), .B(KEYINPUT99), .ZN(new_n906));
  XNOR2_X1  g481(.A(G162), .B(new_n906), .ZN(new_n907));
  XOR2_X1   g482(.A(new_n907), .B(new_n630), .Z(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(G37), .ZN(new_n910));
  INV_X1    g485(.A(new_n908), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n903), .A2(new_n904), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n910), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g489(.A1(new_n609), .A2(new_n615), .A3(new_n870), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n618), .A2(new_n870), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n601), .A2(new_n605), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n566), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n557), .A2(new_n561), .B1(new_n564), .B2(new_n560), .ZN(new_n920));
  OAI211_X1 g495(.A(new_n605), .B(new_n601), .C1(new_n920), .C2(new_n556), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT41), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n919), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n923));
  OAI22_X1  g498(.A1(new_n916), .A2(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n618), .A2(new_n870), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n919), .A2(new_n921), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n915), .A3(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(KEYINPUT104), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G305), .B1(new_n783), .B2(new_n786), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(new_n572), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n783), .A2(new_n786), .A3(G305), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(G290), .B(G166), .ZN(new_n938));
  INV_X1    g513(.A(new_n936), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(new_n933), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(KEYINPUT104), .B2(new_n928), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n930), .B1(new_n924), .B2(new_n927), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n932), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n924), .A2(new_n927), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n929), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n943), .B1(new_n948), .B2(new_n931), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n859), .A2(new_n592), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(G295));
  OAI21_X1  g527(.A(new_n944), .B1(new_n932), .B2(new_n945), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n948), .A2(new_n943), .A3(new_n931), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n592), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n951), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT105), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n950), .A2(new_n958), .A3(new_n951), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(G331));
  NAND2_X1  g535(.A1(G301), .A2(KEYINPUT106), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n868), .A2(new_n869), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n868), .B2(new_n869), .ZN(new_n963));
  OAI21_X1  g538(.A(G168), .B1(KEYINPUT106), .B2(G301), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n964), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n547), .A2(new_n859), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n547), .A2(new_n859), .ZN(new_n968));
  OAI211_X1 g543(.A(KEYINPUT106), .B(G301), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n868), .A2(new_n869), .A3(new_n961), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI22_X1  g546(.A1(new_n965), .A2(new_n971), .B1(new_n923), .B2(new_n922), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n966), .A3(new_n970), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n926), .A3(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n972), .A2(new_n941), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n972), .A2(new_n941), .A3(new_n978), .A4(new_n975), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n910), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n923), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n922), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n922), .A2(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n974), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n941), .B1(new_n987), .B2(new_n975), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(G37), .B1(new_n976), .B2(KEYINPUT107), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n972), .A2(new_n975), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n942), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n990), .A2(new_n991), .A3(new_n979), .A4(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n989), .A2(KEYINPUT44), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n989), .A2(new_n997), .A3(KEYINPUT44), .A4(new_n994), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n977), .A2(new_n993), .A3(new_n910), .A4(new_n979), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n988), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(new_n991), .A3(new_n979), .A4(new_n990), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1000), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n999), .A2(new_n1009), .ZN(G397));
  INV_X1    g585(.A(G1996), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n726), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n827), .A2(new_n829), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n770), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n826), .A2(new_n830), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n471), .A2(new_n478), .A3(G40), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n471), .A2(new_n478), .A3(KEYINPUT111), .A4(G40), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT45), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1023), .B1(G164), .B2(G1384), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(G290), .A2(G1986), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT112), .ZN(new_n1028));
  AOI211_X1 g603(.A(new_n1022), .B(new_n1024), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G290), .A2(G1986), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1017), .A2(new_n1025), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT126), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G286), .A2(G8), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1038), .A2(new_n1024), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n739), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1041));
  INV_X1    g616(.A(G2084), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n888), .A2(new_n1043), .A3(new_n1037), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1036), .B1(new_n1047), .B2(G8), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT45), .B1(new_n888), .B2(new_n1037), .ZN(new_n1049));
  NOR3_X1   g624(.A1(G164), .A2(new_n1023), .A3(G1384), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(G1966), .B1(new_n1051), .B2(new_n1041), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n1044), .A2(new_n1045), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1053), .A2(G2084), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT125), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT125), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1040), .A2(new_n1046), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(G168), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G8), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1035), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1048), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1034), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1061), .A2(KEYINPUT62), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n783), .A2(new_n786), .A3(G1976), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT52), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n497), .A2(new_n500), .ZN(new_n1067));
  AOI21_X1  g642(.A(G1384), .B1(new_n1067), .B2(new_n883), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1020), .A2(new_n1068), .A3(new_n1021), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT114), .A3(G8), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT114), .B1(new_n1069), .B2(G8), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1064), .B(new_n1066), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n583), .A2(new_n584), .ZN(new_n1074));
  NOR2_X1   g649(.A1(KEYINPUT115), .A2(G86), .ZN(new_n1075));
  AND2_X1   g650(.A1(KEYINPUT115), .A2(G86), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n527), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(G1981), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1981), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n579), .A2(new_n1079), .A3(new_n583), .A4(new_n584), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT116), .B1(new_n1078), .B2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(KEYINPUT49), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  AOI211_X1 g658(.A(KEYINPUT116), .B(new_n1083), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1071), .A2(new_n1072), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1073), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1069), .A2(G8), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1070), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1087), .B1(new_n1091), .B2(new_n1064), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1086), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n570), .A2(new_n573), .A3(G8), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT55), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1039), .A2(new_n805), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1044), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1043), .B1(new_n888), .B2(new_n1037), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT118), .B1(new_n1022), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1045), .A2(new_n1101), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1098), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1097), .B1(new_n1103), .B2(new_n696), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1095), .B1(new_n1104), .B2(new_n1059), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT113), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1053), .A2(G2090), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1097), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT55), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1094), .B(new_n1109), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1096), .B(KEYINPUT113), .C1(G2090), .C2(new_n1053), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(G8), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1039), .B2(G2078), .ZN(new_n1114));
  INV_X1    g689(.A(G1961), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1053), .A2(new_n1115), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1113), .A2(G2078), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1114), .B(new_n1116), .C1(new_n1039), .C2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(G171), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1093), .A2(new_n1105), .A3(new_n1112), .A4(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1033), .B1(new_n1063), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1062), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1122), .B(new_n1123), .C1(new_n1124), .C2(new_n1048), .ZN(new_n1125));
  AND4_X1   g700(.A1(new_n1105), .A2(new_n1093), .A3(new_n1112), .A4(new_n1119), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1122), .B1(new_n1124), .B2(new_n1048), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT62), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1121), .A2(new_n1127), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1047), .A2(G8), .A3(G168), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT119), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1047), .A2(new_n1133), .A3(G8), .A4(G168), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(new_n1093), .A3(new_n1105), .A4(new_n1112), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1137), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1108), .A2(G8), .A3(new_n1111), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(new_n1095), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1139), .A2(new_n1112), .A3(new_n1141), .A4(new_n1093), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1138), .A2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1112), .A2(new_n1092), .A3(new_n1086), .ZN(new_n1144));
  INV_X1    g719(.A(G288), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1085), .A2(new_n1065), .A3(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1080), .B(KEYINPUT117), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1091), .B2(new_n1148), .ZN(new_n1149));
  XOR2_X1   g724(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT56), .B(G2072), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1051), .A2(new_n1041), .A3(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1152), .B1(new_n1103), .B2(G1956), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n920), .B(KEYINPUT120), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n556), .A2(KEYINPUT121), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n556), .A2(KEYINPUT121), .ZN(new_n1156));
  NOR3_X1   g731(.A1(new_n1155), .A2(new_n1156), .A3(KEYINPUT57), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1154), .A2(new_n1157), .B1(KEYINPUT57), .B2(G299), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1153), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1158), .B(new_n1152), .C1(new_n1103), .C2(G1956), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1150), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(G1348), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1053), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1041), .A2(new_n1014), .A3(new_n1068), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(KEYINPUT60), .A3(new_n1165), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(new_n609), .A3(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(KEYINPUT123), .B(KEYINPUT58), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(G1341), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1069), .A2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(new_n1039), .B2(G1996), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1174), .A2(KEYINPUT59), .A3(new_n548), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n608), .A2(new_n1164), .A3(KEYINPUT60), .A4(new_n1165), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT59), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1174), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1177), .B1(new_n1178), .B2(new_n547), .ZN(new_n1179));
  NAND4_X1  g754(.A1(new_n1170), .A2(new_n1175), .A3(new_n1176), .A4(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1162), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT122), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1153), .A2(new_n1182), .ZN(new_n1183));
  OAI211_X1 g758(.A(KEYINPUT122), .B(new_n1152), .C1(new_n1103), .C2(G1956), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1183), .A2(new_n1184), .A3(new_n1159), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(KEYINPUT61), .A3(new_n1161), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1166), .A2(new_n609), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g763(.A1(new_n1181), .A2(new_n1186), .B1(new_n1188), .B2(new_n1161), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1093), .A2(new_n1105), .A3(new_n1112), .ZN(new_n1190));
  XNOR2_X1  g765(.A(G301), .B(KEYINPUT54), .ZN(new_n1191));
  AND2_X1   g766(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1018), .A2(new_n1117), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1191), .B1(new_n1051), .B2(new_n1193), .ZN(new_n1194));
  AOI22_X1  g769(.A1(new_n1118), .A2(new_n1191), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1128), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1196));
  OAI211_X1 g771(.A(new_n1143), .B(new_n1149), .C1(new_n1189), .C2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1032), .B1(new_n1130), .B2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1017), .A2(new_n1025), .ZN(new_n1199));
  AND2_X1   g774(.A1(new_n1025), .A2(new_n1030), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(KEYINPUT48), .ZN(new_n1201));
  OR2_X1    g776(.A1(new_n1200), .A2(KEYINPUT48), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1204));
  OAI22_X1  g779(.A1(new_n1204), .A2(new_n1013), .B1(G2067), .B2(new_n770), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1025), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT47), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1015), .A2(new_n727), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1025), .A2(new_n1011), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT46), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1208), .A2(new_n1025), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1211), .B1(new_n1210), .B2(new_n1209), .ZN(new_n1212));
  OAI211_X1 g787(.A(new_n1203), .B(new_n1206), .C1(new_n1207), .C2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1213), .B1(new_n1207), .B2(new_n1212), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1198), .A2(new_n1214), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g790(.A(G229), .ZN(new_n1217));
  INV_X1    g791(.A(G319), .ZN(new_n1218));
  NOR2_X1   g792(.A1(G227), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g793(.A(new_n1219), .B(KEYINPUT127), .ZN(new_n1220));
  AOI21_X1  g794(.A(new_n1220), .B1(new_n646), .B2(new_n648), .ZN(new_n1221));
  AND4_X1   g795(.A1(new_n1217), .A2(new_n1007), .A3(new_n913), .A4(new_n1221), .ZN(G308));
  NAND4_X1  g796(.A1(new_n1217), .A2(new_n1007), .A3(new_n913), .A4(new_n1221), .ZN(G225));
endmodule


