

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  NOR2_X1 U322 ( .A1(n465), .A2(n464), .ZN(n477) );
  XNOR2_X1 U323 ( .A(n469), .B(n468), .ZN(n506) );
  XNOR2_X1 U324 ( .A(n467), .B(KEYINPUT97), .ZN(n468) );
  XOR2_X1 U325 ( .A(n429), .B(n428), .Z(n290) );
  XNOR2_X1 U326 ( .A(n344), .B(n343), .ZN(n346) );
  INV_X1 U327 ( .A(G176GAT), .ZN(n432) );
  XNOR2_X1 U328 ( .A(n346), .B(n345), .ZN(n348) );
  XNOR2_X1 U329 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U330 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U331 ( .A(n435), .B(n434), .ZN(n439) );
  NOR2_X1 U332 ( .A1(n426), .A2(n488), .ZN(n565) );
  XNOR2_X1 U333 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U334 ( .A(n447), .B(n446), .Z(n512) );
  XNOR2_X1 U335 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U336 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U337 ( .A(n454), .B(n453), .ZN(G1349GAT) );
  XNOR2_X1 U338 ( .A(n474), .B(n473), .ZN(G1330GAT) );
  XNOR2_X1 U339 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n291), .B(KEYINPUT13), .ZN(n365) );
  XNOR2_X1 U341 ( .A(G99GAT), .B(G85GAT), .ZN(n292) );
  XNOR2_X1 U342 ( .A(n292), .B(KEYINPUT69), .ZN(n322) );
  XOR2_X1 U343 ( .A(n365), .B(n322), .Z(n297) );
  XOR2_X1 U344 ( .A(G78GAT), .B(G148GAT), .Z(n294) );
  XNOR2_X1 U345 ( .A(G106GAT), .B(G204GAT), .ZN(n293) );
  XNOR2_X1 U346 ( .A(n294), .B(n293), .ZN(n317) );
  XNOR2_X1 U347 ( .A(G176GAT), .B(G92GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n295), .B(G64GAT), .ZN(n396) );
  XNOR2_X1 U349 ( .A(n317), .B(n396), .ZN(n296) );
  XNOR2_X1 U350 ( .A(n297), .B(n296), .ZN(n304) );
  XOR2_X1 U351 ( .A(G120GAT), .B(G71GAT), .Z(n429) );
  XOR2_X1 U352 ( .A(KEYINPUT70), .B(KEYINPUT31), .Z(n299) );
  XNOR2_X1 U353 ( .A(KEYINPUT32), .B(KEYINPUT33), .ZN(n298) );
  XNOR2_X1 U354 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U355 ( .A(n429), .B(n300), .Z(n302) );
  NAND2_X1 U356 ( .A1(G230GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n571) );
  XOR2_X1 U359 ( .A(KEYINPUT41), .B(n571), .Z(n525) );
  INV_X1 U360 ( .A(n525), .ZN(n548) );
  XOR2_X1 U361 ( .A(KEYINPUT86), .B(KEYINPUT24), .Z(n306) );
  XNOR2_X1 U362 ( .A(KEYINPUT22), .B(KEYINPUT84), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n321) );
  XOR2_X1 U364 ( .A(G155GAT), .B(KEYINPUT2), .Z(n308) );
  XNOR2_X1 U365 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U366 ( .A(n308), .B(n307), .ZN(n421) );
  XOR2_X1 U367 ( .A(G50GAT), .B(G162GAT), .Z(n328) );
  XOR2_X1 U368 ( .A(n421), .B(n328), .Z(n310) );
  NAND2_X1 U369 ( .A1(G228GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U371 ( .A(KEYINPUT85), .B(KEYINPUT83), .Z(n312) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U374 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U375 ( .A(G211GAT), .B(KEYINPUT21), .Z(n316) );
  XNOR2_X1 U376 ( .A(G197GAT), .B(G218GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n400) );
  XNOR2_X1 U378 ( .A(n317), .B(n400), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U380 ( .A(n321), .B(n320), .Z(n461) );
  XOR2_X1 U381 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n402) );
  XNOR2_X1 U382 ( .A(G92GAT), .B(n322), .ZN(n324) );
  NAND2_X1 U383 ( .A1(G232GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U384 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U385 ( .A(G36GAT), .B(G190GAT), .Z(n395) );
  XNOR2_X1 U386 ( .A(n325), .B(n395), .ZN(n330) );
  XOR2_X1 U387 ( .A(G29GAT), .B(G43GAT), .Z(n327) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n349) );
  XNOR2_X1 U390 ( .A(n349), .B(n328), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n338) );
  XOR2_X1 U392 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n332) );
  XNOR2_X1 U393 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U395 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n334) );
  XNOR2_X1 U396 ( .A(G134GAT), .B(G106GAT), .ZN(n333) );
  XNOR2_X1 U397 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U398 ( .A(n336), .B(n335), .Z(n337) );
  XOR2_X1 U399 ( .A(n338), .B(n337), .Z(n559) );
  INV_X1 U400 ( .A(n559), .ZN(n534) );
  XOR2_X1 U401 ( .A(G8GAT), .B(G141GAT), .Z(n340) );
  XNOR2_X1 U402 ( .A(G169GAT), .B(G197GAT), .ZN(n339) );
  XNOR2_X1 U403 ( .A(n340), .B(n339), .ZN(n355) );
  XOR2_X1 U404 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n342) );
  XNOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U407 ( .A(G36GAT), .B(G50GAT), .Z(n343) );
  XOR2_X1 U408 ( .A(G113GAT), .B(G1GAT), .Z(n406) );
  XOR2_X1 U409 ( .A(G15GAT), .B(G22GAT), .Z(n362) );
  XNOR2_X1 U410 ( .A(n406), .B(n362), .ZN(n345) );
  AND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n349), .B(KEYINPUT64), .ZN(n351) );
  INV_X1 U414 ( .A(KEYINPUT65), .ZN(n350) );
  XOR2_X1 U415 ( .A(n355), .B(n354), .Z(n523) );
  AND2_X1 U416 ( .A1(n525), .A2(n523), .ZN(n357) );
  XNOR2_X1 U417 ( .A(KEYINPUT106), .B(KEYINPUT46), .ZN(n356) );
  XNOR2_X1 U418 ( .A(n357), .B(n356), .ZN(n358) );
  NOR2_X1 U419 ( .A1(n534), .A2(n358), .ZN(n378) );
  XOR2_X1 U420 ( .A(G64GAT), .B(G155GAT), .Z(n360) );
  XNOR2_X1 U421 ( .A(G78GAT), .B(G211GAT), .ZN(n359) );
  XNOR2_X1 U422 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U423 ( .A(n361), .B(G127GAT), .Z(n364) );
  XNOR2_X1 U424 ( .A(n362), .B(G71GAT), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U426 ( .A(G8GAT), .B(G183GAT), .Z(n393) );
  XOR2_X1 U427 ( .A(n365), .B(n393), .Z(n367) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U430 ( .A(n369), .B(n368), .Z(n377) );
  XOR2_X1 U431 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n371) );
  XNOR2_X1 U432 ( .A(G1GAT), .B(KEYINPUT76), .ZN(n370) );
  XNOR2_X1 U433 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U434 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n373) );
  XNOR2_X1 U435 ( .A(KEYINPUT12), .B(KEYINPUT73), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U438 ( .A(n377), .B(n376), .Z(n530) );
  INV_X1 U439 ( .A(n530), .ZN(n576) );
  NAND2_X1 U440 ( .A1(n378), .A2(n576), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n379), .B(KEYINPUT47), .ZN(n380) );
  XNOR2_X1 U442 ( .A(KEYINPUT107), .B(n380), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n559), .B(KEYINPUT36), .ZN(n579) );
  NOR2_X1 U444 ( .A1(n576), .A2(n579), .ZN(n381) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n381), .Z(n382) );
  NOR2_X1 U446 ( .A1(n571), .A2(n382), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n383), .B(KEYINPUT108), .ZN(n384) );
  INV_X1 U448 ( .A(n523), .ZN(n566) );
  NAND2_X1 U449 ( .A1(n384), .A2(n566), .ZN(n385) );
  NAND2_X1 U450 ( .A1(n386), .A2(n385), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n387), .B(KEYINPUT48), .ZN(n388) );
  XOR2_X1 U452 ( .A(KEYINPUT109), .B(n388), .Z(n542) );
  XOR2_X1 U453 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n390) );
  XNOR2_X1 U454 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n431) );
  XOR2_X1 U456 ( .A(G204GAT), .B(n431), .Z(n392) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U459 ( .A(n394), .B(n393), .Z(n398) );
  XNOR2_X1 U460 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U461 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U462 ( .A(n400), .B(n399), .Z(n510) );
  INV_X1 U463 ( .A(n510), .ZN(n491) );
  NAND2_X1 U464 ( .A1(n542), .A2(n491), .ZN(n401) );
  XNOR2_X1 U465 ( .A(n402), .B(n401), .ZN(n426) );
  XOR2_X1 U466 ( .A(G57GAT), .B(G85GAT), .Z(n404) );
  XNOR2_X1 U467 ( .A(G148GAT), .B(G162GAT), .ZN(n403) );
  XNOR2_X1 U468 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U469 ( .A(n405), .B(G120GAT), .Z(n408) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(n406), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n412) );
  XOR2_X1 U472 ( .A(KEYINPUT91), .B(KEYINPUT93), .Z(n410) );
  XNOR2_X1 U473 ( .A(KEYINPUT87), .B(KEYINPUT89), .ZN(n409) );
  XNOR2_X1 U474 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U476 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n414) );
  XNOR2_X1 U477 ( .A(KEYINPUT92), .B(KEYINPUT88), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n416), .B(n415), .ZN(n425) );
  XOR2_X1 U480 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n418) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U483 ( .A(n419), .B(KEYINPUT90), .Z(n423) );
  XNOR2_X1 U484 ( .A(G134GAT), .B(G127GAT), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n420), .B(KEYINPUT0), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n428), .B(n421), .ZN(n422) );
  XNOR2_X1 U487 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U488 ( .A(n425), .B(n424), .Z(n541) );
  INV_X1 U489 ( .A(n541), .ZN(n488) );
  NAND2_X1 U490 ( .A1(n461), .A2(n565), .ZN(n427) );
  XNOR2_X1 U491 ( .A(n427), .B(KEYINPUT55), .ZN(n448) );
  NAND2_X1 U492 ( .A1(G227GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n290), .B(n430), .ZN(n435) );
  XNOR2_X1 U494 ( .A(n431), .B(KEYINPUT81), .ZN(n433) );
  XOR2_X1 U495 ( .A(G183GAT), .B(G190GAT), .Z(n437) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G99GAT), .ZN(n436) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U498 ( .A(n439), .B(n438), .Z(n447) );
  XOR2_X1 U499 ( .A(KEYINPUT80), .B(KEYINPUT20), .Z(n441) );
  XNOR2_X1 U500 ( .A(KEYINPUT78), .B(KEYINPUT79), .ZN(n440) );
  XNOR2_X1 U501 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U502 ( .A(KEYINPUT82), .B(KEYINPUT77), .Z(n443) );
  XNOR2_X1 U503 ( .A(G113GAT), .B(G15GAT), .ZN(n442) );
  XNOR2_X1 U504 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  INV_X1 U506 ( .A(n512), .ZN(n520) );
  NAND2_X1 U507 ( .A1(n448), .A2(n520), .ZN(n558) );
  NOR2_X1 U508 ( .A1(n548), .A2(n558), .ZN(n454) );
  XOR2_X1 U509 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n450) );
  XNOR2_X1 U510 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT118), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n520), .A2(n491), .ZN(n455) );
  NAND2_X1 U514 ( .A1(n461), .A2(n455), .ZN(n456) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n456), .Z(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT27), .B(n510), .Z(n462) );
  NOR2_X1 U517 ( .A1(n461), .A2(n520), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT26), .ZN(n564) );
  NAND2_X1 U519 ( .A1(n462), .A2(n564), .ZN(n540) );
  NAND2_X1 U520 ( .A1(n458), .A2(n540), .ZN(n459) );
  NAND2_X1 U521 ( .A1(n459), .A2(n541), .ZN(n460) );
  XOR2_X1 U522 ( .A(KEYINPUT94), .B(n460), .Z(n465) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT28), .ZN(n516) );
  AND2_X1 U524 ( .A1(n516), .A2(n462), .ZN(n463) );
  NAND2_X1 U525 ( .A1(n463), .A2(n488), .ZN(n522) );
  NOR2_X1 U526 ( .A1(n520), .A2(n522), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n477), .A2(n579), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n466), .A2(n576), .ZN(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT98), .B(KEYINPUT37), .Z(n467) );
  NOR2_X1 U530 ( .A1(n566), .A2(n571), .ZN(n478) );
  NAND2_X1 U531 ( .A1(n506), .A2(n478), .ZN(n470) );
  XOR2_X1 U532 ( .A(KEYINPUT38), .B(n470), .Z(n495) );
  NAND2_X1 U533 ( .A1(n520), .A2(n495), .ZN(n474) );
  XOR2_X1 U534 ( .A(KEYINPUT100), .B(KEYINPUT40), .Z(n472) );
  XNOR2_X1 U535 ( .A(G43GAT), .B(KEYINPUT101), .ZN(n471) );
  NOR2_X1 U536 ( .A1(n576), .A2(n534), .ZN(n475) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NOR2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n497) );
  NAND2_X1 U539 ( .A1(n478), .A2(n497), .ZN(n486) );
  NOR2_X1 U540 ( .A1(n541), .A2(n486), .ZN(n480) );
  XNOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT95), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U544 ( .A1(n510), .A2(n486), .ZN(n482) );
  XOR2_X1 U545 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  NOR2_X1 U546 ( .A1(n512), .A2(n486), .ZN(n484) );
  XNOR2_X1 U547 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n483) );
  XNOR2_X1 U548 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U549 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  NOR2_X1 U550 ( .A1(n516), .A2(n486), .ZN(n487) );
  XOR2_X1 U551 ( .A(G22GAT), .B(n487), .Z(G1327GAT) );
  XOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  NAND2_X1 U553 ( .A1(n495), .A2(n488), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  XOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT99), .Z(n493) );
  NAND2_X1 U556 ( .A1(n495), .A2(n491), .ZN(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1329GAT) );
  INV_X1 U558 ( .A(n516), .ZN(n494) );
  NAND2_X1 U559 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U561 ( .A1(n523), .A2(n548), .ZN(n507) );
  NAND2_X1 U562 ( .A1(n507), .A2(n497), .ZN(n503) );
  NOR2_X1 U563 ( .A1(n541), .A2(n503), .ZN(n499) );
  XNOR2_X1 U564 ( .A(KEYINPUT102), .B(KEYINPUT42), .ZN(n498) );
  XNOR2_X1 U565 ( .A(n499), .B(n498), .ZN(n500) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n500), .Z(G1332GAT) );
  NOR2_X1 U567 ( .A1(n510), .A2(n503), .ZN(n501) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n501), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n512), .A2(n503), .ZN(n502) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n502), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n516), .A2(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n505), .B(n504), .ZN(G1335GAT) );
  NAND2_X1 U574 ( .A1(n507), .A2(n506), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n541), .A2(n515), .ZN(n509) );
  XNOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(G1336GAT) );
  NOR2_X1 U578 ( .A1(n510), .A2(n515), .ZN(n511) );
  XOR2_X1 U579 ( .A(G92GAT), .B(n511), .Z(G1337GAT) );
  NOR2_X1 U580 ( .A1(n512), .A2(n515), .ZN(n513) );
  XOR2_X1 U581 ( .A(KEYINPUT104), .B(n513), .Z(n514) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(n514), .ZN(G1338GAT) );
  NOR2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT105), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n519), .ZN(G1339GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n542), .ZN(n521) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n535), .A2(n523), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT110), .Z(n527) );
  NAND2_X1 U592 ( .A1(n535), .A2(n525), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n528) );
  XNOR2_X1 U595 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT50), .B(KEYINPUT112), .Z(n532) );
  NAND2_X1 U597 ( .A1(n535), .A2(n530), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n533), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n537) );
  NAND2_X1 U601 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n539) );
  XOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT113), .Z(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(n544), .Z(n552) );
  NOR2_X1 U608 ( .A1(n566), .A2(n552), .ZN(n545) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n547) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n548), .A2(n552), .ZN(n549) );
  XOR2_X1 U614 ( .A(n550), .B(n549), .Z(G1345GAT) );
  NOR2_X1 U615 ( .A1(n576), .A2(n552), .ZN(n551) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n551), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n559), .A2(n552), .ZN(n553) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n553), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n566), .A2(n558), .ZN(n554) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n576), .A2(n558), .ZN(n555) );
  XOR2_X1 U622 ( .A(G183GAT), .B(n555), .Z(G1350GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n557) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n561) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(n561), .B(n560), .Z(G1351GAT) );
  XNOR2_X1 U628 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n563) );
  XNOR2_X1 U630 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(n568) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n578) );
  NOR2_X1 U633 ( .A1(n566), .A2(n578), .ZN(n567) );
  XOR2_X1 U634 ( .A(n568), .B(n567), .Z(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U637 ( .A(n578), .ZN(n572) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XOR2_X1 U642 ( .A(G211GAT), .B(n577), .Z(G1354GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

