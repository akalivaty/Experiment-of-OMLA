//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n547, new_n549, new_n550,
    new_n551, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1287,
    new_n1288, new_n1289, new_n1290;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n460), .A2(new_n461), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n466), .B1(G2105), .B2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2105), .B1(new_n460), .B2(new_n461), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g049(.A(KEYINPUT66), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  XOR2_X1   g052(.A(new_n477), .B(KEYINPUT67), .Z(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT68), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n468), .A2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n478), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(KEYINPUT4), .A2(G138), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT3), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(G102), .A2(G2104), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n459), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n488), .B2(new_n489), .ZN(new_n494));
  AND2_X1   g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  OAI21_X1  g070(.A(G2105), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n492), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT69), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n504), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(G88), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(G50), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n504), .A2(new_n506), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n512), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n512), .B(KEYINPUT71), .C1(new_n513), .C2(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(G166));
  NAND2_X1  g095(.A1(new_n509), .A2(G89), .ZN(new_n521));
  AND2_X1   g096(.A1(G63), .A2(G651), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n514), .A2(new_n522), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT6), .B(G651), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n528), .A2(G51), .A3(G543), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n521), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n514), .A2(G64), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n513), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n514), .A2(G90), .A3(new_n528), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n511), .A2(G52), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(new_n514), .A2(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n513), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n514), .A2(G81), .A3(new_n528), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n511), .A2(G43), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT73), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  INV_X1    g127(.A(G65), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n553), .B1(new_n504), .B2(new_n506), .ZN(new_n554));
  AND2_X1   g129(.A1(G78), .A2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(G651), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n514), .A2(G91), .A3(new_n528), .ZN(new_n557));
  AND2_X1   g132(.A1(KEYINPUT6), .A2(G651), .ZN(new_n558));
  NOR2_X1   g133(.A1(KEYINPUT6), .A2(G651), .ZN(new_n559));
  OAI211_X1 g134(.A(G53), .B(G543), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n556), .A2(new_n557), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n560), .A2(new_n561), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n528), .A2(KEYINPUT74), .A3(G53), .A4(G543), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT9), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT75), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n563), .A2(new_n557), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT9), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .A4(new_n556), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n514), .A2(new_n522), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n524), .A2(new_n526), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n577), .A2(new_n529), .A3(new_n578), .ZN(new_n579));
  AND3_X1   g154(.A1(new_n514), .A2(G89), .A3(new_n528), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n521), .A2(new_n527), .A3(KEYINPUT76), .A4(new_n529), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n581), .A2(new_n582), .ZN(G286));
  INV_X1    g158(.A(G166), .ZN(G303));
  NAND2_X1  g159(.A1(new_n509), .A2(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n511), .A2(G49), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n509), .A2(G86), .B1(new_n511), .B2(G48), .ZN(new_n589));
  INV_X1    g164(.A(G61), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n504), .B2(new_n506), .ZN(new_n591));
  AND2_X1   g166(.A1(G73), .A2(G543), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n589), .A2(new_n593), .ZN(G305));
  AOI22_X1  g169(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(new_n513), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n509), .A2(G85), .B1(new_n511), .B2(G47), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n511), .A2(G54), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n514), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n513), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n509), .A2(G92), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n602), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G286), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(new_n573), .ZN(G297));
  AOI21_X1  g187(.A(new_n611), .B1(new_n610), .B2(new_n573), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g194(.A1(new_n476), .A2(G123), .ZN(new_n620));
  XNOR2_X1  g195(.A(KEYINPUT3), .B(G2104), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(new_n459), .ZN(new_n622));
  INV_X1    g197(.A(G135), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n459), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI22_X1  g200(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n620), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT77), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n628), .A2(G2096), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n629), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n642), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT78), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT17), .ZN(new_n658));
  XOR2_X1   g233(.A(G2067), .B(G2678), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n661), .B1(new_n657), .B2(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(new_n660), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n657), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  OR3_X1    g242(.A1(new_n662), .A2(new_n664), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(G2100), .ZN(new_n669));
  XNOR2_X1  g244(.A(KEYINPUT79), .B(G2096), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(G2100), .ZN(new_n671));
  AND3_X1   g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1956), .B(G2474), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT80), .ZN(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n678), .A2(new_n679), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n687));
  OAI211_X1 g262(.A(new_n685), .B(new_n687), .C1(new_n682), .C2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT81), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n692), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n676), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n690), .A2(new_n692), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n675), .A3(new_n693), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G22), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT83), .Z(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G166), .B2(new_n700), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(G1971), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(G23), .ZN(new_n705));
  INV_X1    g280(.A(G288), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n700), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT33), .B(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT34), .ZN(new_n711));
  INV_X1    g286(.A(G305), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G16), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT32), .ZN(new_n714));
  OR2_X1    g289(.A1(G6), .A2(G16), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g293(.A(G1981), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1981), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n720), .A2(new_n721), .A3(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n703), .A2(G1971), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n710), .A2(new_n711), .A3(new_n723), .A4(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n723), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n704), .A2(new_n724), .A3(new_n709), .ZN(new_n727));
  OAI21_X1  g302(.A(KEYINPUT34), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G24), .B(G290), .S(G16), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1986), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n476), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(G95), .A2(G2105), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(KEYINPUT82), .ZN(new_n735));
  INV_X1    g310(.A(G107), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n463), .B1(new_n736), .B2(G2105), .ZN(new_n737));
  AOI22_X1  g312(.A1(G131), .A2(new_n482), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n740), .B(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n730), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n725), .A2(new_n728), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT36), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT36), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n725), .A2(new_n728), .A3(new_n747), .A4(new_n744), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n731), .A2(G35), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n484), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G2090), .ZN(new_n755));
  NAND2_X1  g330(.A1(G171), .A2(G16), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G5), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1961), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(G1341), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n545), .A2(G16), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G16), .B2(G19), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n759), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G160), .A2(new_n731), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n731), .B1(KEYINPUT24), .B2(G34), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(KEYINPUT24), .B2(G34), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT30), .B(G28), .ZN(new_n770));
  OR2_X1    g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n770), .A2(new_n731), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n769), .B(new_n773), .C1(new_n731), .C2(new_n628), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n767), .A2(new_n768), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n763), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n731), .A2(G33), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n621), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n779), .A2(new_n459), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT86), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT85), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n482), .A2(new_n783), .A3(G139), .ZN(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  OAI21_X1  g360(.A(KEYINPUT85), .B1(new_n622), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT25), .Z(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n780), .B2(new_n781), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n778), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G2072), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n700), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n607), .B2(new_n700), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n700), .A2(G21), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G168), .B2(new_n700), .ZN(new_n801));
  OAI22_X1  g376(.A1(new_n757), .A2(new_n758), .B1(G1966), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n760), .B2(new_n762), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n776), .A2(new_n795), .A3(new_n799), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n731), .A2(G27), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G164), .B2(new_n731), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT90), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n807), .A2(G2078), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n731), .A2(G26), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT28), .ZN(new_n810));
  AOI21_X1  g385(.A(KEYINPUT66), .B1(new_n621), .B2(G2105), .ZN(new_n811));
  INV_X1    g386(.A(new_n475), .ZN(new_n812));
  OAI21_X1  g387(.A(G128), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(G140), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT84), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT84), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n621), .A2(new_n816), .A3(G140), .A4(new_n459), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n819));
  INV_X1    g394(.A(G116), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2105), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n813), .A2(new_n818), .A3(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n810), .B1(new_n824), .B2(new_n731), .ZN(new_n825));
  INV_X1    g400(.A(G2067), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n807), .A2(G2078), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n801), .A2(G1966), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT89), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n808), .A2(new_n827), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n804), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT87), .ZN(new_n833));
  OAI21_X1  g408(.A(G129), .B1(new_n811), .B2(new_n812), .ZN(new_n834));
  NAND3_X1  g409(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT26), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(KEYINPUT26), .A2(G117), .A3(G2104), .A4(G2105), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  OAI211_X1 g414(.A(G141), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n464), .A2(G105), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n833), .B1(new_n834), .B2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G129), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n474), .B2(new_n475), .ZN(new_n846));
  NOR3_X1   g421(.A1(new_n846), .A2(KEYINPUT87), .A3(new_n842), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(G29), .ZN(new_n849));
  NOR2_X1   g424(.A1(G29), .A2(G32), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(KEYINPUT88), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(KEYINPUT88), .B2(new_n849), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT27), .B(G1996), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n853), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n851), .B(new_n855), .C1(KEYINPUT88), .C2(new_n849), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n754), .A2(G2090), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n700), .A2(G20), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT23), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n573), .B2(new_n700), .ZN(new_n860));
  INV_X1    g435(.A(G1956), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  AND4_X1   g437(.A1(new_n755), .A2(new_n832), .A3(new_n857), .A4(new_n862), .ZN(new_n863));
  AND2_X1   g438(.A1(new_n749), .A2(new_n863), .ZN(G311));
  AND3_X1   g439(.A1(new_n749), .A2(KEYINPUT91), .A3(new_n863), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT91), .B1(new_n749), .B2(new_n863), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(G150));
  NAND2_X1  g442(.A1(new_n511), .A2(G55), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n514), .A2(G93), .A3(new_n528), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n513), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT37), .Z(new_n873));
  NAND2_X1  g448(.A1(new_n607), .A2(G559), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n514), .A2(G67), .ZN(new_n876));
  NAND2_X1  g451(.A1(G80), .A2(G543), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n513), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n869), .A2(new_n868), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI22_X1  g455(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n543), .B(new_n542), .C1(new_n881), .C2(new_n513), .ZN(new_n882));
  OAI21_X1  g457(.A(KEYINPUT92), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n545), .A2(new_n884), .A3(new_n871), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(KEYINPUT93), .B1(new_n545), .B2(new_n871), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT93), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n880), .A2(new_n888), .A3(new_n882), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  OR2_X1    g466(.A1(new_n875), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n875), .A2(new_n891), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT94), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n894), .ZN(new_n897));
  AOI21_X1  g472(.A(G860), .B1(new_n897), .B2(KEYINPUT39), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(KEYINPUT95), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(KEYINPUT95), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n873), .B1(new_n900), .B2(new_n901), .ZN(G145));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT101), .B(G37), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n733), .A2(new_n738), .ZN(new_n908));
  OAI21_X1  g483(.A(G130), .B1(new_n811), .B2(new_n812), .ZN(new_n909));
  INV_X1    g484(.A(new_n631), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n459), .A2(G118), .ZN(new_n911));
  OAI21_X1  g486(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n913), .B1(new_n482), .B2(G142), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(G130), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(new_n474), .B2(new_n475), .ZN(new_n917));
  INV_X1    g492(.A(G142), .ZN(new_n918));
  OAI22_X1  g493(.A1(new_n622), .A2(new_n918), .B1(new_n911), .B2(new_n912), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n631), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n908), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n908), .B1(new_n915), .B2(new_n920), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n907), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g498(.A1(new_n917), .A2(new_n919), .A3(new_n631), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n910), .B1(new_n909), .B2(new_n914), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n739), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n908), .A2(new_n915), .A3(new_n920), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n906), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n923), .A2(KEYINPUT100), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n923), .A2(new_n928), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT100), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n823), .B1(new_n844), .B2(new_n847), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT96), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n500), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n492), .A2(new_n496), .A3(KEYINPUT96), .A4(new_n499), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n834), .A2(new_n833), .A3(new_n843), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT87), .B1(new_n846), .B2(new_n842), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n821), .B1(new_n476), .B2(G128), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n818), .A4(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n933), .A2(new_n937), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n937), .B1(new_n933), .B2(new_n941), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT97), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n788), .A2(new_n792), .A3(new_n944), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n782), .A2(new_n787), .ZN(new_n947));
  OAI21_X1  g522(.A(KEYINPUT97), .B1(new_n947), .B2(new_n791), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n937), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n844), .A2(new_n847), .A3(new_n823), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n938), .A2(new_n939), .B1(new_n818), .B2(new_n940), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n933), .A2(new_n941), .A3(new_n937), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n929), .B(new_n932), .C1(new_n946), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n945), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n945), .A2(new_n948), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(new_n942), .B2(new_n943), .ZN(new_n960));
  AND3_X1   g535(.A1(new_n923), .A2(KEYINPUT100), .A3(new_n928), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT100), .B1(new_n923), .B2(new_n928), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n958), .B(new_n960), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n956), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n627), .B(G160), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(new_n484), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n905), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n960), .A2(new_n930), .A3(new_n958), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT102), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n960), .A2(new_n958), .A3(new_n970), .A4(new_n930), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n961), .A2(new_n962), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n960), .A2(new_n958), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n967), .A2(KEYINPUT103), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT103), .B1(new_n967), .B2(new_n976), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n903), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(new_n976), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n967), .A2(new_n976), .A3(KEYINPUT103), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT40), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g559(.A1(new_n979), .A2(new_n984), .ZN(G395));
  NAND2_X1  g560(.A1(new_n616), .A2(KEYINPUT104), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n607), .A2(new_n987), .A3(new_n614), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n891), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n883), .A2(new_n885), .B1(new_n887), .B2(new_n889), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n991), .A2(new_n986), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n607), .A2(new_n568), .A3(new_n572), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n605), .A2(new_n606), .ZN(new_n995));
  INV_X1    g570(.A(new_n602), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n568), .A2(new_n572), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT41), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n994), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n607), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n573), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n607), .A2(new_n568), .A3(new_n572), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT41), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT105), .B1(new_n993), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n998), .B1(new_n994), .B2(new_n997), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1001), .A2(KEYINPUT41), .A3(new_n1002), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1008), .A2(new_n1009), .A3(new_n990), .A4(new_n992), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n993), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1005), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT42), .ZN(new_n1014));
  AOI21_X1  g589(.A(G288), .B1(new_n518), .B2(new_n519), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n518), .A2(new_n519), .A3(G288), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G290), .A2(new_n712), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n596), .A2(G305), .A3(new_n597), .ZN(new_n1019));
  AOI22_X1  g594(.A1(new_n1016), .A2(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n1015), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1005), .A2(new_n1025), .A3(new_n1010), .A4(new_n1012), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1014), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1024), .B1(new_n1014), .B2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g603(.A(G868), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(G868), .B2(new_n880), .ZN(G295));
  OAI21_X1  g605(.A(new_n1029), .B1(G868), .B2(new_n880), .ZN(G331));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT43), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1024), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n581), .A2(G171), .A3(new_n1035), .A4(new_n582), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n581), .A2(G171), .A3(new_n582), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1037), .B(KEYINPUT106), .C1(new_n530), .C2(G171), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n891), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n581), .A2(G171), .A3(new_n582), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT106), .B1(G171), .B2(new_n530), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n991), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1039), .A2(new_n1011), .A3(new_n1043), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1039), .A2(new_n1043), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1034), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n991), .A2(new_n1042), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n991), .A2(new_n1042), .ZN(new_n1048));
  OAI22_X1  g623(.A1(new_n1047), .A2(new_n1048), .B1(new_n999), .B2(new_n1003), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1039), .A2(new_n1011), .A3(new_n1043), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n1024), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1046), .A2(new_n904), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1033), .B1(new_n1052), .B2(KEYINPUT109), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1046), .A2(new_n1051), .A3(new_n1054), .A4(new_n904), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1032), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1051), .ZN(new_n1057));
  INV_X1    g632(.A(G37), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1046), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1057), .B1(new_n1059), .B2(KEYINPUT107), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT107), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1046), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1060), .A2(KEYINPUT108), .A3(new_n1033), .A4(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1024), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT107), .B1(new_n1064), .B2(G37), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(new_n1062), .A3(new_n1033), .A4(new_n1051), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT108), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1056), .A2(new_n1063), .A3(new_n1068), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1065), .A2(new_n1062), .A3(KEYINPUT43), .A4(new_n1051), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1052), .A2(new_n1033), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1070), .A2(new_n1032), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(G397));
  INV_X1    g648(.A(G1384), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n500), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT110), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT45), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n500), .A2(new_n1078), .A3(new_n1074), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(G160), .A2(G40), .ZN(new_n1081));
  OR3_X1    g656(.A1(new_n1080), .A2(G1996), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT46), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  XOR2_X1   g659(.A(new_n1084), .B(KEYINPUT127), .Z(new_n1085));
  NOR2_X1   g660(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n823), .B(new_n826), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n848), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1082), .A2(new_n1083), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1085), .A2(KEYINPUT47), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n848), .B(G1996), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n1087), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n908), .A2(new_n742), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n739), .A2(new_n741), .ZN(new_n1094));
  NOR3_X1   g669(.A1(new_n1092), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1086), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1096), .A2(G1986), .A3(G290), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT48), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1092), .A2(new_n742), .A3(new_n908), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1100), .B1(new_n826), .B2(new_n824), .ZN(new_n1101));
  OAI22_X1  g676(.A1(new_n1097), .A2(new_n1099), .B1(new_n1101), .B2(new_n1096), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT47), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1090), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT111), .B(G1971), .Z(new_n1106));
  NAND3_X1  g681(.A1(new_n500), .A2(KEYINPUT45), .A3(new_n1074), .ZN(new_n1107));
  INV_X1    g682(.A(G40), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1108), .B(new_n466), .C1(G2105), .C2(new_n470), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(KEYINPUT45), .B1(new_n500), .B2(new_n1074), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1106), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1075), .A2(KEYINPUT50), .ZN(new_n1113));
  INV_X1    g688(.A(G2090), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT50), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n500), .A2(new_n1115), .A3(new_n1074), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1113), .A2(new_n1114), .A3(new_n1109), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1112), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G8), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n518), .A2(G8), .A3(new_n519), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT55), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n518), .A2(KEYINPUT55), .A3(G8), .A4(new_n519), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n509), .A2(G86), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n511), .A2(G48), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n593), .A2(new_n1127), .A3(new_n721), .A4(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT113), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT113), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n589), .A2(new_n1131), .A3(new_n593), .A4(new_n721), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(G305), .A2(G1981), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1133), .A2(KEYINPUT49), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT114), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT49), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1133), .A2(new_n1134), .A3(new_n1140), .A4(KEYINPUT49), .ZN(new_n1141));
  INV_X1    g716(.A(G8), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1075), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1142), .B1(new_n1143), .B2(new_n1109), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1136), .A2(new_n1139), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n706), .A2(G1976), .ZN(new_n1146));
  XNOR2_X1  g721(.A(KEYINPUT112), .B(G1976), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT52), .B1(G288), .B2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1146), .B(G8), .C1(new_n1075), .C2(new_n1081), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT52), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1124), .A2(new_n1118), .A3(G8), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1126), .A2(new_n1145), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1966), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1113), .A2(new_n768), .A3(new_n1109), .A4(new_n1116), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(G8), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1159), .A2(G286), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1105), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1124), .A2(new_n1118), .A3(G8), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1124), .B1(G8), .B2(new_n1118), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT63), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1159), .A2(new_n1165), .A3(G286), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n1167));
  AND3_X1   g742(.A1(new_n1145), .A2(new_n1152), .A3(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1167), .B1(new_n1145), .B2(new_n1152), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1164), .B(new_n1166), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1161), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1110), .ZN(new_n1172));
  INV_X1    g747(.A(G2078), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1172), .A2(KEYINPUT121), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1174), .A2(new_n1173), .A3(new_n1109), .A4(new_n1107), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT121), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1175), .A2(new_n1178), .A3(KEYINPUT53), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1113), .A2(new_n1109), .A3(new_n1116), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1180), .A2(new_n1176), .B1(new_n1181), .B2(new_n758), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(G171), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1154), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT51), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1186), .B(G8), .C1(new_n1158), .C2(new_n530), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n530), .A2(G8), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1188), .B1(new_n1158), .B2(new_n1190), .ZN(new_n1191));
  AOI211_X1 g766(.A(KEYINPUT120), .B(new_n1189), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1187), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI211_X1 g768(.A(new_n1186), .B(new_n1190), .C1(new_n1158), .C2(G8), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1189), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1196));
  XNOR2_X1  g771(.A(new_n1196), .B(new_n1188), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1159), .A2(KEYINPUT51), .A3(new_n1189), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1187), .ZN(new_n1200));
  NAND3_X1  g775(.A1(new_n1185), .A2(new_n1195), .A3(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1144), .ZN(new_n1202));
  INV_X1    g777(.A(G1976), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1145), .A2(new_n1203), .A3(new_n706), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n1204), .B2(new_n1133), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(KEYINPUT115), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1145), .A2(new_n1152), .A3(new_n1167), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n1205), .B1(new_n1209), .B2(new_n1162), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1171), .A2(new_n1201), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT54), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n462), .A2(KEYINPUT122), .A3(new_n465), .ZN(new_n1213));
  OR2_X1    g788(.A1(new_n1173), .A2(KEYINPUT124), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1173), .A2(KEYINPUT124), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1214), .A2(KEYINPUT53), .A3(G40), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1216), .B1(new_n466), .B2(new_n1217), .ZN(new_n1218));
  AOI22_X1  g793(.A1(new_n621), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1219));
  OAI21_X1  g794(.A(G2105), .B1(new_n1219), .B2(KEYINPUT123), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT123), .ZN(new_n1221));
  NOR2_X1   g796(.A1(new_n470), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g797(.A(new_n1213), .B(new_n1218), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1223), .B1(new_n1143), .B2(KEYINPUT45), .ZN(new_n1224));
  AND3_X1   g799(.A1(new_n1080), .A2(new_n1224), .A3(KEYINPUT125), .ZN(new_n1225));
  AOI21_X1  g800(.A(KEYINPUT125), .B1(new_n1080), .B2(new_n1224), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1181), .A2(new_n758), .ZN(new_n1229));
  NAND3_X1  g804(.A1(new_n1228), .A2(G301), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g806(.A(G301), .B1(new_n1179), .B2(new_n1182), .ZN(new_n1232));
  OAI21_X1  g807(.A(new_n1212), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1182), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1234), .A2(G171), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1179), .A2(G301), .A3(new_n1182), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1235), .A2(KEYINPUT54), .A3(new_n1236), .ZN(new_n1237));
  NOR3_X1   g812(.A1(new_n1206), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1238));
  OAI211_X1 g813(.A(new_n1199), .B(new_n1187), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1239));
  NAND4_X1  g814(.A1(new_n1233), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  OR2_X1    g815(.A1(new_n1240), .A2(KEYINPUT126), .ZN(new_n1241));
  NOR2_X1   g816(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1242));
  AOI22_X1  g817(.A1(new_n1181), .A2(new_n798), .B1(new_n826), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1243), .A2(KEYINPUT60), .ZN(new_n1244));
  NOR2_X1   g819(.A1(new_n1244), .A2(new_n607), .ZN(new_n1245));
  XOR2_X1   g820(.A(KEYINPUT58), .B(G1341), .Z(new_n1246));
  OAI21_X1  g821(.A(new_n1246), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1247));
  NAND3_X1  g822(.A1(new_n1174), .A2(new_n1109), .A3(new_n1107), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1247), .B1(new_n1248), .B2(G1996), .ZN(new_n1249));
  AOI21_X1  g824(.A(KEYINPUT59), .B1(new_n1249), .B2(new_n545), .ZN(new_n1250));
  AND3_X1   g825(.A1(new_n1249), .A2(KEYINPUT59), .A3(new_n545), .ZN(new_n1251));
  NOR3_X1   g826(.A1(new_n1245), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  OR2_X1    g827(.A1(new_n1243), .A2(KEYINPUT60), .ZN(new_n1253));
  NAND3_X1  g828(.A1(new_n1253), .A2(new_n607), .A3(new_n1244), .ZN(new_n1254));
  NAND3_X1  g829(.A1(new_n569), .A2(new_n571), .A3(new_n556), .ZN(new_n1255));
  NOR2_X1   g830(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1256));
  NAND2_X1  g831(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1257));
  XOR2_X1   g832(.A(new_n1257), .B(KEYINPUT118), .Z(new_n1258));
  INV_X1    g833(.A(new_n1258), .ZN(new_n1259));
  OR3_X1    g834(.A1(new_n1255), .A2(new_n1256), .A3(new_n1259), .ZN(new_n1260));
  OAI21_X1  g835(.A(new_n1259), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1261));
  NAND2_X1  g836(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1262), .A2(KEYINPUT119), .ZN(new_n1263));
  XNOR2_X1  g838(.A(KEYINPUT56), .B(G2072), .ZN(new_n1264));
  NAND3_X1  g839(.A1(new_n1172), .A2(new_n1174), .A3(new_n1264), .ZN(new_n1265));
  NAND2_X1  g840(.A1(new_n1181), .A2(new_n861), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g842(.A(KEYINPUT119), .ZN(new_n1268));
  NAND3_X1  g843(.A1(new_n1260), .A2(new_n1268), .A3(new_n1261), .ZN(new_n1269));
  NAND3_X1  g844(.A1(new_n1263), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g845(.A1(new_n1262), .A2(new_n1265), .A3(new_n1266), .ZN(new_n1271));
  NAND3_X1  g846(.A1(new_n1270), .A2(KEYINPUT61), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g847(.A(KEYINPUT61), .ZN(new_n1273));
  INV_X1    g848(.A(new_n1271), .ZN(new_n1274));
  AOI21_X1  g849(.A(new_n1262), .B1(new_n1266), .B2(new_n1265), .ZN(new_n1275));
  OAI21_X1  g850(.A(new_n1273), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND4_X1  g851(.A1(new_n1252), .A2(new_n1254), .A3(new_n1272), .A4(new_n1276), .ZN(new_n1277));
  INV_X1    g852(.A(new_n1270), .ZN(new_n1278));
  NOR2_X1   g853(.A1(new_n1243), .A2(new_n1000), .ZN(new_n1279));
  AOI21_X1  g854(.A(new_n1278), .B1(new_n1271), .B2(new_n1279), .ZN(new_n1280));
  AOI22_X1  g855(.A1(new_n1240), .A2(KEYINPUT126), .B1(new_n1277), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g856(.A(new_n1211), .B1(new_n1241), .B2(new_n1281), .ZN(new_n1282));
  XOR2_X1   g857(.A(G290), .B(G1986), .Z(new_n1283));
  AOI21_X1  g858(.A(new_n1096), .B1(new_n1095), .B2(new_n1283), .ZN(new_n1284));
  OAI21_X1  g859(.A(new_n1104), .B1(new_n1282), .B2(new_n1284), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g860(.A1(new_n982), .A2(new_n983), .ZN(new_n1287));
  AND2_X1   g861(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1288));
  OAI211_X1 g862(.A(G319), .B(new_n654), .C1(new_n672), .C2(new_n673), .ZN(new_n1289));
  AOI21_X1  g863(.A(new_n1289), .B1(new_n696), .B2(new_n698), .ZN(new_n1290));
  AND3_X1   g864(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(G308));
  NAND3_X1  g865(.A1(new_n1287), .A2(new_n1288), .A3(new_n1290), .ZN(G225));
endmodule


