

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744;

  NOR2_X1 U371 ( .A1(n672), .A2(n580), .ZN(n581) );
  INV_X1 U372 ( .A(G953), .ZN(n730) );
  XNOR2_X2 U373 ( .A(n472), .B(n471), .ZN(n541) );
  NOR2_X2 U374 ( .A1(G902), .A2(n619), .ZN(n472) );
  OR2_X1 U375 ( .A1(n721), .A2(n616), .ZN(n652) );
  OR2_X1 U376 ( .A1(n567), .A2(n663), .ZN(n392) );
  NOR2_X1 U377 ( .A1(n743), .A2(n744), .ZN(n602) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n426) );
  NAND2_X1 U379 ( .A1(n608), .A2(n649), .ZN(n729) );
  XNOR2_X1 U380 ( .A(n596), .B(KEYINPUT40), .ZN(n743) );
  NOR2_X1 U381 ( .A1(n681), .A2(n686), .ZN(n358) );
  NOR2_X1 U382 ( .A1(n525), .A2(n524), .ZN(n597) );
  XNOR2_X1 U383 ( .A(n515), .B(n514), .ZN(n557) );
  INV_X1 U384 ( .A(KEYINPUT30), .ZN(n369) );
  NAND2_X1 U385 ( .A1(n386), .A2(n385), .ZN(n608) );
  NOR2_X1 U386 ( .A1(n391), .A2(n605), .ZN(n389) );
  NAND2_X1 U387 ( .A1(n603), .A2(n392), .ZN(n391) );
  NOR2_X1 U388 ( .A1(n517), .A2(n362), .ZN(n535) );
  NOR2_X1 U389 ( .A1(n690), .A2(n371), .ZN(n539) );
  NOR2_X1 U390 ( .A1(n606), .A2(n595), .ZN(n596) );
  BUF_X1 U391 ( .A(n538), .Z(n371) );
  XNOR2_X1 U392 ( .A(n373), .B(n372), .ZN(n690) );
  XNOR2_X1 U393 ( .A(n358), .B(n598), .ZN(n679) );
  XNOR2_X1 U394 ( .A(n370), .B(n369), .ZN(n572) );
  BUF_X1 U395 ( .A(n557), .Z(n516) );
  XNOR2_X1 U396 ( .A(n481), .B(n431), .ZN(n727) );
  XNOR2_X1 U397 ( .A(n363), .B(G125), .ZN(n460) );
  INV_X2 U398 ( .A(G143), .ZN(n374) );
  XNOR2_X1 U399 ( .A(KEYINPUT4), .B(KEYINPUT64), .ZN(n430) );
  INV_X1 U400 ( .A(G146), .ZN(n363) );
  XNOR2_X2 U401 ( .A(n526), .B(KEYINPUT70), .ZN(n529) );
  NOR2_X2 U402 ( .A1(n557), .A2(n666), .ZN(n526) );
  XNOR2_X1 U403 ( .A(n435), .B(n434), .ZN(n570) );
  XNOR2_X1 U404 ( .A(n459), .B(n458), .ZN(n538) );
  XNOR2_X1 U405 ( .A(n497), .B(n496), .ZN(n582) );
  XNOR2_X1 U406 ( .A(n727), .B(G146), .ZN(n495) );
  OR2_X1 U407 ( .A1(n729), .A2(n615), .ZN(n616) );
  NAND2_X1 U408 ( .A1(n412), .A2(n449), .ZN(n406) );
  NAND2_X1 U409 ( .A1(KEYINPUT68), .A2(KEYINPUT19), .ZN(n407) );
  NAND2_X1 U410 ( .A1(n410), .A2(n409), .ZN(n408) );
  NAND2_X1 U411 ( .A1(n412), .A2(KEYINPUT19), .ZN(n409) );
  NAND2_X1 U412 ( .A1(KEYINPUT68), .A2(n449), .ZN(n410) );
  XNOR2_X1 U413 ( .A(n381), .B(KEYINPUT105), .ZN(n380) );
  NAND2_X1 U414 ( .A1(n533), .A2(n680), .ZN(n382) );
  XNOR2_X1 U415 ( .A(G113), .B(G143), .ZN(n465) );
  XOR2_X1 U416 ( .A(G104), .B(G122), .Z(n466) );
  NAND2_X1 U417 ( .A1(n575), .A2(n683), .ZN(n448) );
  XNOR2_X1 U418 ( .A(n549), .B(KEYINPUT45), .ZN(n413) );
  XNOR2_X1 U419 ( .A(n582), .B(n498), .ZN(n663) );
  INV_X1 U420 ( .A(KEYINPUT33), .ZN(n372) );
  XNOR2_X1 U421 ( .A(n488), .B(n354), .ZN(n517) );
  NOR2_X1 U422 ( .A1(n538), .A2(n487), .ZN(n488) );
  BUF_X1 U423 ( .A(n563), .Z(n362) );
  XNOR2_X1 U424 ( .A(n448), .B(n412), .ZN(n411) );
  NAND2_X1 U425 ( .A1(n529), .A2(n582), .ZN(n574) );
  NAND2_X1 U426 ( .A1(n378), .A2(n376), .ZN(n375) );
  NOR2_X1 U427 ( .A1(n377), .A2(n714), .ZN(n376) );
  NAND2_X1 U428 ( .A1(n710), .A2(n356), .ZN(n378) );
  NOR2_X1 U429 ( .A1(n355), .A2(G472), .ZN(n377) );
  XNOR2_X1 U430 ( .A(G101), .B(G107), .ZN(n493) );
  XNOR2_X1 U431 ( .A(n661), .B(n660), .ZN(n420) );
  INV_X1 U432 ( .A(KEYINPUT85), .ZN(n660) );
  NAND2_X1 U433 ( .A1(n407), .A2(n406), .ZN(n405) );
  XNOR2_X1 U434 ( .A(n394), .B(n393), .ZN(n424) );
  XNOR2_X1 U435 ( .A(G116), .B(G131), .ZN(n393) );
  XNOR2_X1 U436 ( .A(n395), .B(KEYINPUT95), .ZN(n394) );
  XNOR2_X1 U437 ( .A(KEYINPUT5), .B(KEYINPUT77), .ZN(n395) );
  OR2_X1 U438 ( .A1(n604), .A2(KEYINPUT48), .ZN(n388) );
  XNOR2_X1 U439 ( .A(n364), .B(n425), .ZN(n438) );
  XNOR2_X1 U440 ( .A(n361), .B(KEYINPUT90), .ZN(n364) );
  XNOR2_X1 U441 ( .A(G119), .B(KEYINPUT3), .ZN(n361) );
  XOR2_X1 U442 ( .A(G902), .B(KEYINPUT15), .Z(n611) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n450) );
  XNOR2_X1 U444 ( .A(n591), .B(KEYINPUT38), .ZN(n684) );
  INV_X1 U445 ( .A(KEYINPUT76), .ZN(n530) );
  OR2_X1 U446 ( .A1(G237), .A2(G902), .ZN(n447) );
  NAND2_X1 U447 ( .A1(n570), .A2(n683), .ZN(n370) );
  XNOR2_X1 U448 ( .A(n360), .B(KEYINPUT6), .ZN(n559) );
  XNOR2_X1 U449 ( .A(G140), .B(KEYINPUT23), .ZN(n502) );
  XNOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT93), .ZN(n507) );
  XNOR2_X1 U451 ( .A(KEYINPUT8), .B(KEYINPUT71), .ZN(n477) );
  XNOR2_X1 U452 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n473) );
  XOR2_X1 U453 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n474) );
  XNOR2_X1 U454 ( .A(n467), .B(n421), .ZN(n468) );
  XNOR2_X1 U455 ( .A(n489), .B(n417), .ZN(n491) );
  NAND2_X1 U456 ( .A1(n721), .A2(n656), .ZN(n657) );
  XNOR2_X1 U457 ( .A(n594), .B(n593), .ZN(n606) );
  XNOR2_X1 U458 ( .A(KEYINPUT88), .B(KEYINPUT39), .ZN(n593) );
  AND2_X1 U459 ( .A1(n592), .A2(n684), .ZN(n594) );
  INV_X1 U460 ( .A(n559), .ZN(n550) );
  XNOR2_X1 U461 ( .A(n367), .B(n366), .ZN(n567) );
  INV_X1 U462 ( .A(KEYINPUT36), .ZN(n366) );
  NOR2_X1 U463 ( .A1(n566), .A2(n591), .ZN(n367) );
  NOR2_X1 U464 ( .A1(n577), .A2(n576), .ZN(n635) );
  NOR2_X1 U465 ( .A1(n584), .A2(n599), .ZN(n637) );
  NAND2_X1 U466 ( .A1(n411), .A2(n449), .ZN(n579) );
  OR2_X1 U467 ( .A1(n411), .A2(n449), .ZN(n578) );
  NAND2_X1 U468 ( .A1(n416), .A2(n353), .ZN(n415) );
  INV_X1 U469 ( .A(n574), .ZN(n569) );
  NOR2_X1 U470 ( .A1(n379), .A2(n375), .ZN(n618) );
  NOR2_X1 U471 ( .A1(n710), .A2(n355), .ZN(n379) );
  XNOR2_X1 U472 ( .A(n709), .B(n708), .ZN(n400) );
  XNOR2_X1 U473 ( .A(n707), .B(n706), .ZN(n397) );
  NOR2_X1 U474 ( .A1(n714), .A2(n704), .ZN(n705) );
  XNOR2_X1 U475 ( .A(n419), .B(n418), .ZN(G75) );
  XNOR2_X1 U476 ( .A(KEYINPUT119), .B(KEYINPUT53), .ZN(n418) );
  NAND2_X1 U477 ( .A1(n420), .A2(n423), .ZN(n419) );
  XOR2_X1 U478 ( .A(n442), .B(n460), .Z(n350) );
  AND2_X1 U479 ( .A1(n390), .A2(n604), .ZN(n351) );
  AND2_X1 U480 ( .A1(G210), .A2(n447), .ZN(n352) );
  AND2_X1 U481 ( .A1(n672), .A2(n516), .ZN(n353) );
  XOR2_X1 U482 ( .A(KEYINPUT66), .B(KEYINPUT22), .Z(n354) );
  XOR2_X1 U483 ( .A(n433), .B(KEYINPUT62), .Z(n355) );
  NOR2_X1 U484 ( .A1(G952), .A2(n730), .ZN(n714) );
  AND2_X1 U485 ( .A1(n355), .A2(G472), .ZN(n356) );
  INV_X1 U486 ( .A(KEYINPUT48), .ZN(n605) );
  XNOR2_X1 U487 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n357) );
  XNOR2_X1 U488 ( .A(n439), .B(n438), .ZN(n716) );
  XNOR2_X1 U489 ( .A(n359), .B(n350), .ZN(n445) );
  XNOR2_X1 U490 ( .A(n443), .B(n444), .ZN(n359) );
  BUF_X1 U491 ( .A(n570), .Z(n360) );
  XNOR2_X1 U492 ( .A(n417), .B(KEYINPUT16), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n368), .B(n508), .ZN(n509) );
  NAND2_X1 U494 ( .A1(n547), .A2(n548), .ZN(n414) );
  NOR2_X2 U495 ( .A1(n544), .A2(n522), .ZN(n523) );
  NAND2_X1 U496 ( .A1(n391), .A2(n605), .ZN(n365) );
  XNOR2_X2 U497 ( .A(n446), .B(n352), .ZN(n575) );
  NOR2_X1 U498 ( .A1(n590), .A2(n589), .ZN(n604) );
  NAND2_X1 U499 ( .A1(n365), .A2(n388), .ZN(n387) );
  XNOR2_X1 U500 ( .A(n428), .B(n429), .ZN(n432) );
  XNOR2_X1 U501 ( .A(n506), .B(n507), .ZN(n368) );
  INV_X1 U502 ( .A(n529), .ZN(n662) );
  XNOR2_X1 U503 ( .A(n716), .B(n445), .ZN(n701) );
  NOR2_X2 U504 ( .A1(n740), .A2(n742), .ZN(n544) );
  NAND2_X1 U505 ( .A1(n537), .A2(n550), .ZN(n373) );
  XNOR2_X1 U506 ( .A(n531), .B(n530), .ZN(n537) );
  XNOR2_X2 U507 ( .A(n441), .B(G134), .ZN(n481) );
  XNOR2_X2 U508 ( .A(n374), .B(G128), .ZN(n441) );
  AND2_X4 U509 ( .A1(n700), .A2(n652), .ZN(n710) );
  AND2_X1 U510 ( .A1(n383), .A2(n380), .ZN(n546) );
  NAND2_X1 U511 ( .A1(n382), .A2(n741), .ZN(n381) );
  NAND2_X1 U512 ( .A1(n739), .A2(KEYINPUT44), .ZN(n383) );
  XNOR2_X2 U513 ( .A(n384), .B(KEYINPUT35), .ZN(n739) );
  NAND2_X1 U514 ( .A1(n542), .A2(n568), .ZN(n384) );
  INV_X1 U515 ( .A(n650), .ZN(n390) );
  NAND2_X1 U516 ( .A1(n387), .A2(n390), .ZN(n385) );
  NAND2_X1 U517 ( .A1(n389), .A2(n351), .ZN(n386) );
  INV_X1 U518 ( .A(n392), .ZN(n647) );
  NOR2_X1 U519 ( .A1(n396), .A2(n714), .ZN(G54) );
  XNOR2_X1 U520 ( .A(n398), .B(n397), .ZN(n396) );
  NAND2_X1 U521 ( .A1(n710), .A2(G469), .ZN(n398) );
  NOR2_X1 U522 ( .A1(n399), .A2(n714), .ZN(G63) );
  XNOR2_X1 U523 ( .A(n401), .B(n400), .ZN(n399) );
  NAND2_X1 U524 ( .A1(n710), .A2(G478), .ZN(n401) );
  NAND2_X2 U525 ( .A1(n614), .A2(n613), .ZN(n700) );
  XNOR2_X1 U526 ( .A(n424), .B(KEYINPUT94), .ZN(n429) );
  NAND2_X1 U527 ( .A1(n403), .A2(n402), .ZN(n457) );
  NAND2_X1 U528 ( .A1(n448), .A2(n405), .ZN(n402) );
  NAND2_X1 U529 ( .A1(n404), .A2(n408), .ZN(n403) );
  INV_X1 U530 ( .A(n448), .ZN(n404) );
  INV_X1 U531 ( .A(KEYINPUT68), .ZN(n412) );
  XNOR2_X2 U532 ( .A(n414), .B(n413), .ZN(n721) );
  XNOR2_X2 U533 ( .A(n415), .B(KEYINPUT107), .ZN(n740) );
  XNOR2_X1 U534 ( .A(n535), .B(KEYINPUT106), .ZN(n416) );
  XNOR2_X2 U535 ( .A(G104), .B(G110), .ZN(n417) );
  XNOR2_X1 U536 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U537 ( .A(n701), .B(n357), .ZN(n702) );
  XOR2_X1 U538 ( .A(n466), .B(n465), .Z(n421) );
  XOR2_X1 U539 ( .A(n621), .B(n620), .Z(n422) );
  AND2_X1 U540 ( .A1(n698), .A2(n697), .ZN(n423) );
  XNOR2_X1 U541 ( .A(n438), .B(n427), .ZN(n428) );
  XNOR2_X1 U542 ( .A(n469), .B(n468), .ZN(n619) );
  XNOR2_X1 U543 ( .A(n432), .B(n495), .ZN(n433) );
  INV_X1 U544 ( .A(KEYINPUT1), .ZN(n498) );
  XNOR2_X1 U545 ( .A(n470), .B(G475), .ZN(n471) );
  INV_X1 U546 ( .A(KEYINPUT63), .ZN(n617) );
  XNOR2_X1 U547 ( .A(G101), .B(G113), .ZN(n425) );
  XOR2_X1 U548 ( .A(KEYINPUT79), .B(n426), .Z(n464) );
  NAND2_X1 U549 ( .A1(n464), .A2(G210), .ZN(n427) );
  INV_X1 U550 ( .A(n430), .ZN(n440) );
  XNOR2_X1 U551 ( .A(G137), .B(n440), .ZN(n431) );
  NOR2_X1 U552 ( .A1(G902), .A2(n433), .ZN(n435) );
  INV_X1 U553 ( .A(G472), .ZN(n434) );
  INV_X1 U554 ( .A(n570), .ZN(n672) );
  XNOR2_X1 U555 ( .A(G116), .B(G122), .ZN(n436) );
  XNOR2_X1 U556 ( .A(n436), .B(G107), .ZN(n476) );
  XNOR2_X1 U557 ( .A(n437), .B(n476), .ZN(n439) );
  XNOR2_X1 U558 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U559 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n442) );
  NAND2_X1 U560 ( .A1(G224), .A2(n730), .ZN(n444) );
  INV_X1 U561 ( .A(n611), .ZN(n484) );
  NAND2_X1 U562 ( .A1(n701), .A2(n484), .ZN(n446) );
  NAND2_X1 U563 ( .A1(G214), .A2(n447), .ZN(n683) );
  INV_X1 U564 ( .A(KEYINPUT19), .ZN(n449) );
  NOR2_X1 U565 ( .A1(G898), .A2(n730), .ZN(n715) );
  XNOR2_X1 U566 ( .A(n450), .B(KEYINPUT14), .ZN(n451) );
  XOR2_X1 U567 ( .A(KEYINPUT75), .B(n451), .Z(n453) );
  NAND2_X1 U568 ( .A1(G902), .A2(n453), .ZN(n551) );
  INV_X1 U569 ( .A(n551), .ZN(n452) );
  NAND2_X1 U570 ( .A1(n715), .A2(n452), .ZN(n455) );
  NAND2_X1 U571 ( .A1(G952), .A2(n453), .ZN(n695) );
  NOR2_X1 U572 ( .A1(G953), .A2(n695), .ZN(n454) );
  XNOR2_X1 U573 ( .A(KEYINPUT91), .B(n454), .ZN(n554) );
  NAND2_X1 U574 ( .A1(n455), .A2(n554), .ZN(n456) );
  NAND2_X1 U575 ( .A1(n457), .A2(n456), .ZN(n459) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(KEYINPUT69), .Z(n458) );
  XOR2_X1 U577 ( .A(G131), .B(G140), .Z(n489) );
  XNOR2_X1 U578 ( .A(n460), .B(KEYINPUT10), .ZN(n506) );
  XNOR2_X1 U579 ( .A(n489), .B(n506), .ZN(n726) );
  XOR2_X1 U580 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n462) );
  XNOR2_X1 U581 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n461) );
  XNOR2_X1 U582 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U583 ( .A(n726), .B(n463), .Z(n469) );
  NAND2_X1 U584 ( .A1(G214), .A2(n464), .ZN(n467) );
  XNOR2_X1 U585 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n470) );
  INV_X1 U586 ( .A(n541), .ZN(n525) );
  XNOR2_X1 U587 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U588 ( .A(n476), .B(n475), .Z(n480) );
  NAND2_X1 U589 ( .A1(n730), .A2(G234), .ZN(n478) );
  XNOR2_X1 U590 ( .A(n478), .B(n477), .ZN(n499) );
  NAND2_X1 U591 ( .A1(G217), .A2(n499), .ZN(n479) );
  XNOR2_X1 U592 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U593 ( .A(n482), .B(n481), .ZN(n709) );
  NOR2_X1 U594 ( .A1(n709), .A2(G902), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n483), .B(G478), .ZN(n540) );
  INV_X1 U596 ( .A(n540), .ZN(n524) );
  NAND2_X1 U597 ( .A1(n484), .A2(G234), .ZN(n485) );
  XNOR2_X1 U598 ( .A(n485), .B(KEYINPUT20), .ZN(n511) );
  NAND2_X1 U599 ( .A1(n511), .A2(G221), .ZN(n486) );
  XNOR2_X1 U600 ( .A(KEYINPUT21), .B(n486), .ZN(n666) );
  INV_X1 U601 ( .A(n666), .ZN(n555) );
  NAND2_X1 U602 ( .A1(n597), .A2(n555), .ZN(n487) );
  NAND2_X1 U603 ( .A1(G227), .A2(n730), .ZN(n490) );
  XNOR2_X1 U604 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n495), .B(n494), .ZN(n707) );
  NOR2_X1 U607 ( .A1(G902), .A2(n707), .ZN(n497) );
  XNOR2_X1 U608 ( .A(KEYINPUT73), .B(G469), .ZN(n496) );
  INV_X1 U609 ( .A(n663), .ZN(n563) );
  NAND2_X1 U610 ( .A1(n499), .A2(G221), .ZN(n510) );
  XOR2_X1 U611 ( .A(G110), .B(G128), .Z(n501) );
  XNOR2_X1 U612 ( .A(G119), .B(G137), .ZN(n500) );
  XNOR2_X1 U613 ( .A(n501), .B(n500), .ZN(n505) );
  XOR2_X1 U614 ( .A(KEYINPUT92), .B(KEYINPUT74), .Z(n503) );
  XNOR2_X1 U615 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U616 ( .A(n505), .B(n504), .ZN(n508) );
  XNOR2_X1 U617 ( .A(n510), .B(n509), .ZN(n712) );
  NOR2_X1 U618 ( .A1(n712), .A2(G902), .ZN(n515) );
  XOR2_X1 U619 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n513) );
  NAND2_X1 U620 ( .A1(n511), .A2(G217), .ZN(n512) );
  XNOR2_X1 U621 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U622 ( .A(KEYINPUT103), .B(n516), .Z(n667) );
  INV_X1 U623 ( .A(n667), .ZN(n518) );
  NOR2_X1 U624 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U625 ( .A1(n519), .A2(n362), .ZN(n520) );
  NOR2_X1 U626 ( .A1(n520), .A2(n550), .ZN(n521) );
  XNOR2_X1 U627 ( .A(n521), .B(KEYINPUT32), .ZN(n742) );
  INV_X1 U628 ( .A(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U629 ( .A(n523), .B(KEYINPUT65), .ZN(n548) );
  NAND2_X1 U630 ( .A1(n524), .A2(n541), .ZN(n644) );
  XNOR2_X1 U631 ( .A(KEYINPUT102), .B(n644), .ZN(n607) );
  NAND2_X1 U632 ( .A1(n525), .A2(n540), .ZN(n595) );
  NAND2_X1 U633 ( .A1(n607), .A2(n595), .ZN(n680) );
  NOR2_X1 U634 ( .A1(n371), .A2(n360), .ZN(n527) );
  NAND2_X1 U635 ( .A1(n569), .A2(n527), .ZN(n528) );
  XNOR2_X1 U636 ( .A(KEYINPUT96), .B(n528), .ZN(n626) );
  NAND2_X1 U637 ( .A1(n563), .A2(n529), .ZN(n531) );
  NAND2_X1 U638 ( .A1(n360), .A2(n537), .ZN(n675) );
  NOR2_X1 U639 ( .A1(n675), .A2(n371), .ZN(n532) );
  XNOR2_X1 U640 ( .A(n532), .B(KEYINPUT31), .ZN(n643) );
  NAND2_X1 U641 ( .A1(n626), .A2(n643), .ZN(n533) );
  NOR2_X1 U642 ( .A1(n667), .A2(n550), .ZN(n534) );
  NAND2_X1 U643 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U644 ( .A(KEYINPUT104), .B(n536), .ZN(n741) );
  XNOR2_X1 U645 ( .A(n539), .B(KEYINPUT34), .ZN(n542) );
  NOR2_X1 U646 ( .A1(n541), .A2(n540), .ZN(n568) );
  NOR2_X1 U647 ( .A1(n739), .A2(KEYINPUT44), .ZN(n543) );
  NAND2_X1 U648 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X1 U649 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U650 ( .A(KEYINPUT86), .ZN(n549) );
  XNOR2_X1 U651 ( .A(KEYINPUT108), .B(n595), .ZN(n640) );
  NOR2_X1 U652 ( .A1(G900), .A2(n551), .ZN(n552) );
  NAND2_X1 U653 ( .A1(G953), .A2(n552), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n571) );
  NAND2_X1 U655 ( .A1(n555), .A2(n571), .ZN(n556) );
  XOR2_X1 U656 ( .A(KEYINPUT72), .B(n556), .Z(n558) );
  NAND2_X1 U657 ( .A1(n558), .A2(n557), .ZN(n580) );
  NOR2_X1 U658 ( .A1(n559), .A2(n580), .ZN(n560) );
  XNOR2_X1 U659 ( .A(n560), .B(KEYINPUT109), .ZN(n561) );
  NOR2_X1 U660 ( .A1(n640), .A2(n561), .ZN(n562) );
  NAND2_X1 U661 ( .A1(n562), .A2(n683), .ZN(n566) );
  NOR2_X1 U662 ( .A1(n362), .A2(n566), .ZN(n564) );
  XNOR2_X1 U663 ( .A(n564), .B(KEYINPUT43), .ZN(n565) );
  NOR2_X1 U664 ( .A1(n575), .A2(n565), .ZN(n650) );
  INV_X1 U665 ( .A(n575), .ZN(n591) );
  INV_X1 U666 ( .A(n568), .ZN(n577) );
  NAND2_X1 U667 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X2 U668 ( .A1(n574), .A2(n573), .ZN(n592) );
  NAND2_X1 U669 ( .A1(n575), .A2(n592), .ZN(n576) );
  XNOR2_X1 U670 ( .A(n635), .B(KEYINPUT83), .ZN(n586) );
  AND2_X1 U671 ( .A1(n579), .A2(n578), .ZN(n584) );
  XNOR2_X1 U672 ( .A(KEYINPUT28), .B(n581), .ZN(n583) );
  NAND2_X1 U673 ( .A1(n583), .A2(n582), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n637), .A2(n680), .ZN(n588) );
  NAND2_X1 U675 ( .A1(KEYINPUT47), .A2(n588), .ZN(n585) );
  NAND2_X1 U676 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U677 ( .A(n587), .B(KEYINPUT82), .ZN(n590) );
  NOR2_X1 U678 ( .A1(n588), .A2(KEYINPUT47), .ZN(n589) );
  INV_X1 U679 ( .A(n597), .ZN(n686) );
  NAND2_X1 U680 ( .A1(n684), .A2(n683), .ZN(n681) );
  XNOR2_X1 U681 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n598) );
  NOR2_X1 U682 ( .A1(n599), .A2(n679), .ZN(n600) );
  XNOR2_X1 U683 ( .A(n600), .B(KEYINPUT42), .ZN(n744) );
  XOR2_X1 U684 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n601) );
  XNOR2_X1 U685 ( .A(n602), .B(n601), .ZN(n603) );
  OR2_X1 U686 ( .A1(n607), .A2(n606), .ZN(n649) );
  XNOR2_X1 U687 ( .A(n729), .B(KEYINPUT78), .ZN(n609) );
  NOR2_X1 U688 ( .A1(n721), .A2(n609), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n610), .A2(n611), .ZN(n614) );
  NAND2_X1 U690 ( .A1(KEYINPUT2), .A2(n611), .ZN(n612) );
  XOR2_X1 U691 ( .A(n612), .B(KEYINPUT67), .Z(n613) );
  INV_X1 U692 ( .A(KEYINPUT2), .ZN(n615) );
  XNOR2_X1 U693 ( .A(n618), .B(n617), .ZN(G57) );
  NAND2_X1 U694 ( .A1(n710), .A2(G475), .ZN(n622) );
  XOR2_X1 U695 ( .A(KEYINPUT89), .B(KEYINPUT120), .Z(n621) );
  XNOR2_X1 U696 ( .A(n619), .B(KEYINPUT59), .ZN(n620) );
  XNOR2_X1 U697 ( .A(n622), .B(n422), .ZN(n623) );
  NOR2_X2 U698 ( .A1(n623), .A2(n714), .ZN(n624) );
  XNOR2_X1 U699 ( .A(n624), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U700 ( .A1(n626), .A2(n640), .ZN(n625) );
  XOR2_X1 U701 ( .A(G104), .B(n625), .Z(G6) );
  NOR2_X1 U702 ( .A1(n644), .A2(n626), .ZN(n630) );
  XOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n628) );
  XNOR2_X1 U704 ( .A(G107), .B(KEYINPUT111), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n630), .B(n629), .ZN(G9) );
  XOR2_X1 U707 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n633) );
  INV_X1 U708 ( .A(n644), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n637), .A2(n631), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U711 ( .A(G128), .B(n634), .ZN(G30) );
  XOR2_X1 U712 ( .A(G143), .B(n635), .Z(G45) );
  XOR2_X1 U713 ( .A(G146), .B(KEYINPUT113), .Z(n639) );
  INV_X1 U714 ( .A(n640), .ZN(n636) );
  NAND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U716 ( .A(n639), .B(n638), .ZN(G48) );
  NOR2_X1 U717 ( .A1(n640), .A2(n643), .ZN(n641) );
  XOR2_X1 U718 ( .A(KEYINPUT114), .B(n641), .Z(n642) );
  XNOR2_X1 U719 ( .A(G113), .B(n642), .ZN(G15) );
  NOR2_X1 U720 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U721 ( .A(G116), .B(KEYINPUT115), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(G18) );
  XNOR2_X1 U723 ( .A(G125), .B(n647), .ZN(n648) );
  XNOR2_X1 U724 ( .A(n648), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U725 ( .A(G134), .B(n649), .ZN(G36) );
  XOR2_X1 U726 ( .A(G140), .B(n650), .Z(G42) );
  OR2_X1 U727 ( .A1(n615), .A2(KEYINPUT81), .ZN(n651) );
  NAND2_X1 U728 ( .A1(n729), .A2(n651), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U730 ( .A1(KEYINPUT81), .A2(n615), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n655), .A2(n654), .ZN(n659) );
  XNOR2_X1 U732 ( .A(KEYINPUT2), .B(KEYINPUT81), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(KEYINPUT84), .ZN(n658) );
  NAND2_X1 U734 ( .A1(n659), .A2(n658), .ZN(n661) );
  OR2_X1 U735 ( .A1(n690), .A2(n679), .ZN(n698) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(KEYINPUT50), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT117), .B(n665), .ZN(n671) );
  NAND2_X1 U739 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT116), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT49), .B(n669), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U744 ( .A(n674), .B(KEYINPUT118), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U746 ( .A(KEYINPUT51), .B(n677), .ZN(n678) );
  NOR2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n692) );
  INV_X1 U748 ( .A(n680), .ZN(n682) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n688) );
  NOR2_X1 U750 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U755 ( .A(n693), .B(KEYINPUT52), .ZN(n694) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U757 ( .A1(G953), .A2(n696), .ZN(n697) );
  AND2_X1 U758 ( .A1(n652), .A2(G210), .ZN(n699) );
  NAND2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n703) );
  XNOR2_X1 U760 ( .A(KEYINPUT56), .B(n705), .ZN(G51) );
  XOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n706) );
  XOR2_X1 U762 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n708) );
  NAND2_X1 U763 ( .A1(G217), .A2(n710), .ZN(n711) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  NOR2_X1 U765 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U766 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n725) );
  NAND2_X1 U769 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U770 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n720), .A2(G898), .ZN(n723) );
  OR2_X1 U772 ( .A1(n721), .A2(G953), .ZN(n722) );
  NAND2_X1 U773 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U774 ( .A(n725), .B(n724), .Z(G69) );
  XNOR2_X1 U775 ( .A(n726), .B(KEYINPUT125), .ZN(n728) );
  XNOR2_X1 U776 ( .A(n728), .B(n727), .ZN(n732) );
  XNOR2_X1 U777 ( .A(n732), .B(n729), .ZN(n731) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(n738) );
  XNOR2_X1 U779 ( .A(KEYINPUT126), .B(n732), .ZN(n733) );
  XNOR2_X1 U780 ( .A(G227), .B(n733), .ZN(n734) );
  NAND2_X1 U781 ( .A1(G900), .A2(n734), .ZN(n735) );
  XOR2_X1 U782 ( .A(KEYINPUT127), .B(n735), .Z(n736) );
  NAND2_X1 U783 ( .A1(G953), .A2(n736), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n738), .A2(n737), .ZN(G72) );
  XOR2_X1 U785 ( .A(n739), .B(G122), .Z(G24) );
  XOR2_X1 U786 ( .A(G110), .B(n740), .Z(G12) );
  XNOR2_X1 U787 ( .A(G101), .B(n741), .ZN(G3) );
  XOR2_X1 U788 ( .A(G119), .B(n742), .Z(G21) );
  XOR2_X1 U789 ( .A(n743), .B(G131), .Z(G33) );
  XOR2_X1 U790 ( .A(G137), .B(n744), .Z(G39) );
endmodule

