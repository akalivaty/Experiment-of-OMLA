//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT84), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  AND3_X1   g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n195));
  OAI21_X1  g009(.A(G107), .B1(new_n189), .B2(KEYINPUT3), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(KEYINPUT3), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT85), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT4), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT85), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(new_n196), .A4(new_n197), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n199), .A2(new_n200), .A3(G101), .A4(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT69), .B1(KEYINPUT2), .B2(G113), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR3_X1   g020(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n208));
  INV_X1    g022(.A(G113), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n206), .A2(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n211));
  XNOR2_X1  g025(.A(G116), .B(G119), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(KEYINPUT2), .A2(G113), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT69), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n208), .A3(new_n209), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n217), .B2(new_n205), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n211), .B1(new_n218), .B2(new_n212), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n204), .A2(new_n214), .A3(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n199), .A2(G101), .A3(new_n203), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n201), .A2(new_n224), .A3(new_n196), .A4(new_n197), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(KEYINPUT4), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n223), .A2(KEYINPUT86), .A3(new_n226), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n222), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(G104), .B1(new_n192), .B2(new_n194), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT87), .B1(new_n189), .B2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n191), .A3(G104), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n225), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT5), .ZN(new_n240));
  INV_X1    g054(.A(G119), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(G116), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT92), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n243), .B(G113), .C1(new_n240), .C2(new_n213), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n218), .A2(new_n212), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n239), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n188), .B1(new_n231), .B2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n204), .A2(new_n214), .A3(new_n221), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n223), .A2(KEYINPUT86), .A3(new_n226), .ZN(new_n250));
  AOI21_X1  g064(.A(KEYINPUT86), .B1(new_n223), .B2(new_n226), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n246), .A3(new_n187), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g073(.A1(KEYINPUT67), .A2(G128), .ZN(new_n260));
  NOR2_X1   g074(.A1(KEYINPUT67), .A2(G128), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT1), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n263), .B1(G143), .B2(new_n255), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n259), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n257), .B2(G146), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n255), .A2(KEYINPUT64), .A3(G143), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT1), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .A4(new_n258), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  OR2_X1    g089(.A1(KEYINPUT0), .A2(G128), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n259), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n275), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n267), .A2(new_n268), .A3(new_n278), .A4(new_n258), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G125), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G953), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G224), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT93), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n282), .B(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n288), .B(new_n188), .C1(new_n231), .C2(new_n247), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n254), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n187), .B(KEYINPUT8), .Z(new_n291));
  NAND2_X1  g105(.A1(new_n244), .A2(new_n245), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n238), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n291), .B1(new_n293), .B2(new_n246), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n286), .B(KEYINPUT94), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT7), .ZN(new_n296));
  INV_X1    g110(.A(new_n286), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n282), .B2(new_n297), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n274), .A2(new_n281), .B1(KEYINPUT7), .B2(new_n297), .ZN(new_n299));
  NOR3_X1   g113(.A1(new_n294), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(G902), .B1(new_n300), .B2(new_n253), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(KEYINPUT95), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n304), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n290), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(G952), .A3(new_n283), .ZN(new_n310));
  XNOR2_X1  g124(.A(KEYINPUT21), .B(G898), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(new_n314), .B(KEYINPUT102), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  INV_X1    g130(.A(G237), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n317), .A2(new_n283), .A3(G214), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n257), .ZN(new_n319));
  NOR2_X1   g133(.A1(G237), .A2(G953), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(G143), .A3(G214), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(KEYINPUT96), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT18), .ZN(new_n323));
  INV_X1    g137(.A(G131), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n319), .A2(KEYINPUT96), .A3(new_n326), .A4(new_n321), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n273), .A2(G140), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n255), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n330), .A2(new_n331), .ZN(new_n335));
  OR2_X1    g149(.A1(new_n335), .A2(new_n255), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n321), .ZN(new_n339));
  AOI21_X1  g153(.A(G143), .B1(new_n320), .B2(G214), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT17), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n319), .A2(new_n324), .A3(new_n321), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT78), .A4(KEYINPUT16), .ZN(new_n345));
  AND3_X1   g159(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n255), .B(new_n345), .C1(new_n346), .C2(new_n348), .ZN(new_n351));
  OAI211_X1 g165(.A(KEYINPUT17), .B(G131), .C1(new_n339), .C2(new_n340), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n344), .A2(new_n350), .A3(new_n351), .A4(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G113), .B(G122), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT98), .B(G104), .ZN(new_n355));
  OR2_X1    g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n355), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT99), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n356), .A2(new_n360), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AND3_X1   g176(.A1(new_n338), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n358), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n338), .B2(new_n353), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n316), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(G475), .ZN(new_n367));
  NOR2_X1   g181(.A1(G475), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n341), .A2(new_n343), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT19), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n330), .B(new_n331), .C1(KEYINPUT97), .C2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n371), .B(new_n255), .C1(new_n335), .C2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n350), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n364), .B1(new_n338), .B2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n368), .B1(new_n363), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT20), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n338), .A2(new_n374), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n358), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n338), .A2(new_n353), .A3(new_n362), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n378), .B1(new_n382), .B2(new_n368), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n315), .B(new_n367), .C1(new_n377), .C2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT100), .ZN(new_n385));
  INV_X1    g199(.A(G116), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n385), .B1(new_n386), .B2(G122), .ZN(new_n387));
  INV_X1    g201(.A(G122), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT100), .A3(G116), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(G122), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n192), .A2(new_n194), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(KEYINPUT14), .ZN(new_n396));
  OR3_X1    g210(.A1(new_n388), .A2(KEYINPUT14), .A3(G116), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n390), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n393), .A2(new_n395), .B1(new_n398), .B2(G107), .ZN(new_n399));
  OR2_X1    g213(.A1(KEYINPUT67), .A2(G128), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT67), .A2(G128), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(G143), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT101), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n269), .A2(G143), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n402), .B2(new_n405), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n406), .A2(new_n407), .A3(G134), .ZN(new_n408));
  INV_X1    g222(.A(G134), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n260), .A2(new_n261), .A3(new_n257), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT101), .B1(new_n410), .B2(new_n404), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n399), .B1(new_n408), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n392), .A2(new_n394), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n395), .A2(new_n390), .A3(new_n391), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n409), .A3(new_n412), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n404), .B(KEYINPUT13), .ZN(new_n419));
  OAI21_X1  g233(.A(G134), .B1(new_n419), .B2(new_n410), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT9), .B(G234), .ZN(new_n422));
  INV_X1    g236(.A(G217), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n422), .A2(new_n423), .A3(G953), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n414), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n424), .B1(new_n414), .B2(new_n421), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n316), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT15), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G478), .ZN(new_n429));
  INV_X1    g243(.A(new_n424), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n398), .A2(G107), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n416), .ZN(new_n432));
  OAI21_X1  g246(.A(G134), .B1(new_n406), .B2(new_n407), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n418), .B2(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n417), .A2(new_n418), .A3(new_n420), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n414), .A2(new_n421), .A3(new_n424), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n428), .A2(G478), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n316), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n429), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT103), .B1(new_n384), .B2(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n429), .A2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n376), .A2(KEYINPUT20), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n382), .A2(new_n378), .A3(new_n368), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n444), .A2(new_n445), .B1(G475), .B2(new_n366), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT103), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n443), .A2(new_n446), .A3(new_n447), .A4(new_n315), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n442), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(G214), .B1(G237), .B2(G902), .ZN(new_n450));
  XOR2_X1   g264(.A(new_n450), .B(KEYINPUT91), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n308), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT74), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n221), .A2(new_n214), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n277), .A2(new_n279), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT11), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n409), .B2(G137), .ZN(new_n458));
  INV_X1    g272(.A(G137), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT11), .A3(G134), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n409), .A2(G137), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G131), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n458), .A2(new_n460), .A3(new_n324), .A4(new_n461), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n456), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n265), .A2(new_n271), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n409), .A2(G137), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n459), .A2(G134), .ZN(new_n469));
  OAI21_X1  g283(.A(G131), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n467), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n455), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT28), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n320), .A2(G210), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n475), .B(KEYINPUT27), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT26), .B(G101), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n280), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n277), .A2(KEYINPUT65), .A3(new_n279), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n465), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n464), .A2(new_n470), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT66), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n464), .A2(new_n470), .A3(KEYINPUT66), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n467), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n455), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT71), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n456), .A2(new_n465), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n471), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n456), .B2(new_n465), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n488), .B1(new_n493), .B2(new_n455), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n474), .B(new_n478), .C1(new_n494), .C2(new_n473), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT29), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n455), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n463), .A2(new_n464), .ZN(new_n499));
  OAI21_X1  g313(.A(KEYINPUT71), .B1(new_n499), .B2(new_n280), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n500), .A2(KEYINPUT30), .A3(new_n490), .A4(new_n471), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT68), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n487), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT68), .B(KEYINPUT30), .C1(new_n482), .C2(new_n487), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n498), .B(new_n501), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n500), .A2(new_n455), .A3(new_n490), .A4(new_n471), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n478), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n454), .B1(new_n497), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n474), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n280), .A2(new_n479), .B1(new_n464), .B2(new_n463), .ZN(new_n512));
  AOI22_X1  g326(.A1(new_n483), .A2(new_n484), .B1(new_n265), .B2(new_n271), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n481), .B1(new_n513), .B2(new_n486), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n508), .B1(new_n455), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n515), .B2(KEYINPUT28), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT29), .B1(new_n516), .B2(new_n478), .ZN(new_n517));
  INV_X1    g331(.A(new_n478), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n501), .A2(new_n498), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n503), .A2(new_n502), .A3(new_n504), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT68), .B1(new_n514), .B2(KEYINPUT30), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n508), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n518), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n517), .A2(new_n524), .A3(KEYINPUT74), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT75), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n472), .A2(new_n526), .A3(new_n473), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n472), .B2(new_n473), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n498), .B1(new_n491), .B2(new_n492), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n508), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT28), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n529), .A2(new_n532), .A3(KEYINPUT29), .A4(new_n478), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n533), .A2(new_n316), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n510), .A2(new_n525), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G472), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n508), .A2(KEYINPUT72), .A3(new_n478), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT72), .B1(new_n508), .B2(new_n478), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT31), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n539), .A2(new_n522), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n508), .A2(new_n478), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n508), .A2(KEYINPUT72), .A3(new_n478), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT31), .B1(new_n546), .B2(new_n507), .ZN(new_n547));
  OAI22_X1  g361(.A1(new_n541), .A2(new_n547), .B1(new_n516), .B2(new_n478), .ZN(new_n548));
  NOR2_X1   g362(.A1(G472), .A2(G902), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(KEYINPUT32), .A3(new_n549), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n516), .A2(new_n478), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n540), .B1(new_n539), .B2(new_n522), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(KEYINPUT31), .A3(new_n507), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n549), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n552), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n536), .A2(new_n550), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G234), .ZN(new_n560));
  OAI21_X1  g374(.A(G217), .B1(new_n560), .B2(G902), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT76), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n262), .A2(G119), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n241), .A2(G128), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT24), .B(G110), .Z(new_n565));
  NAND3_X1  g379(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n330), .A2(new_n331), .A3(KEYINPUT16), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(new_n347), .C1(KEYINPUT16), .C2(new_n330), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n255), .B1(new_n568), .B2(new_n345), .ZN(new_n569));
  INV_X1    g383(.A(new_n351), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n241), .A2(G128), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n564), .B1(new_n572), .B2(KEYINPUT23), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n400), .A2(KEYINPUT23), .A3(G119), .A4(new_n401), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT77), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n262), .A2(new_n576), .A3(KEYINPUT23), .A4(G119), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n573), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(G110), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n565), .B1(new_n563), .B2(new_n564), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n581), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n350), .A2(new_n334), .ZN(new_n583));
  OAI22_X1  g397(.A1(new_n571), .A2(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(G221), .A2(G234), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT80), .B1(new_n585), .B2(G953), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n587), .A2(new_n283), .A3(G221), .A4(G234), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT22), .B(G137), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(new_n586), .A3(new_n588), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  OAI221_X1 g409(.A(new_n566), .B1(new_n578), .B2(new_n579), .C1(new_n569), .C2(new_n570), .ZN(new_n596));
  AOI211_X1 g410(.A(G110), .B(new_n573), .C1(new_n575), .C2(new_n577), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n350), .B(new_n334), .C1(new_n597), .C2(new_n581), .ZN(new_n598));
  INV_X1    g412(.A(new_n594), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT25), .B1(new_n601), .B2(new_n316), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT25), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n603), .B(G902), .C1(new_n595), .C2(new_n600), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n562), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT81), .ZN(new_n606));
  INV_X1    g420(.A(new_n601), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n562), .A2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n562), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n584), .A2(new_n594), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n599), .B1(new_n596), .B2(new_n598), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n316), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n603), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n601), .A2(KEYINPUT25), .A3(new_n316), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n611), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n607), .A2(new_n609), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT81), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n610), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G221), .B1(new_n422), .B2(G902), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n621), .B(KEYINPUT82), .Z(new_n622));
  INV_X1    g436(.A(G469), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(new_n316), .ZN(new_n624));
  XNOR2_X1  g438(.A(G110), .B(G140), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n283), .A2(G227), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n204), .A2(new_n456), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n628), .B1(new_n229), .B2(new_n230), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n272), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n239), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n267), .A2(new_n268), .A3(new_n258), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n264), .A2(new_n269), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n271), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n225), .A3(new_n237), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n630), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n629), .A2(new_n465), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g453(.A1(new_n204), .A2(new_n456), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n250), .B2(new_n251), .ZN(new_n641));
  AOI22_X1  g455(.A1(new_n631), .A2(new_n239), .B1(new_n636), .B2(new_n630), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n499), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n627), .B1(new_n639), .B2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT12), .B1(new_n465), .B2(KEYINPUT89), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n238), .A2(new_n272), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n646), .A2(KEYINPUT88), .A3(new_n636), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n465), .B1(new_n646), .B2(KEYINPUT88), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n467), .B1(new_n225), .B2(new_n237), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT88), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n499), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n645), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n646), .A2(new_n636), .A3(KEYINPUT88), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n649), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n641), .A2(new_n499), .A3(new_n642), .ZN(new_n657));
  INV_X1    g471(.A(new_n627), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n644), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n624), .B1(new_n660), .B2(new_n623), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n627), .B(KEYINPUT83), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n657), .A2(KEYINPUT90), .A3(new_n658), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n465), .B1(new_n629), .B2(new_n638), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(KEYINPUT90), .B1(new_n657), .B2(new_n658), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n664), .B(G469), .C1(new_n667), .C2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n622), .B1(new_n661), .B2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n453), .A2(new_n559), .A3(new_n620), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G101), .ZN(G3));
  INV_X1    g486(.A(new_n659), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n658), .B1(new_n666), .B2(new_n657), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n623), .B(new_n316), .C1(new_n673), .C2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n624), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n675), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n622), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n619), .A2(new_n677), .A3(new_n610), .A4(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n451), .B1(new_n302), .B2(new_n303), .ZN(new_n680));
  AOI21_X1  g494(.A(G478), .B1(new_n438), .B2(new_n316), .ZN(new_n681));
  NOR2_X1   g495(.A1(KEYINPUT104), .A2(KEYINPUT33), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(KEYINPUT104), .A2(KEYINPUT33), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n683), .B(new_n684), .C1(new_n425), .C2(new_n426), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT33), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n436), .A2(new_n686), .A3(new_n687), .A4(new_n437), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n316), .A2(G478), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n681), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n446), .ZN(new_n693));
  INV_X1    g507(.A(new_n303), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n290), .A2(new_n301), .A3(new_n694), .ZN(new_n695));
  AND4_X1   g509(.A1(new_n315), .A2(new_n680), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n556), .B2(G902), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n548), .A2(new_n549), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n679), .A2(new_n696), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT34), .B(G104), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G6));
  NOR2_X1   g517(.A1(new_n384), .A2(new_n443), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n680), .A2(new_n695), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n679), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT35), .B(G107), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G9));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT36), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n710), .B1(new_n594), .B2(new_n711), .ZN(new_n712));
  AOI211_X1 g526(.A(KEYINPUT105), .B(KEYINPUT36), .C1(new_n592), .C2(new_n593), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n584), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n596), .A2(new_n598), .A3(new_n714), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n709), .B1(new_n718), .B2(new_n609), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(KEYINPUT106), .A3(new_n608), .A4(new_n717), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n605), .A2(new_n721), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n697), .A2(new_n698), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n453), .A2(new_n670), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT37), .B(G110), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(KEYINPUT107), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n724), .B(new_n726), .ZN(G12));
  INV_X1    g541(.A(new_n695), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n694), .B1(new_n290), .B2(new_n301), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n310), .B(KEYINPUT108), .Z(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(G900), .B2(new_n313), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n446), .A2(new_n441), .A3(new_n731), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n728), .A2(new_n729), .A3(new_n732), .A4(new_n451), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n559), .A2(new_n733), .A3(new_n670), .A4(new_n722), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G128), .ZN(G30));
  XNOR2_X1  g549(.A(new_n308), .B(KEYINPUT38), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n731), .B(KEYINPUT39), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n670), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(KEYINPUT40), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n719), .A2(new_n720), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n615), .A2(new_n616), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n742), .B2(new_n562), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n443), .A2(new_n446), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n452), .A3(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n737), .A2(new_n740), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n539), .A2(new_n522), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n518), .B2(new_n531), .ZN(new_n748));
  OAI21_X1  g562(.A(G472), .B1(new_n748), .B2(G902), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n550), .A2(new_n558), .A3(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n550), .A2(new_n558), .A3(new_n749), .A4(KEYINPUT109), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n739), .A2(KEYINPUT40), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n746), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G143), .ZN(G45));
  AND2_X1   g571(.A1(new_n550), .A2(new_n558), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n743), .B1(new_n758), .B2(new_n536), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  INV_X1    g574(.A(new_n731), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n692), .A2(new_n446), .A3(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n680), .A2(new_n760), .A3(new_n695), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n302), .A2(new_n303), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n762), .A3(new_n452), .A4(new_n695), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT110), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n759), .A2(new_n670), .A3(new_n763), .A4(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G146), .ZN(G48));
  OAI21_X1  g582(.A(new_n316), .B1(new_n673), .B2(new_n674), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(G469), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n678), .A3(new_n675), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n696), .A2(new_n559), .A3(new_n620), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(KEYINPUT41), .B(G113), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G15));
  NAND4_X1  g589(.A1(new_n559), .A2(new_n705), .A3(new_n620), .A4(new_n772), .ZN(new_n776));
  XNOR2_X1  g590(.A(KEYINPUT111), .B(G116), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G18));
  NAND3_X1  g592(.A1(new_n764), .A2(new_n452), .A3(new_n695), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n771), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n559), .A3(new_n449), .A4(new_n722), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G119), .ZN(G21));
  XOR2_X1   g596(.A(KEYINPUT112), .B(G472), .Z(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n556), .B2(G902), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n529), .A2(new_n532), .ZN(new_n785));
  OAI22_X1  g599(.A1(new_n541), .A2(new_n547), .B1(new_n478), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n549), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n617), .A2(new_n618), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n678), .A2(new_n770), .A3(new_n675), .A4(new_n744), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n728), .A2(new_n729), .A3(new_n451), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n789), .A2(new_n315), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT113), .B(G122), .Z(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G24));
  AND4_X1   g608(.A1(new_n722), .A2(new_n784), .A3(new_n787), .A4(new_n762), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n780), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G125), .ZN(G27));
  INV_X1    g611(.A(KEYINPUT32), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n556), .B2(new_n557), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n550), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(G472), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n533), .A2(new_n316), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n517), .A2(new_n524), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n802), .B1(new_n803), .B2(new_n454), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n801), .B1(new_n804), .B2(new_n525), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n788), .B1(new_n800), .B2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n290), .A2(new_n301), .A3(new_n306), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n306), .B1(new_n290), .B2(new_n301), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n807), .A2(new_n808), .A3(new_n451), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n670), .A2(new_n809), .A3(new_n762), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT42), .B1(new_n806), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n677), .A2(new_n678), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n305), .A2(new_n452), .A3(new_n307), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n762), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT42), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n814), .A2(new_n559), .A3(new_n620), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n324), .ZN(G33));
  NAND2_X1  g633(.A1(new_n559), .A2(new_n620), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n670), .A2(new_n809), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n820), .A2(new_n732), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n409), .ZN(G36));
  OAI21_X1  g637(.A(new_n367), .B1(new_n377), .B2(new_n383), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n692), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT43), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT43), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n699), .A2(new_n722), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n809), .B1(new_n830), .B2(KEYINPUT44), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(KEYINPUT44), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n832), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  INV_X1    g651(.A(new_n675), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT45), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n623), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n676), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT46), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n838), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(KEYINPUT46), .A3(new_n676), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n678), .ZN(new_n848));
  INV_X1    g662(.A(new_n738), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n622), .B1(new_n845), .B2(new_n846), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(KEYINPUT114), .A3(new_n738), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n836), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n459), .ZN(G39));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n848), .B1(new_n855), .B2(KEYINPUT47), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT116), .B(KEYINPUT47), .Z(new_n857));
  NAND2_X1  g671(.A1(new_n851), .A2(new_n857), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n559), .A2(new_n620), .A3(new_n813), .A4(new_n815), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT117), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(G140), .ZN(G42));
  NAND3_X1  g676(.A1(new_n559), .A2(new_n670), .A3(new_n722), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n766), .A2(new_n763), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n734), .B(new_n796), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT120), .B1(new_n722), .B2(new_n761), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n743), .A2(new_n867), .A3(new_n731), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n670), .A3(new_n791), .A4(new_n744), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n870), .B1(new_n752), .B2(new_n753), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT52), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n734), .A2(new_n796), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n867), .B1(new_n743), .B2(new_n731), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n617), .A2(new_n741), .A3(KEYINPUT120), .A4(new_n761), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n680), .A2(new_n695), .A3(new_n744), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n877), .A2(new_n812), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n754), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n873), .A2(new_n874), .A3(new_n767), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n872), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n315), .B(new_n452), .C1(new_n807), .C2(new_n808), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  OR3_X1    g698(.A1(new_n692), .A2(new_n446), .A3(KEYINPUT118), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n692), .B2(new_n446), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n429), .A2(KEYINPUT119), .A3(new_n440), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT119), .B1(new_n429), .B2(new_n440), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n446), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n679), .A2(new_n884), .A3(new_n700), .A4(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n671), .A2(new_n891), .A3(new_n724), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n795), .ZN(new_n895));
  NOR4_X1   g709(.A1(new_n887), .A2(new_n888), .A3(new_n824), .A4(new_n761), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n550), .A2(new_n558), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n722), .B(new_n896), .C1(new_n897), .C2(new_n805), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n821), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n822), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n734), .A2(new_n796), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT52), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n882), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n773), .A2(new_n781), .A3(new_n776), .A4(new_n792), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n818), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n905), .A2(new_n906), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT123), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n910), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n908), .A4(new_n907), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n904), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n818), .A2(new_n822), .A3(new_n899), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n905), .A2(new_n892), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n872), .A3(new_n918), .A4(new_n881), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n919), .A2(KEYINPUT121), .A3(new_n893), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT121), .B1(new_n919), .B2(new_n893), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n915), .B(new_n916), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n893), .ZN(new_n923));
  AOI21_X1  g737(.A(KEYINPUT53), .B1(new_n901), .B2(KEYINPUT52), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(new_n806), .ZN(new_n928));
  INV_X1    g742(.A(new_n730), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n827), .A2(new_n929), .A3(new_n829), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n813), .A2(new_n771), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n928), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT48), .ZN(new_n934));
  INV_X1    g748(.A(new_n754), .ZN(new_n935));
  INV_X1    g749(.A(new_n620), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n936), .A2(new_n310), .A3(new_n771), .A4(new_n813), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n935), .A2(new_n937), .A3(new_n693), .ZN(new_n938));
  INV_X1    g752(.A(G952), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n931), .A2(new_n789), .ZN(new_n940));
  AOI211_X1 g754(.A(new_n939), .B(G953), .C1(new_n940), .C2(new_n780), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n809), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n856), .A2(new_n858), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n660), .A2(new_n623), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n946), .A2(new_n838), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n622), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n940), .A2(new_n451), .A3(new_n737), .A4(new_n772), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT50), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n935), .A2(new_n937), .A3(new_n446), .A4(new_n692), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(KEYINPUT50), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n784), .A2(new_n787), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n931), .A2(new_n722), .A3(new_n954), .A4(new_n932), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n943), .B1(new_n949), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n942), .B1(new_n957), .B2(KEYINPUT51), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n927), .B(new_n958), .C1(KEYINPUT51), .C2(new_n957), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(G952), .B2(G953), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT49), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n947), .A2(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n947), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n788), .A2(new_n678), .A3(new_n452), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n826), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n935), .A2(new_n737), .A3(new_n962), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n960), .A2(new_n966), .ZN(G75));
  NOR2_X1   g781(.A1(new_n283), .A2(G952), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n923), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n919), .A2(KEYINPUT121), .A3(new_n893), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n316), .B1(new_n973), .B2(new_n915), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT56), .B1(new_n974), .B2(G210), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n254), .A2(new_n289), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n287), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT55), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n969), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n980), .B1(new_n975), .B2(new_n979), .ZN(G51));
  AOI21_X1  g795(.A(new_n916), .B1(new_n973), .B2(new_n915), .ZN(new_n982));
  INV_X1    g796(.A(new_n922), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n624), .B(KEYINPUT57), .Z(new_n985));
  OAI22_X1  g799(.A1(new_n984), .A2(new_n985), .B1(new_n674), .B2(new_n673), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n974), .B(new_n841), .C1(new_n840), .C2(new_n839), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n968), .B1(new_n986), .B2(new_n987), .ZN(G54));
  NAND3_X1  g802(.A1(new_n974), .A2(KEYINPUT58), .A3(G475), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(new_n381), .A3(new_n380), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n974), .A2(KEYINPUT58), .A3(G475), .A4(new_n382), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n990), .A2(new_n991), .A3(new_n969), .ZN(G60));
  INV_X1    g806(.A(new_n689), .ZN(new_n993));
  NAND2_X1  g807(.A1(G478), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT59), .Z(new_n995));
  NOR2_X1   g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n982), .B2(new_n983), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n998), .A3(new_n969), .ZN(new_n999));
  INV_X1    g813(.A(new_n996), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT54), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(new_n922), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT125), .B1(new_n1003), .B2(new_n968), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n993), .B1(new_n927), .B2(new_n995), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n999), .A2(new_n1004), .A3(new_n1005), .ZN(G63));
  NAND2_X1  g820(.A1(G217), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT60), .Z(new_n1008));
  NAND2_X1  g822(.A1(new_n1001), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n968), .B1(new_n1009), .B2(new_n607), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1010), .B1(new_n718), .B2(new_n1009), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1010), .B(KEYINPUT61), .C1(new_n718), .C2(new_n1009), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(G66));
  INV_X1    g829(.A(G224), .ZN(new_n1016));
  OAI21_X1  g830(.A(G953), .B1(new_n311), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n918), .B2(G953), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n976), .B1(G898), .B2(new_n283), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1018), .B(new_n1019), .ZN(G69));
  AOI21_X1  g834(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n818), .A2(new_n822), .ZN(new_n1023));
  NOR3_X1   g837(.A1(new_n853), .A2(new_n865), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n850), .A2(new_n852), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1025), .A2(new_n791), .A3(new_n744), .A4(new_n928), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n861), .A2(new_n1024), .A3(new_n283), .A4(new_n1026), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n371), .B1(new_n335), .B2(new_n372), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1028), .B(new_n1029), .Z(new_n1030));
  AOI21_X1  g844(.A(new_n1030), .B1(G900), .B2(G953), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT126), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1022), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n890), .A2(new_n809), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n820), .A2(new_n739), .A3(new_n1035), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n853), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n756), .A2(new_n767), .A3(new_n873), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n861), .A2(new_n1037), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n283), .ZN(new_n1042));
  AOI22_X1  g856(.A1(new_n1042), .A2(new_n1030), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1034), .B(new_n1043), .ZN(G72));
  NAND2_X1  g858(.A1(G472), .A2(G902), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT63), .Z(new_n1046));
  INV_X1    g860(.A(new_n918), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n1046), .B1(new_n1041), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g862(.A(new_n1048), .B(new_n478), .C1(new_n523), .C2(new_n522), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n861), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1046), .B1(new_n1050), .B2(new_n1047), .ZN(new_n1051));
  NAND4_X1  g865(.A1(new_n1051), .A2(new_n508), .A3(new_n518), .A4(new_n507), .ZN(new_n1052));
  INV_X1    g866(.A(new_n1046), .ZN(new_n1053));
  INV_X1    g867(.A(new_n747), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1053), .B1(new_n1054), .B2(new_n524), .ZN(new_n1055));
  AOI21_X1  g869(.A(new_n968), .B1(new_n925), .B2(new_n1055), .ZN(new_n1056));
  AND3_X1   g870(.A1(new_n1049), .A2(new_n1052), .A3(new_n1056), .ZN(G57));
endmodule


