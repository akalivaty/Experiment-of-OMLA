//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:24 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  AOI21_X1  g004(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n191));
  NAND2_X1  g005(.A1(KEYINPUT18), .A2(G131), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G214), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n197), .B2(new_n189), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT80), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT64), .B(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n199), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT96), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n199), .A2(new_n212), .A3(KEYINPUT96), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n190), .A2(new_n191), .A3(G131), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n219), .B1(new_n197), .B2(new_n189), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT17), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT99), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n207), .A2(KEYINPUT16), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n201), .A2(KEYINPUT16), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(G146), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(G146), .B1(new_n225), .B2(new_n226), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n229), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT99), .A3(new_n227), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n223), .A2(new_n230), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n217), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G113), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(G104), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n217), .A2(new_n238), .A3(new_n234), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G902), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n187), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(G475), .A2(G902), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n245), .B(KEYINPUT100), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n199), .A2(new_n212), .A3(KEYINPUT96), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT96), .B1(new_n199), .B2(new_n212), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n227), .B1(new_n218), .B2(new_n220), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT19), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n206), .A2(new_n208), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n204), .A2(KEYINPUT19), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n209), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT97), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n252), .A2(KEYINPUT97), .A3(new_n209), .A4(new_n253), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(KEYINPUT98), .B(new_n239), .C1(new_n249), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n241), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n256), .A2(new_n257), .ZN(new_n261));
  INV_X1    g075(.A(new_n250), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n217), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT98), .B1(new_n264), .B2(new_n239), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n246), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT20), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT20), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n268), .B(new_n246), .C1(new_n260), .C2(new_n265), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n244), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G953), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(G952), .ZN(new_n272));
  NAND2_X1  g086(.A1(G234), .A2(G237), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(G902), .A3(G953), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  XNOR2_X1  g091(.A(KEYINPUT21), .B(G898), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT9), .B(G234), .ZN(new_n281));
  INV_X1    g095(.A(G217), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n281), .A2(new_n282), .A3(G953), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT106), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G107), .ZN(new_n286));
  INV_X1    g100(.A(G116), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G116), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(new_n290), .A3(G122), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT101), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT101), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n288), .A2(new_n290), .A3(new_n293), .A4(G122), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n287), .A2(G122), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT102), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT102), .ZN(new_n299));
  AOI211_X1 g113(.A(new_n299), .B(new_n296), .C1(new_n292), .C2(new_n294), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n286), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G128), .B(G143), .ZN(new_n302));
  INV_X1    g116(.A(G134), .ZN(new_n303));
  XNOR2_X1  g117(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT104), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT14), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n307), .B1(new_n292), .B2(new_n294), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n308), .B2(new_n296), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT70), .B(G116), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n293), .B1(new_n310), .B2(G122), .ZN(new_n311));
  AND4_X1   g125(.A1(new_n293), .A2(new_n288), .A3(new_n290), .A4(G122), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT14), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(KEYINPUT104), .A3(new_n297), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT105), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n292), .A2(new_n315), .A3(new_n307), .A4(new_n294), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT105), .B1(new_n295), .B2(KEYINPUT14), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n309), .A2(new_n314), .A3(new_n316), .A4(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n305), .B1(G107), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT103), .B(KEYINPUT13), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(G134), .C1(G128), .C2(new_n196), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n304), .B(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(new_n298), .ZN(new_n323));
  INV_X1    g137(.A(new_n300), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G107), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n322), .B1(new_n325), .B2(new_n301), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n285), .B1(new_n319), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n318), .A2(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n301), .A3(new_n304), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n301), .ZN(new_n330));
  INV_X1    g144(.A(new_n322), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n329), .A2(new_n332), .A3(new_n284), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n243), .ZN(new_n335));
  INV_X1    g149(.A(G478), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(KEYINPUT15), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n334), .B(new_n243), .C1(KEYINPUT15), .C2(new_n336), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n270), .A2(new_n280), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT107), .ZN(new_n341));
  AND2_X1   g155(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT107), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n342), .A2(new_n343), .A3(new_n280), .A4(new_n270), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n346));
  INV_X1    g160(.A(G119), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G128), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(new_n347), .A3(G128), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n349), .B(new_n351), .C1(new_n347), .C2(G128), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT79), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT24), .B(G110), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G128), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT23), .A3(G119), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n347), .A2(G128), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n348), .B(new_n358), .C1(new_n359), .C2(KEYINPUT23), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n360), .A2(G110), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n227), .B(new_n210), .C1(new_n356), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n353), .A2(new_n355), .ZN(new_n363));
  AOI22_X1  g177(.A1(new_n231), .A2(new_n227), .B1(G110), .B2(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n271), .A2(G221), .A3(G234), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT81), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT22), .B(G137), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n365), .A3(new_n370), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n346), .B1(new_n374), .B2(G902), .ZN(new_n375));
  INV_X1    g189(.A(new_n346), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n372), .A2(new_n243), .A3(new_n373), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(G234), .ZN(new_n380));
  OAI21_X1  g194(.A(G217), .B1(new_n380), .B2(G902), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT77), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n374), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n243), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G146), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(KEYINPUT64), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT64), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G146), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n392), .A3(G143), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n196), .A2(G146), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n357), .A2(KEYINPUT1), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n357), .B1(new_n393), .B2(KEYINPUT1), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n196), .A2(G146), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n390), .A2(new_n392), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n196), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n396), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT72), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(KEYINPUT72), .B(new_n396), .C1(new_n397), .C2(new_n400), .ZN(new_n404));
  INV_X1    g218(.A(G137), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT66), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT66), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G137), .ZN(new_n408));
  AOI21_X1  g222(.A(G134), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n303), .A2(G137), .ZN(new_n410));
  OAI21_X1  g224(.A(G131), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT68), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n413), .B(G131), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT11), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT65), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n416), .B(new_n418), .C1(new_n303), .C2(G137), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n417), .A2(new_n303), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n406), .A3(new_n408), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n303), .A2(G137), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n219), .A4(new_n422), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n403), .A2(new_n404), .A3(new_n412), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n398), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n426), .B1(new_n209), .B2(G143), .ZN(new_n427));
  AND2_X1   g241(.A1(KEYINPUT0), .A2(G128), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT0), .A2(G128), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n393), .A2(new_n394), .A3(new_n428), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n219), .A2(KEYINPUT67), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT66), .B(G137), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n434), .A2(new_n420), .B1(new_n303), .B2(G137), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n433), .B1(new_n435), .B2(new_n419), .ZN(new_n436));
  AND4_X1   g250(.A1(new_n419), .A2(new_n421), .A3(new_n422), .A4(new_n433), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n431), .B(new_n432), .C1(new_n436), .C2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n425), .A2(KEYINPUT30), .A3(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n401), .A2(new_n412), .A3(new_n423), .A4(new_n414), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT30), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT69), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n445));
  INV_X1    g259(.A(G113), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(KEYINPUT69), .A2(KEYINPUT2), .A3(G113), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n445), .B2(new_n446), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n288), .A2(new_n290), .A3(G119), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n287), .A2(G119), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT71), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n450), .A2(KEYINPUT71), .A3(new_n452), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n449), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n451), .B1(new_n310), .B2(G119), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n449), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n439), .A2(new_n443), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n425), .A2(new_n461), .A3(new_n438), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT26), .B(G101), .Z(new_n465));
  NAND2_X1  g279(.A1(new_n188), .A2(G210), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n464), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT31), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n463), .A2(KEYINPUT31), .A3(new_n464), .A4(new_n470), .ZN(new_n474));
  INV_X1    g288(.A(new_n464), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n461), .B1(new_n438), .B2(new_n440), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT28), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT28), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n464), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT74), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT74), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n464), .A2(new_n481), .A3(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n473), .A2(new_n474), .B1(new_n483), .B2(new_n469), .ZN(new_n484));
  NOR2_X1   g298(.A1(G472), .A2(G902), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n485), .B(KEYINPUT75), .Z(new_n486));
  OAI21_X1  g300(.A(KEYINPUT32), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n473), .A2(new_n474), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(new_n469), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT32), .ZN(new_n491));
  INV_X1    g305(.A(new_n486), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n461), .B1(new_n425), .B2(new_n438), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT28), .B1(new_n475), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n469), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n496), .A2(new_n480), .A3(new_n482), .A4(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(new_n243), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n463), .A2(new_n464), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n469), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT76), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT76), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n501), .A2(new_n504), .A3(new_n469), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n497), .B1(new_n483), .B2(new_n469), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G472), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n388), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G210), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G110), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT8), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT3), .B1(new_n237), .B2(G107), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT3), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n286), .A3(G104), .ZN(new_n517));
  INV_X1    g331(.A(G101), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n237), .A2(G107), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n515), .A2(new_n517), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n286), .A2(G104), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n237), .A2(G107), .ZN(new_n522));
  OAI21_X1  g336(.A(G101), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT84), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT84), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT92), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT5), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n446), .B1(new_n451), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n450), .A2(KEYINPUT5), .A3(new_n452), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n531), .A2(new_n532), .B1(new_n458), .B2(new_n449), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n528), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n455), .A2(KEYINPUT5), .A3(new_n456), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n460), .B1(new_n535), .B2(new_n531), .ZN(new_n536));
  INV_X1    g350(.A(new_n524), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n520), .A2(new_n523), .A3(new_n526), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n526), .B1(new_n520), .B2(new_n523), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n532), .A2(new_n531), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n459), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT92), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n514), .B1(new_n538), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n393), .A2(KEYINPUT1), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G128), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n393), .A2(new_n394), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n548), .A2(new_n427), .B1(new_n549), .B2(new_n395), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n202), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n202), .B1(new_n431), .B2(new_n432), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT91), .B(G224), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n555), .A2(new_n271), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n558), .B1(new_n552), .B2(KEYINPUT93), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n554), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n551), .A2(new_n553), .A3(KEYINPUT93), .A4(new_n558), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT94), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n546), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n535), .A2(new_n531), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n528), .A3(new_n459), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n515), .A2(new_n517), .A3(new_n519), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT83), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n515), .A2(new_n517), .A3(KEYINPUT83), .A4(new_n519), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(G101), .A3(new_n570), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n520), .A2(KEYINPUT4), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n518), .A2(KEYINPUT4), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n573), .B(new_n575), .C1(new_n457), .C2(new_n460), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n566), .A2(new_n576), .A3(new_n513), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n564), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n544), .B(new_n534), .C1(new_n537), .C2(new_n536), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(new_n514), .B1(new_n560), .B2(new_n561), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n563), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n243), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n566), .A2(new_n576), .ZN(new_n583));
  INV_X1    g397(.A(new_n513), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(KEYINPUT6), .A3(new_n577), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n554), .B(new_n556), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n513), .B1(new_n566), .B2(new_n576), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT90), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT89), .B(KEYINPUT6), .Z(new_n590));
  AND3_X1   g404(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n586), .B(new_n587), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n512), .B1(new_n582), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n596));
  INV_X1    g410(.A(new_n577), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n580), .B2(new_n563), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n546), .A2(new_n562), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(KEYINPUT94), .ZN(new_n600));
  AOI21_X1  g414(.A(G902), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n511), .A3(new_n593), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n595), .A2(new_n596), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G214), .B1(G237), .B2(G902), .ZN(new_n604));
  OAI211_X1 g418(.A(KEYINPUT95), .B(new_n512), .C1(new_n582), .C2(new_n594), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n345), .A2(new_n510), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(G221), .B1(new_n281), .B2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(G110), .B(G140), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n271), .A2(G227), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT10), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n525), .B2(new_n527), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(new_n403), .A3(new_n404), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n436), .A2(new_n437), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n431), .A2(new_n432), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n573), .A3(new_n575), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n393), .A2(new_n394), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT1), .ZN(new_n621));
  OAI21_X1  g435(.A(G128), .B1(new_n398), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n396), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n537), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n614), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n616), .A2(new_n617), .A3(new_n619), .A4(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT85), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n575), .A2(new_n431), .A3(new_n432), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n630), .A2(new_n573), .B1(new_n625), .B2(new_n614), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(KEYINPUT85), .A3(new_n617), .A4(new_n616), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT12), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n541), .A2(new_n550), .B1(new_n537), .B2(new_n624), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n634), .B1(new_n635), .B2(new_n617), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n625), .B1(new_n528), .B2(new_n401), .ZN(new_n637));
  INV_X1    g451(.A(new_n617), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(KEYINPUT12), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n633), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT86), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n633), .A2(KEYINPUT86), .A3(new_n640), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n613), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n612), .B1(new_n629), .B2(new_n632), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n631), .A2(new_n616), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n638), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(KEYINPUT87), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  AOI221_X4 g465(.A(new_n642), .B1(new_n636), .B2(new_n639), .C1(new_n629), .C2(new_n632), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT86), .B1(new_n633), .B2(new_n640), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n612), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT87), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n654), .A2(new_n655), .A3(new_n649), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n651), .A2(G469), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(G469), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n243), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n633), .A2(new_n648), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n612), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n646), .A2(new_n640), .ZN(new_n662));
  AOI21_X1  g476(.A(G902), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n659), .B1(new_n663), .B2(new_n658), .ZN(new_n664));
  AOI211_X1 g478(.A(KEYINPUT88), .B(new_n609), .C1(new_n657), .C2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT88), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n657), .A2(new_n664), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n666), .B1(new_n667), .B2(new_n608), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n607), .B1(new_n665), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G101), .ZN(G3));
  AOI22_X1  g484(.A1(new_n379), .A2(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n484), .B2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n490), .A2(new_n492), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n671), .B(new_n675), .C1(new_n668), .C2(new_n665), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n336), .A2(G902), .ZN(new_n677));
  AOI21_X1  g491(.A(KEYINPUT33), .B1(new_n334), .B2(KEYINPUT108), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT33), .ZN(new_n680));
  AOI211_X1 g494(.A(new_n679), .B(new_n680), .C1(new_n327), .C2(new_n333), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n677), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n335), .A2(new_n336), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n270), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n595), .A2(new_n602), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n604), .A3(new_n280), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n676), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(KEYINPUT34), .B(G104), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  NAND2_X1  g504(.A1(new_n338), .A2(new_n339), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n270), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n676), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(KEYINPUT35), .B(G107), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G9));
  NOR2_X1   g509(.A1(new_n371), .A2(KEYINPUT36), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n366), .B(new_n696), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n379), .A2(new_n382), .B1(new_n386), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n345), .A2(new_n606), .A3(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(new_n675), .C1(new_n665), .C2(new_n668), .ZN(new_n701));
  XOR2_X1   g515(.A(KEYINPUT37), .B(G110), .Z(new_n702));
  XNOR2_X1  g516(.A(new_n701), .B(new_n702), .ZN(G12));
  NAND2_X1  g517(.A1(new_n494), .A2(new_n509), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n275), .B1(new_n277), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n692), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n604), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n595), .B2(new_n602), .ZN(new_n709));
  AND4_X1   g523(.A1(new_n704), .A2(new_n707), .A3(new_n709), .A4(new_n699), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n668), .B2(new_n665), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  NAND2_X1  g526(.A1(new_n603), .A2(new_n605), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n469), .B1(new_n475), .B2(new_n495), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n471), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g530(.A(G902), .B1(new_n716), .B2(KEYINPUT109), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n717), .B1(KEYINPUT109), .B2(new_n716), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G472), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n494), .A2(KEYINPUT110), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT110), .B1(new_n494), .B2(new_n719), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n244), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT98), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n249), .A2(new_n258), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n724), .B1(new_n725), .B2(new_n238), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n241), .A3(new_n259), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n268), .B1(new_n727), .B2(new_n246), .ZN(new_n728));
  INV_X1    g542(.A(new_n269), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n723), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n691), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n698), .A2(new_n604), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n714), .A2(new_n722), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT40), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n706), .B(KEYINPUT39), .Z(new_n735));
  OAI211_X1 g549(.A(new_n734), .B(new_n735), .C1(new_n668), .C2(new_n665), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n735), .B1(new_n668), .B2(new_n665), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT40), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G143), .ZN(G45));
  INV_X1    g554(.A(new_n706), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n684), .A2(KEYINPUT111), .A3(new_n709), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n698), .B1(new_n494), .B2(new_n509), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n684), .A2(new_n741), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n686), .A2(new_n604), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n744), .B(new_n748), .C1(new_n668), .C2(new_n665), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  INV_X1    g564(.A(new_n687), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n663), .A2(new_n658), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n663), .A2(new_n658), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n752), .A2(new_n608), .A3(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n510), .A2(new_n751), .A3(new_n684), .A4(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(KEYINPUT41), .B(G113), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G15));
  NOR2_X1   g571(.A1(new_n687), .A2(new_n692), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n510), .A3(new_n754), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT112), .B(G116), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G18));
  NAND4_X1  g575(.A1(new_n345), .A2(new_n743), .A3(new_n709), .A4(new_n754), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G119), .ZN(G21));
  NOR2_X1   g577(.A1(new_n747), .A2(new_n731), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n496), .A2(new_n480), .A3(new_n482), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n469), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n488), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT113), .A3(new_n492), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n473), .A2(new_n474), .B1(new_n765), .B2(new_n469), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n486), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n671), .A2(new_n672), .A3(new_n768), .A4(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n764), .A2(new_n772), .A3(new_n280), .A4(new_n754), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  INV_X1    g588(.A(new_n754), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n747), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n699), .A2(new_n672), .A3(new_n768), .A4(new_n771), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n746), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  AOI21_X1  g594(.A(new_n708), .B1(new_n603), .B2(new_n605), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n654), .A2(G469), .A3(new_n649), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n609), .B1(new_n664), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  AOI211_X1 g598(.A(new_n706), .B(new_n270), .C1(new_n682), .C2(new_n683), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(KEYINPUT42), .A3(new_n510), .A4(new_n785), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n510), .A2(new_n785), .A3(new_n783), .A4(new_n781), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n786), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G131), .ZN(G33));
  AND4_X1   g605(.A1(new_n510), .A2(new_n707), .A3(new_n783), .A4(new_n781), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(new_n303), .ZN(G36));
  AOI21_X1  g607(.A(KEYINPUT45), .B1(new_n651), .B2(new_n656), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT114), .B1(new_n794), .B2(new_n658), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT45), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n654), .A2(new_n655), .A3(new_n649), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n655), .B1(new_n654), .B2(new_n649), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT114), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n799), .A2(new_n800), .A3(G469), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n654), .A2(KEYINPUT45), .A3(new_n649), .ZN(new_n802));
  XOR2_X1   g616(.A(new_n802), .B(KEYINPUT115), .Z(new_n803));
  NAND3_X1  g617(.A1(new_n795), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n659), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT46), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n805), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n808), .A2(new_n753), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n675), .A2(new_n698), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n682), .A2(new_n683), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n730), .A2(KEYINPUT117), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n270), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT43), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n682), .A2(new_n819), .A3(new_n683), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n730), .A2(KEYINPUT43), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n811), .A2(new_n817), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT44), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n817), .A2(new_n811), .A3(new_n822), .A4(KEYINPUT44), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n825), .A2(new_n781), .A3(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n810), .A2(new_n608), .A3(new_n735), .A4(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G137), .ZN(G39));
  XOR2_X1   g643(.A(KEYINPUT118), .B(KEYINPUT47), .Z(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n810), .A2(new_n608), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n781), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n833), .A2(new_n746), .A3(new_n704), .A4(new_n671), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT119), .ZN(new_n835));
  INV_X1    g649(.A(new_n753), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n806), .B2(new_n807), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n609), .B1(new_n837), .B2(new_n809), .ZN(new_n838));
  NOR2_X1   g652(.A1(KEYINPUT118), .A2(KEYINPUT47), .ZN(new_n839));
  OAI211_X1 g653(.A(new_n832), .B(new_n835), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n840), .B(G140), .ZN(G42));
  AND2_X1   g655(.A1(new_n752), .A2(new_n753), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(KEYINPUT49), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(KEYINPUT49), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n671), .A2(new_n608), .A3(new_n604), .ZN(new_n846));
  NOR4_X1   g660(.A1(new_n844), .A2(new_n845), .A3(new_n816), .A4(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n714), .A3(new_n722), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n817), .A2(new_n822), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n275), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n775), .A2(new_n833), .ZN(new_n851));
  INV_X1    g665(.A(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n777), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n850), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n775), .A2(new_n604), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n714), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n854), .A2(new_n857), .A3(KEYINPUT50), .A4(new_n772), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n849), .A2(new_n275), .A3(new_n772), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n856), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n851), .A2(new_n722), .A3(new_n671), .A4(new_n275), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n812), .A2(new_n730), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n863), .A2(KEYINPUT122), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n863), .B2(new_n865), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n862), .A2(KEYINPUT51), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n843), .A2(new_n608), .ZN(new_n870));
  INV_X1    g684(.A(new_n839), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n804), .A2(KEYINPUT46), .A3(new_n805), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT46), .B1(new_n804), .B2(new_n805), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n872), .A2(new_n873), .A3(new_n836), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n871), .B1(new_n874), .B2(new_n609), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n870), .B1(new_n875), .B2(new_n832), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n860), .A2(new_n833), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n869), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n854), .A2(new_n772), .A3(new_n776), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n880), .B(new_n272), .C1(new_n685), .C2(new_n863), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n854), .A2(new_n510), .A3(new_n851), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(KEYINPUT48), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n862), .A2(new_n868), .ZN(new_n886));
  INV_X1    g700(.A(new_n870), .ZN(new_n887));
  AOI211_X1 g701(.A(new_n609), .B(new_n830), .C1(new_n837), .C2(new_n809), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n839), .B1(new_n810), .B2(new_n608), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n886), .B1(new_n890), .B2(new_n877), .ZN(new_n891));
  OAI211_X1 g705(.A(new_n879), .B(new_n885), .C1(new_n891), .C2(KEYINPUT51), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT54), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n711), .A2(new_n779), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n783), .A2(new_n698), .A3(new_n741), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n764), .C1(new_n721), .C2(new_n720), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n894), .A2(KEYINPUT52), .A3(new_n749), .A4(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n749), .A2(new_n711), .A3(new_n779), .A4(new_n896), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n792), .B1(new_n786), .B2(new_n789), .ZN(new_n902));
  AND4_X1   g716(.A1(new_n755), .A2(new_n762), .A3(new_n773), .A4(new_n759), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n778), .A2(new_n784), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n691), .A2(new_n730), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n743), .A2(new_n905), .A3(new_n741), .A4(new_n781), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n907), .B1(new_n665), .B2(new_n668), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n902), .A2(new_n903), .A3(new_n904), .A4(new_n908), .ZN(new_n909));
  AOI22_X1  g723(.A1(new_n685), .A2(KEYINPUT120), .B1(new_n691), .B2(new_n270), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n910), .B1(KEYINPUT120), .B2(new_n685), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n713), .A2(new_n708), .A3(new_n279), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n701), .B(new_n669), .C1(new_n676), .C2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n901), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n901), .A2(KEYINPUT121), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n901), .B(new_n915), .C1(KEYINPUT121), .C2(KEYINPUT53), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n893), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n901), .A2(new_n915), .A3(KEYINPUT53), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT53), .B1(new_n901), .B2(new_n915), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT54), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n892), .A2(new_n921), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(G952), .A2(G953), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n848), .B1(new_n925), .B2(new_n926), .ZN(G75));
  XNOR2_X1  g741(.A(new_n898), .B(KEYINPUT52), .ZN(new_n928));
  INV_X1    g742(.A(new_n668), .ZN(new_n929));
  INV_X1    g743(.A(new_n665), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n906), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n762), .A2(new_n773), .A3(new_n759), .A4(new_n755), .ZN(new_n932));
  INV_X1    g746(.A(new_n904), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n701), .A2(new_n669), .ZN(new_n935));
  OR2_X1    g749(.A1(new_n913), .A2(new_n676), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n935), .A3(new_n936), .A4(new_n902), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n918), .B1(new_n928), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n901), .A2(new_n915), .A3(KEYINPUT53), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(G210), .A3(G902), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n587), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT55), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n945), .B1(new_n941), .B2(new_n942), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n271), .A2(G952), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(G51));
  XNOR2_X1  g763(.A(new_n659), .B(KEYINPUT57), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n893), .B1(new_n938), .B2(new_n939), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n924), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n661), .A2(new_n662), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n953), .B(KEYINPUT123), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n940), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n956), .A2(new_n243), .A3(new_n804), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n948), .B1(new_n955), .B2(new_n957), .ZN(G54));
  NAND4_X1  g772(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n959));
  INV_X1    g773(.A(new_n727), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n962), .A3(new_n948), .ZN(G60));
  NAND2_X1  g777(.A1(G478), .A2(G902), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT59), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n678), .B2(new_n681), .ZN(new_n966));
  OAI21_X1  g780(.A(KEYINPUT54), .B1(new_n922), .B2(new_n923), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n938), .A2(new_n893), .A3(new_n939), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n965), .B1(new_n921), .B2(new_n924), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n678), .A2(new_n681), .ZN(new_n971));
  AOI211_X1 g785(.A(new_n948), .B(new_n969), .C1(new_n970), .C2(new_n971), .ZN(G63));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT60), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n974), .B1(new_n938), .B2(new_n939), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n975), .A2(new_n384), .ZN(new_n976));
  INV_X1    g790(.A(new_n948), .ZN(new_n977));
  INV_X1    g791(.A(new_n974), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n697), .B(new_n978), .C1(new_n922), .C2(new_n923), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n976), .A2(KEYINPUT61), .A3(new_n977), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(new_n977), .C1(new_n975), .C2(new_n384), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n980), .A2(new_n983), .ZN(G66));
  INV_X1    g798(.A(new_n278), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n271), .B1(new_n985), .B2(new_n555), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n914), .A2(new_n932), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n986), .B1(new_n988), .B2(new_n271), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n943), .B1(G898), .B2(new_n271), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n989), .B(new_n990), .Z(G69));
  NAND2_X1  g805(.A1(new_n439), .A2(new_n443), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n252), .A2(new_n253), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n911), .A2(new_n510), .A3(new_n781), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(new_n737), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n828), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT124), .ZN(new_n999));
  AND3_X1   g813(.A1(new_n749), .A2(new_n711), .A3(new_n779), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n739), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n739), .A2(KEYINPUT62), .A3(new_n1000), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT124), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n828), .A2(new_n1006), .A3(new_n997), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n999), .A2(new_n1005), .A3(new_n840), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n995), .B1(new_n1009), .B2(G953), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n838), .A2(new_n510), .A3(new_n735), .A4(new_n764), .ZN(new_n1011));
  AND3_X1   g825(.A1(new_n894), .A2(new_n749), .A3(new_n902), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1011), .A2(new_n828), .A3(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(G953), .B1(new_n1013), .B2(new_n840), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n705), .A2(G953), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT125), .Z(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n994), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(G227), .A2(G900), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(G953), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1010), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n828), .A2(new_n1012), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1022), .A2(new_n840), .A3(new_n1011), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(new_n271), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1024), .A2(new_n1016), .ZN(new_n1025));
  OAI211_X1 g839(.A(G953), .B(new_n1019), .C1(new_n1025), .C2(new_n995), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1021), .A2(new_n1026), .ZN(G72));
  NAND4_X1  g841(.A1(new_n1022), .A2(new_n840), .A3(new_n987), .A4(new_n1011), .ZN(new_n1028));
  NAND2_X1  g842(.A1(G472), .A2(G902), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT63), .Z(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(KEYINPUT126), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT126), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1028), .A2(new_n1033), .A3(new_n1030), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n501), .A2(new_n470), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1030), .B1(new_n1008), .B2(new_n988), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n469), .B1(new_n463), .B2(new_n464), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n919), .A2(new_n920), .ZN(new_n1040));
  NAND3_X1  g854(.A1(new_n503), .A2(new_n471), .A3(new_n505), .ZN(new_n1041));
  AND2_X1   g855(.A1(new_n1041), .A2(new_n1030), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n948), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g857(.A1(new_n1036), .A2(new_n1039), .A3(new_n1043), .ZN(G57));
endmodule


