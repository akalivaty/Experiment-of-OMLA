

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(n546), .A2(G2105), .ZN(n595) );
  OR2_X1 U553 ( .A1(n742), .A2(n741), .ZN(n747) );
  XNOR2_X1 U554 ( .A(n757), .B(KEYINPUT107), .ZN(n758) );
  XNOR2_X1 U555 ( .A(n759), .B(n758), .ZN(n775) );
  NOR2_X1 U556 ( .A1(G651), .A2(n617), .ZN(n635) );
  XOR2_X1 U557 ( .A(KEYINPUT17), .B(n543), .Z(n880) );
  NOR2_X1 U558 ( .A1(G651), .A2(G543), .ZN(n639) );
  AND2_X1 U559 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U560 ( .A(G57), .ZN(G237) );
  INV_X1 U561 ( .A(G108), .ZN(G238) );
  INV_X1 U562 ( .A(G120), .ZN(G236) );
  XOR2_X1 U563 ( .A(KEYINPUT0), .B(G543), .Z(n617) );
  NAND2_X1 U564 ( .A1(n635), .A2(G52), .ZN(n518) );
  XNOR2_X1 U565 ( .A(n518), .B(KEYINPUT68), .ZN(n522) );
  INV_X1 U566 ( .A(G651), .ZN(n523) );
  NOR2_X1 U567 ( .A1(G543), .A2(n523), .ZN(n519) );
  XOR2_X1 U568 ( .A(KEYINPUT1), .B(n519), .Z(n634) );
  NAND2_X1 U569 ( .A1(G64), .A2(n634), .ZN(n520) );
  XOR2_X1 U570 ( .A(KEYINPUT67), .B(n520), .Z(n521) );
  NAND2_X1 U571 ( .A1(n522), .A2(n521), .ZN(n530) );
  XNOR2_X1 U572 ( .A(KEYINPUT9), .B(KEYINPUT70), .ZN(n528) );
  NOR2_X1 U573 ( .A1(n617), .A2(n523), .ZN(n643) );
  NAND2_X1 U574 ( .A1(n643), .A2(G77), .ZN(n526) );
  NAND2_X1 U575 ( .A1(n639), .A2(G90), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT69), .B(n524), .Z(n525) );
  NAND2_X1 U577 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U578 ( .A(n528), .B(n527), .Z(n529) );
  NOR2_X1 U579 ( .A1(n530), .A2(n529), .ZN(G171) );
  INV_X1 U580 ( .A(G171), .ZN(G301) );
  NAND2_X1 U581 ( .A1(G89), .A2(n639), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n531), .B(KEYINPUT4), .ZN(n532) );
  XNOR2_X1 U583 ( .A(n532), .B(KEYINPUT80), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G76), .A2(n643), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT5), .ZN(n540) );
  NAND2_X1 U587 ( .A1(G63), .A2(n634), .ZN(n537) );
  NAND2_X1 U588 ( .A1(G51), .A2(n635), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U590 ( .A(KEYINPUT6), .B(n538), .Z(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n541), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U593 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U594 ( .A(G2104), .B(KEYINPUT64), .Z(n546) );
  NAND2_X1 U595 ( .A1(G101), .A2(n595), .ZN(n542) );
  XOR2_X1 U596 ( .A(KEYINPUT23), .B(n542), .Z(n545) );
  NOR2_X1 U597 ( .A1(G2105), .A2(G2104), .ZN(n543) );
  NAND2_X1 U598 ( .A1(n880), .A2(G137), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n545), .A2(n544), .ZN(n685) );
  AND2_X1 U600 ( .A1(G2105), .A2(n546), .ZN(n888) );
  NAND2_X1 U601 ( .A1(G125), .A2(n888), .ZN(n548) );
  AND2_X1 U602 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U603 ( .A1(G113), .A2(n885), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n683) );
  NOR2_X1 U605 ( .A1(n685), .A2(n683), .ZN(G160) );
  XOR2_X1 U606 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n550) );
  NAND2_X1 U607 ( .A1(G7), .A2(G661), .ZN(n549) );
  XNOR2_X1 U608 ( .A(n550), .B(n549), .ZN(G223) );
  INV_X1 U609 ( .A(G223), .ZN(n826) );
  NAND2_X1 U610 ( .A1(n826), .A2(G567), .ZN(n551) );
  XOR2_X1 U611 ( .A(KEYINPUT11), .B(n551), .Z(G234) );
  XOR2_X1 U612 ( .A(KEYINPUT76), .B(KEYINPUT14), .Z(n553) );
  NAND2_X1 U613 ( .A1(G56), .A2(n634), .ZN(n552) );
  XNOR2_X1 U614 ( .A(n553), .B(n552), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n643), .A2(G68), .ZN(n554) );
  XNOR2_X1 U616 ( .A(KEYINPUT78), .B(n554), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT77), .B(KEYINPUT12), .Z(n556) );
  NAND2_X1 U618 ( .A1(G81), .A2(n639), .ZN(n555) );
  XNOR2_X1 U619 ( .A(n556), .B(n555), .ZN(n557) );
  NAND2_X1 U620 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT13), .B(n559), .Z(n560) );
  NOR2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n635), .A2(G43), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n562), .ZN(n707) );
  INV_X1 U625 ( .A(n707), .ZN(n966) );
  XOR2_X1 U626 ( .A(G860), .B(KEYINPUT79), .Z(n584) );
  NAND2_X1 U627 ( .A1(n966), .A2(n584), .ZN(G153) );
  NAND2_X1 U628 ( .A1(G868), .A2(G301), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G92), .A2(n639), .ZN(n565) );
  NAND2_X1 U630 ( .A1(G54), .A2(n635), .ZN(n564) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G79), .A2(n643), .ZN(n567) );
  NAND2_X1 U633 ( .A1(G66), .A2(n634), .ZN(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT15), .ZN(n969) );
  INV_X1 U637 ( .A(G868), .ZN(n654) );
  NAND2_X1 U638 ( .A1(n969), .A2(n654), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(G284) );
  NAND2_X1 U640 ( .A1(G65), .A2(n634), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G53), .A2(n635), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n581) );
  NAND2_X1 U643 ( .A1(n639), .A2(G91), .ZN(n575) );
  XNOR2_X1 U644 ( .A(KEYINPUT71), .B(n575), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n643), .A2(G78), .ZN(n576) );
  XOR2_X1 U646 ( .A(KEYINPUT72), .B(n576), .Z(n577) );
  NOR2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U648 ( .A(n579), .B(KEYINPUT73), .ZN(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n965) );
  XOR2_X1 U650 ( .A(n965), .B(KEYINPUT74), .Z(G299) );
  NOR2_X1 U651 ( .A1(G299), .A2(G868), .ZN(n583) );
  NOR2_X1 U652 ( .A1(G286), .A2(n654), .ZN(n582) );
  NOR2_X1 U653 ( .A1(n583), .A2(n582), .ZN(G297) );
  INV_X1 U654 ( .A(G559), .ZN(n602) );
  NOR2_X1 U655 ( .A1(n584), .A2(n602), .ZN(n585) );
  NOR2_X1 U656 ( .A1(n969), .A2(n585), .ZN(n586) );
  XOR2_X1 U657 ( .A(KEYINPUT16), .B(n586), .Z(G148) );
  NOR2_X1 U658 ( .A1(n969), .A2(n654), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT81), .ZN(n588) );
  NOR2_X1 U660 ( .A1(G559), .A2(n588), .ZN(n590) );
  NOR2_X1 U661 ( .A1(G868), .A2(n707), .ZN(n589) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(G282) );
  XNOR2_X1 U663 ( .A(G2100), .B(KEYINPUT83), .ZN(n601) );
  NAND2_X1 U664 ( .A1(G123), .A2(n888), .ZN(n591) );
  XNOR2_X1 U665 ( .A(n591), .B(KEYINPUT18), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT82), .ZN(n594) );
  NAND2_X1 U667 ( .A1(G111), .A2(n885), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n599) );
  NAND2_X1 U669 ( .A1(G135), .A2(n880), .ZN(n597) );
  NAND2_X1 U670 ( .A1(G99), .A2(n595), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n920) );
  XNOR2_X1 U673 ( .A(n920), .B(G2096), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(G156) );
  OR2_X1 U675 ( .A1(n602), .A2(n969), .ZN(n603) );
  XNOR2_X1 U676 ( .A(n603), .B(n707), .ZN(n652) );
  NOR2_X1 U677 ( .A1(n652), .A2(G860), .ZN(n612) );
  NAND2_X1 U678 ( .A1(G80), .A2(n643), .ZN(n605) );
  NAND2_X1 U679 ( .A1(G67), .A2(n634), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n605), .A2(n604), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G93), .A2(n639), .ZN(n606) );
  XNOR2_X1 U682 ( .A(KEYINPUT85), .B(n606), .ZN(n607) );
  NOR2_X1 U683 ( .A1(n608), .A2(n607), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n635), .A2(G55), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n610), .A2(n609), .ZN(n655) );
  XOR2_X1 U686 ( .A(n655), .B(KEYINPUT84), .Z(n611) );
  XNOR2_X1 U687 ( .A(n612), .B(n611), .ZN(G145) );
  NAND2_X1 U688 ( .A1(G49), .A2(n635), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G74), .A2(G651), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U691 ( .A1(n634), .A2(n615), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT86), .ZN(n619) );
  NAND2_X1 U693 ( .A1(G87), .A2(n617), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n619), .A2(n618), .ZN(G288) );
  NAND2_X1 U695 ( .A1(G75), .A2(n643), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G88), .A2(n639), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G62), .A2(n634), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G50), .A2(n635), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U701 ( .A1(n625), .A2(n624), .ZN(G166) );
  NAND2_X1 U702 ( .A1(G61), .A2(n634), .ZN(n627) );
  NAND2_X1 U703 ( .A1(G48), .A2(n635), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n631) );
  XOR2_X1 U705 ( .A(KEYINPUT2), .B(KEYINPUT87), .Z(n629) );
  NAND2_X1 U706 ( .A1(n643), .A2(G73), .ZN(n628) );
  XOR2_X1 U707 ( .A(n629), .B(n628), .Z(n630) );
  NOR2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n639), .A2(G86), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(G305) );
  NAND2_X1 U711 ( .A1(G60), .A2(n634), .ZN(n637) );
  NAND2_X1 U712 ( .A1(G47), .A2(n635), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U714 ( .A(KEYINPUT66), .B(n638), .ZN(n642) );
  NAND2_X1 U715 ( .A1(G85), .A2(n639), .ZN(n640) );
  XNOR2_X1 U716 ( .A(KEYINPUT65), .B(n640), .ZN(n641) );
  NOR2_X1 U717 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U718 ( .A1(n643), .A2(G72), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(G290) );
  XNOR2_X1 U720 ( .A(G299), .B(KEYINPUT19), .ZN(n647) );
  XNOR2_X1 U721 ( .A(G288), .B(G166), .ZN(n646) );
  XNOR2_X1 U722 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n648), .B(G305), .ZN(n649) );
  XNOR2_X1 U724 ( .A(n649), .B(n655), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n650), .B(G290), .ZN(n896) );
  XNOR2_X1 U726 ( .A(n896), .B(KEYINPUT88), .ZN(n651) );
  XNOR2_X1 U727 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n653), .A2(G868), .ZN(n657) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(KEYINPUT20), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(KEYINPUT89), .ZN(n660) );
  NAND2_X1 U734 ( .A1(n660), .A2(G2090), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(KEYINPUT90), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(KEYINPUT21), .ZN(n663) );
  NAND2_X1 U737 ( .A1(n663), .A2(G2072), .ZN(G158) );
  XOR2_X1 U738 ( .A(KEYINPUT91), .B(G44), .Z(n664) );
  XNOR2_X1 U739 ( .A(KEYINPUT3), .B(n664), .ZN(G218) );
  NOR2_X1 U740 ( .A1(G236), .A2(G238), .ZN(n665) );
  NAND2_X1 U741 ( .A1(G69), .A2(n665), .ZN(n666) );
  NOR2_X1 U742 ( .A1(n666), .A2(G237), .ZN(n667) );
  XNOR2_X1 U743 ( .A(n667), .B(KEYINPUT93), .ZN(n831) );
  NAND2_X1 U744 ( .A1(n831), .A2(G567), .ZN(n673) );
  NAND2_X1 U745 ( .A1(G132), .A2(G82), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n668), .B(KEYINPUT22), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT92), .ZN(n670) );
  NOR2_X1 U748 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U749 ( .A1(G96), .A2(n671), .ZN(n832) );
  NAND2_X1 U750 ( .A1(n832), .A2(G2106), .ZN(n672) );
  NAND2_X1 U751 ( .A1(n673), .A2(n672), .ZN(n833) );
  NAND2_X1 U752 ( .A1(G661), .A2(G483), .ZN(n674) );
  XNOR2_X1 U753 ( .A(KEYINPUT94), .B(n674), .ZN(n675) );
  NOR2_X1 U754 ( .A1(n833), .A2(n675), .ZN(n830) );
  NAND2_X1 U755 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U756 ( .A1(G126), .A2(n888), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G138), .A2(n880), .ZN(n676) );
  NAND2_X1 U758 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U759 ( .A1(G114), .A2(n885), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G102), .A2(n595), .ZN(n678) );
  NAND2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U762 ( .A1(n681), .A2(n680), .ZN(G164) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U764 ( .A(G1986), .B(G290), .ZN(n973) );
  NOR2_X1 U765 ( .A1(G164), .A2(G1384), .ZN(n701) );
  INV_X1 U766 ( .A(G40), .ZN(n682) );
  OR2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n684) );
  OR2_X1 U768 ( .A1(n685), .A2(n684), .ZN(n698) );
  NOR2_X1 U769 ( .A1(n701), .A2(n698), .ZN(n686) );
  XNOR2_X1 U770 ( .A(KEYINPUT95), .B(n686), .ZN(n804) );
  INV_X1 U771 ( .A(n804), .ZN(n820) );
  NAND2_X1 U772 ( .A1(n973), .A2(n820), .ZN(n810) );
  XNOR2_X1 U773 ( .A(G2067), .B(KEYINPUT37), .ZN(n687) );
  XNOR2_X1 U774 ( .A(n687), .B(KEYINPUT96), .ZN(n818) );
  NAND2_X1 U775 ( .A1(G140), .A2(n880), .ZN(n689) );
  NAND2_X1 U776 ( .A1(G104), .A2(n595), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n691) );
  XOR2_X1 U778 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n690) );
  XNOR2_X1 U779 ( .A(n691), .B(n690), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G128), .A2(n888), .ZN(n693) );
  NAND2_X1 U781 ( .A1(G116), .A2(n885), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U783 ( .A(KEYINPUT35), .B(n694), .Z(n695) );
  NOR2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U785 ( .A(KEYINPUT36), .B(n697), .ZN(n859) );
  NOR2_X1 U786 ( .A1(n818), .A2(n859), .ZN(n918) );
  NAND2_X1 U787 ( .A1(n820), .A2(n918), .ZN(n816) );
  INV_X1 U788 ( .A(n816), .ZN(n808) );
  XOR2_X1 U789 ( .A(n698), .B(KEYINPUT100), .Z(n700) );
  NAND2_X1 U790 ( .A1(n701), .A2(n700), .ZN(n749) );
  NOR2_X1 U791 ( .A1(G2084), .A2(n749), .ZN(n699) );
  XOR2_X1 U792 ( .A(KEYINPUT101), .B(n699), .Z(n734) );
  NAND2_X1 U793 ( .A1(n734), .A2(G8), .ZN(n746) );
  NAND2_X1 U794 ( .A1(G8), .A2(n749), .ZN(n776) );
  NOR2_X1 U795 ( .A1(G1966), .A2(n776), .ZN(n744) );
  AND2_X2 U796 ( .A1(n701), .A2(n700), .ZN(n726) );
  NAND2_X1 U797 ( .A1(n726), .A2(G1996), .ZN(n702) );
  XNOR2_X1 U798 ( .A(n702), .B(KEYINPUT26), .ZN(n704) );
  NAND2_X1 U799 ( .A1(G1341), .A2(n749), .ZN(n703) );
  NAND2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U801 ( .A(KEYINPUT104), .B(n705), .Z(n708) );
  NAND2_X1 U802 ( .A1(n966), .A2(n708), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n706), .A2(n969), .ZN(n715) );
  NOR2_X1 U804 ( .A1(n707), .A2(n969), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n709), .A2(n708), .ZN(n713) );
  NOR2_X1 U806 ( .A1(n726), .A2(G1348), .ZN(n711) );
  NOR2_X1 U807 ( .A1(G2067), .A2(n749), .ZN(n710) );
  NOR2_X1 U808 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U810 ( .A1(n715), .A2(n714), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n726), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n716), .B(KEYINPUT27), .ZN(n718) );
  XNOR2_X1 U813 ( .A(G1956), .B(KEYINPUT103), .ZN(n998) );
  NOR2_X1 U814 ( .A1(n998), .A2(n726), .ZN(n717) );
  NOR2_X1 U815 ( .A1(n718), .A2(n717), .ZN(n721) );
  NAND2_X1 U816 ( .A1(n965), .A2(n721), .ZN(n719) );
  NAND2_X1 U817 ( .A1(n720), .A2(n719), .ZN(n724) );
  NOR2_X1 U818 ( .A1(n965), .A2(n721), .ZN(n722) );
  XOR2_X1 U819 ( .A(n722), .B(KEYINPUT28), .Z(n723) );
  NAND2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U821 ( .A(n725), .B(KEYINPUT29), .ZN(n731) );
  NAND2_X1 U822 ( .A1(G1961), .A2(n749), .ZN(n728) );
  XOR2_X1 U823 ( .A(KEYINPUT25), .B(G2078), .Z(n941) );
  NAND2_X1 U824 ( .A1(n726), .A2(n941), .ZN(n727) );
  NAND2_X1 U825 ( .A1(n728), .A2(n727), .ZN(n732) );
  NOR2_X1 U826 ( .A1(G301), .A2(n732), .ZN(n729) );
  XNOR2_X1 U827 ( .A(n729), .B(KEYINPUT102), .ZN(n730) );
  NOR2_X1 U828 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X1 U829 ( .A1(G301), .A2(n732), .ZN(n733) );
  XNOR2_X1 U830 ( .A(n733), .B(KEYINPUT105), .ZN(n739) );
  NOR2_X1 U831 ( .A1(n744), .A2(n734), .ZN(n735) );
  NAND2_X1 U832 ( .A1(G8), .A2(n735), .ZN(n736) );
  XNOR2_X1 U833 ( .A(KEYINPUT30), .B(n736), .ZN(n737) );
  NOR2_X1 U834 ( .A1(n737), .A2(G168), .ZN(n738) );
  NOR2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U836 ( .A(n740), .B(KEYINPUT31), .ZN(n741) );
  INV_X1 U837 ( .A(n747), .ZN(n743) );
  NOR2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U839 ( .A1(n746), .A2(n745), .ZN(n773) );
  NAND2_X1 U840 ( .A1(n747), .A2(G286), .ZN(n756) );
  INV_X1 U841 ( .A(G8), .ZN(n754) );
  NOR2_X1 U842 ( .A1(G1971), .A2(n776), .ZN(n748) );
  XNOR2_X1 U843 ( .A(n748), .B(KEYINPUT106), .ZN(n751) );
  NOR2_X1 U844 ( .A1(n749), .A2(G2090), .ZN(n750) );
  NOR2_X1 U845 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U846 ( .A1(n752), .A2(G303), .ZN(n753) );
  OR2_X1 U847 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n759) );
  XOR2_X1 U849 ( .A(KEYINPUT32), .B(KEYINPUT108), .Z(n757) );
  NAND2_X1 U850 ( .A1(n773), .A2(n775), .ZN(n761) );
  NOR2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n765) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n760) );
  NOR2_X1 U853 ( .A1(n765), .A2(n760), .ZN(n975) );
  NAND2_X1 U854 ( .A1(n761), .A2(n975), .ZN(n762) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n974) );
  NAND2_X1 U856 ( .A1(n762), .A2(n974), .ZN(n763) );
  NOR2_X1 U857 ( .A1(n763), .A2(n776), .ZN(n764) );
  OR2_X1 U858 ( .A1(n764), .A2(KEYINPUT33), .ZN(n770) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n981) );
  INV_X1 U860 ( .A(n981), .ZN(n768) );
  NAND2_X1 U861 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  NOR2_X1 U862 ( .A1(n776), .A2(n766), .ZN(n767) );
  NOR2_X1 U863 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U864 ( .A1(n770), .A2(n769), .ZN(n787) );
  NOR2_X1 U865 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XOR2_X1 U866 ( .A(n771), .B(KEYINPUT24), .Z(n772) );
  NOR2_X1 U867 ( .A1(n776), .A2(n772), .ZN(n785) );
  AND2_X1 U868 ( .A1(n773), .A2(n776), .ZN(n774) );
  NAND2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n782) );
  INV_X1 U870 ( .A(n776), .ZN(n780) );
  NOR2_X1 U871 ( .A1(G2090), .A2(G303), .ZN(n777) );
  XOR2_X1 U872 ( .A(KEYINPUT109), .B(n777), .Z(n778) );
  NAND2_X1 U873 ( .A1(G8), .A2(n778), .ZN(n779) );
  OR2_X1 U874 ( .A1(n780), .A2(n779), .ZN(n781) );
  AND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U876 ( .A(n783), .B(KEYINPUT110), .Z(n784) );
  NOR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n806) );
  NAND2_X1 U879 ( .A1(G119), .A2(n888), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G131), .A2(n880), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n792) );
  NAND2_X1 U882 ( .A1(n885), .A2(G107), .ZN(n790) );
  XOR2_X1 U883 ( .A(KEYINPUT98), .B(n790), .Z(n791) );
  NOR2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n595), .A2(G95), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n862) );
  XOR2_X1 U887 ( .A(KEYINPUT99), .B(G1991), .Z(n942) );
  AND2_X1 U888 ( .A1(n862), .A2(n942), .ZN(n803) );
  NAND2_X1 U889 ( .A1(G141), .A2(n880), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G117), .A2(n885), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n595), .A2(G105), .ZN(n797) );
  XOR2_X1 U893 ( .A(KEYINPUT38), .B(n797), .Z(n798) );
  NOR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n888), .A2(G129), .ZN(n800) );
  NAND2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n863) );
  AND2_X1 U897 ( .A1(n863), .A2(G1996), .ZN(n802) );
  NOR2_X1 U898 ( .A1(n803), .A2(n802), .ZN(n922) );
  NOR2_X1 U899 ( .A1(n922), .A2(n804), .ZN(n813) );
  INV_X1 U900 ( .A(n813), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n823) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n863), .ZN(n932) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n942), .A2(n862), .ZN(n924) );
  NOR2_X1 U907 ( .A1(n811), .A2(n924), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n932), .A2(n814), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n818), .A2(n859), .ZN(n916) );
  NAND2_X1 U913 ( .A1(n819), .A2(n916), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n825) );
  XOR2_X1 U916 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n824) );
  XNOR2_X1 U917 ( .A(n825), .B(n824), .ZN(G329) );
  NAND2_X1 U918 ( .A1(G2106), .A2(n826), .ZN(G217) );
  NAND2_X1 U919 ( .A1(G15), .A2(G2), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT112), .B(n827), .Z(n828) );
  NAND2_X1 U921 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U925 ( .A(G132), .ZN(G219) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n833), .ZN(G319) );
  XOR2_X1 U930 ( .A(G2096), .B(G2100), .Z(n835) );
  XNOR2_X1 U931 ( .A(KEYINPUT42), .B(G2678), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U933 ( .A(KEYINPUT43), .B(G2072), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2090), .B(G2067), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1986), .B(G1971), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1981), .B(G1976), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U942 ( .A(G1991), .B(G1966), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1956), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U946 ( .A(KEYINPUT113), .B(G2474), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U948 ( .A(G1961), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G136), .A2(n880), .ZN(n853) );
  NAND2_X1 U951 ( .A1(G112), .A2(n885), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U953 ( .A1(n888), .A2(G124), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U955 ( .A1(G100), .A2(n595), .ZN(n855) );
  NAND2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U957 ( .A1(n858), .A2(n857), .ZN(G162) );
  XNOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n859), .B(KEYINPUT119), .ZN(n860) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n867) );
  XNOR2_X1 U961 ( .A(n920), .B(n862), .ZN(n865) );
  XOR2_X1 U962 ( .A(G160), .B(n863), .Z(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U964 ( .A(n867), .B(n866), .Z(n869) );
  XNOR2_X1 U965 ( .A(G164), .B(G162), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n869), .B(n868), .ZN(n894) );
  NAND2_X1 U967 ( .A1(n880), .A2(G139), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n870), .B(KEYINPUT116), .ZN(n872) );
  NAND2_X1 U969 ( .A1(G103), .A2(n595), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U971 ( .A(n873), .B(KEYINPUT117), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G127), .A2(n888), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G115), .A2(n885), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U975 ( .A(KEYINPUT47), .B(n876), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(KEYINPUT118), .ZN(n927) );
  NAND2_X1 U978 ( .A1(n880), .A2(G142), .ZN(n881) );
  XOR2_X1 U979 ( .A(KEYINPUT115), .B(n881), .Z(n883) );
  NAND2_X1 U980 ( .A1(n595), .A2(G106), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(KEYINPUT45), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G118), .A2(n885), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n891) );
  NAND2_X1 U985 ( .A1(n888), .A2(G130), .ZN(n889) );
  XOR2_X1 U986 ( .A(KEYINPUT114), .B(n889), .Z(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n927), .B(n892), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U990 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U991 ( .A(n969), .B(n896), .ZN(n898) );
  XNOR2_X1 U992 ( .A(G286), .B(n966), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(G301), .ZN(n900) );
  NOR2_X1 U995 ( .A1(G37), .A2(n900), .ZN(G397) );
  XOR2_X1 U996 ( .A(G2451), .B(G2430), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2438), .B(G2443), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n908) );
  XOR2_X1 U999 ( .A(G2435), .B(G2454), .Z(n904) );
  XNOR2_X1 U1000 ( .A(G1348), .B(G1341), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n906) );
  XOR2_X1 U1002 ( .A(G2446), .B(G2427), .Z(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1004 ( .A(n908), .B(n907), .Z(n909) );
  NAND2_X1 U1005 ( .A1(G14), .A2(n909), .ZN(n915) );
  NAND2_X1 U1006 ( .A1(G319), .A2(n915), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G69), .ZN(G235) );
  INV_X1 U1015 ( .A(n915), .ZN(G401) );
  INV_X1 U1016 ( .A(n916), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n926) );
  XOR2_X1 U1018 ( .A(G2084), .B(G160), .Z(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n937) );
  XOR2_X1 U1023 ( .A(G164), .B(G2078), .Z(n929) );
  XNOR2_X1 U1024 ( .A(G2072), .B(n927), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n930), .ZN(n935) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1029 ( .A(KEYINPUT51), .B(n933), .Z(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n938), .ZN(n939) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n961) );
  NAND2_X1 U1034 ( .A1(n939), .A2(n961), .ZN(n940) );
  NAND2_X1 U1035 ( .A1(n940), .A2(G29), .ZN(n1023) );
  XOR2_X1 U1036 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n954) );
  XNOR2_X1 U1037 ( .A(n941), .B(G27), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(n942), .B(G25), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(G2067), .B(G26), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G1996), .B(G32), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1043 ( .A1(G28), .A2(n947), .ZN(n950) );
  XNOR2_X1 U1044 ( .A(G33), .B(G2072), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT120), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n954), .B(n953), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G2084), .B(G34), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT54), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G35), .B(G2090), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1054 ( .A(n961), .B(n960), .ZN(n963) );
  INV_X1 U1055 ( .A(G29), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n964), .ZN(n1021) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XOR2_X1 U1059 ( .A(n965), .B(G1956), .Z(n968) );
  XOR2_X1 U1060 ( .A(n966), .B(G1341), .Z(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n988) );
  XNOR2_X1 U1062 ( .A(G171), .B(G1961), .ZN(n971) );
  XOR2_X1 U1063 ( .A(G1348), .B(n969), .Z(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n980) );
  NAND2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n977) );
  AND2_X1 U1067 ( .A1(G303), .A2(G1971), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XOR2_X1 U1069 ( .A(KEYINPUT123), .B(n978), .Z(n979) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n986) );
  XNOR2_X1 U1071 ( .A(G168), .B(G1966), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n983), .B(KEYINPUT57), .ZN(n984) );
  XOR2_X1 U1074 ( .A(KEYINPUT122), .B(n984), .Z(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1076 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1077 ( .A1(n990), .A2(n989), .ZN(n1019) );
  INV_X1 U1078 ( .A(G16), .ZN(n1017) );
  XOR2_X1 U1079 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n997) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n992) );
  XNOR2_X1 U1081 ( .A(G24), .B(G1986), .ZN(n991) );
  NOR2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n995) );
  XOR2_X1 U1083 ( .A(G1976), .B(KEYINPUT126), .Z(n993) );
  XNOR2_X1 U1084 ( .A(G23), .B(n993), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(n997), .B(n996), .ZN(n1014) );
  XOR2_X1 U1087 ( .A(G1961), .B(G5), .Z(n1009) );
  XOR2_X1 U1088 ( .A(G1981), .B(G6), .Z(n1000) );
  XNOR2_X1 U1089 ( .A(n998), .B(G20), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(n1001), .B(G4), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(G1341), .B(KEYINPUT124), .Z(n1002) );
  XNOR2_X1 U1094 ( .A(G19), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G21), .B(G1966), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT125), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(KEYINPUT61), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1024), .Z(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

