//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(new_n203), .A2(G50), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G1), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n209), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT0), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT65), .Z(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT66), .ZN(new_n225));
  OR2_X1    g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT64), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n226), .A2(new_n227), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(new_n214), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n211), .B(new_n217), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NOR2_X1   g0050(.A1(new_n209), .A2(G1), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT70), .ZN(new_n252));
  INV_X1    g0052(.A(G50), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n212), .A2(G13), .A3(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n208), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n254), .A2(new_n259), .B1(new_n253), .B2(new_n256), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n209), .A2(G33), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g0063(.A(KEYINPUT8), .B(G58), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n258), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n260), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  AND2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT68), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n273), .B1(new_n276), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n276), .A2(new_n282), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(G222), .A3(new_n273), .ZN(new_n286));
  INV_X1    g0086(.A(G77), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n284), .B(new_n286), .C1(new_n287), .C2(new_n285), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n208), .B1(G33), .B2(G41), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(G1), .A3(G13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n295), .A3(G274), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n289), .A2(new_n293), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(G226), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n290), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n272), .B1(new_n301), .B2(G169), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n300), .A2(G179), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n272), .B(KEYINPUT9), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n301), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G190), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n307), .A2(KEYINPUT10), .A3(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n304), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n298), .ZN(new_n313));
  INV_X1    g0113(.A(G244), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n296), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n285), .A2(G232), .A3(new_n273), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n285), .A2(G238), .A3(G1698), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n276), .A2(new_n282), .A3(G107), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n315), .B1(new_n319), .B2(new_n289), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G190), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n252), .A2(new_n287), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(new_n259), .B1(new_n287), .B2(new_n256), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n264), .A2(new_n269), .B1(new_n209), .B2(new_n287), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(new_n261), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n258), .B1(new_n324), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n321), .B(new_n329), .C1(new_n306), .C2(new_n320), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n328), .B1(new_n320), .B2(G169), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT71), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n320), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(KEYINPUT71), .B(new_n328), .C1(new_n320), .C2(G169), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n312), .A2(new_n330), .A3(new_n337), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n263), .A2(new_n287), .B1(new_n209), .B2(G68), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n268), .A2(G50), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT74), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n342), .B1(new_n209), .B2(G68), .C1(new_n263), .C2(new_n287), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n258), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT11), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n252), .A2(new_n202), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT12), .B1(new_n255), .B2(G68), .ZN(new_n350));
  OR3_X1    g0150(.A1(new_n255), .A2(KEYINPUT12), .A3(G68), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n349), .A2(new_n259), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT14), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n283), .B2(G232), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n285), .A2(G226), .A3(new_n273), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n295), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(G238), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n296), .B1(new_n313), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(KEYINPUT13), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n274), .A2(new_n275), .A3(KEYINPUT68), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n364));
  OAI211_X1 g0164(.A(G232), .B(G1698), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n358), .A2(new_n365), .A3(new_n355), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n289), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT13), .ZN(new_n368));
  INV_X1    g0168(.A(new_n361), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n367), .A2(KEYINPUT72), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n362), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n361), .B1(new_n366), .B2(new_n289), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT72), .B1(new_n372), .B2(new_n368), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n354), .B(G169), .C1(new_n371), .C2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT73), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n377), .A3(new_n368), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n376), .A2(G179), .A3(new_n362), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n375), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n382), .A2(new_n362), .A3(new_n370), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n354), .B1(new_n383), .B2(G169), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n353), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(G200), .B1(new_n371), .B2(new_n373), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n348), .A2(new_n352), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT11), .B1(new_n344), .B2(new_n258), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n376), .A2(G190), .A3(new_n362), .A4(new_n378), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n385), .A2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n252), .A2(new_n264), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n259), .B1(new_n256), .B2(new_n264), .ZN(new_n394));
  XNOR2_X1  g0194(.A(G58), .B(G68), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n268), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT75), .B(G33), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n275), .B1(new_n398), .B2(KEYINPUT3), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n397), .B1(new_n399), .B2(new_n209), .ZN(new_n400));
  AND2_X1   g0200(.A1(KEYINPUT75), .A2(G33), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT75), .A2(G33), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT3), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n403), .A2(new_n397), .A3(new_n209), .A4(new_n279), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G68), .ZN(new_n405));
  OAI211_X1 g0205(.A(KEYINPUT16), .B(new_n396), .C1(new_n400), .C2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n258), .ZN(new_n407));
  XNOR2_X1  g0207(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n276), .A2(new_n282), .A3(new_n397), .A4(new_n209), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n281), .A2(new_n209), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n401), .A2(new_n402), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n277), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n410), .B(G68), .C1(new_n397), .C2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n409), .B1(new_n414), .B2(new_n396), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n394), .B1(new_n407), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g0216(.A1(G223), .A2(G1698), .ZN(new_n417));
  INV_X1    g0217(.A(G226), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G1698), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n403), .B2(new_n279), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n278), .A2(new_n220), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n289), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT77), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n298), .A2(G232), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n425), .A2(new_n334), .A3(new_n296), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n289), .C1(new_n421), .C2(new_n422), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(G169), .ZN(new_n430));
  INV_X1    g0230(.A(new_n423), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n425), .A2(new_n296), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n416), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT18), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT18), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n416), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n425), .A2(new_n308), .A3(new_n296), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n424), .A2(new_n440), .A3(new_n428), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n306), .B1(new_n431), .B2(new_n432), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n439), .B1(new_n416), .B2(new_n443), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n414), .A2(new_n396), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n258), .B(new_n406), .C1(new_n445), .C2(new_n409), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n441), .A2(new_n442), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(KEYINPUT17), .A4(new_n394), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n436), .A2(new_n438), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  AND3_X1   g0250(.A1(new_n338), .A2(new_n392), .A3(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT4), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(new_n314), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n273), .B(new_n455), .C1(new_n363), .C2(new_n364), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n273), .A2(G244), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n403), .B2(new_n279), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n460), .B2(KEYINPUT4), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n289), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT5), .B(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n292), .A2(G1), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(G274), .A3(new_n295), .A4(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n289), .B1(new_n464), .B2(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G257), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n462), .A2(G190), .A3(new_n465), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT78), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n454), .B1(new_n399), .B2(new_n459), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n470), .A2(new_n453), .A3(new_n458), .A4(new_n456), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(new_n289), .B1(G257), .B2(new_n466), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT78), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n472), .A2(new_n473), .A3(G190), .A4(new_n465), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  INV_X1    g0276(.A(G107), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n222), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n268), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n410), .B1(new_n397), .B2(new_n413), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n477), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n258), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n256), .A2(new_n222), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n212), .A2(G33), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n255), .A2(new_n488), .A3(new_n208), .A4(new_n257), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(new_n222), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n462), .A2(new_n465), .A3(new_n467), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(G200), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n472), .A2(new_n334), .A3(new_n465), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n493), .A2(new_n430), .B1(new_n486), .B2(new_n491), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n475), .A2(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT84), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n221), .A2(new_n273), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n223), .A2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n501), .B1(new_n403), .B2(new_n279), .ZN(new_n502));
  INV_X1    g0302(.A(G294), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n412), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n498), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n398), .A2(G294), .ZN(new_n506));
  OAI211_X1 g0306(.A(KEYINPUT84), .B(new_n506), .C1(new_n399), .C2(new_n501), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n507), .A3(new_n289), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n466), .A2(G264), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n508), .A2(new_n465), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n306), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT85), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT85), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n510), .A2(new_n513), .A3(new_n306), .ZN(new_n514));
  INV_X1    g0314(.A(new_n510), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n308), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n258), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT75), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n278), .ZN(new_n520));
  NAND2_X1  g0320(.A1(KEYINPUT75), .A2(G33), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n277), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n209), .B(G87), .C1(new_n522), .C2(new_n275), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n220), .A2(KEYINPUT22), .A3(G20), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n523), .A2(KEYINPUT22), .B1(new_n285), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT83), .B1(new_n209), .B2(G107), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  OR2_X1    g0329(.A1(KEYINPUT79), .A2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT79), .A2(G116), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n398), .ZN(new_n533));
  OAI211_X1 g0333(.A(new_n528), .B(new_n529), .C1(new_n533), .C2(G20), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT24), .B1(new_n525), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n534), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT22), .ZN(new_n538));
  AOI21_X1  g0338(.A(G20), .B1(new_n403), .B2(new_n279), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n538), .B1(new_n539), .B2(G87), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n285), .A2(new_n524), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n536), .B(new_n537), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n518), .B1(new_n535), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n477), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT25), .B1(new_n256), .B2(new_n477), .ZN(new_n546));
  OAI22_X1  g0346(.A1(new_n545), .A2(new_n546), .B1(new_n477), .B2(new_n489), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n517), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n497), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n360), .A2(new_n273), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n314), .A2(G1698), .ZN(new_n552));
  AND2_X1   g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n522), .B2(new_n275), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n295), .B1(new_n554), .B2(new_n533), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n295), .B(G250), .C1(G1), .C2(new_n292), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n295), .A2(G274), .A3(new_n464), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT80), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n551), .A2(new_n552), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n560), .B1(new_n403), .B2(new_n279), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n530), .A2(new_n531), .B1(new_n520), .B2(new_n521), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n289), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT80), .ZN(new_n564));
  INV_X1    g0364(.A(new_n558), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n559), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n403), .A2(new_n279), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n209), .A3(G68), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n479), .A2(new_n220), .B1(new_n355), .B2(new_n209), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT19), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G97), .ZN(new_n572));
  OAI22_X1  g0372(.A1(new_n570), .A2(new_n571), .B1(new_n261), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n518), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n325), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n255), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n489), .A2(new_n325), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n567), .A2(new_n334), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n559), .A2(new_n430), .A3(new_n566), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n308), .B1(new_n559), .B2(new_n566), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n489), .A2(new_n220), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n574), .A2(new_n576), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n559), .A2(G200), .A3(new_n566), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n583), .C2(new_n584), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n582), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n510), .A2(new_n430), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n508), .A2(new_n334), .A3(new_n465), .A4(new_n509), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n592), .B(new_n593), .C1(new_n543), .C2(new_n547), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  MUX2_X1   g0395(.A(G257), .B(G264), .S(G1698), .Z(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n522), .B2(new_n275), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n276), .A2(new_n282), .A3(G303), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n295), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(KEYINPUT5), .A2(G41), .ZN(new_n600));
  NOR2_X1   g0400(.A1(KEYINPUT5), .A2(G41), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n464), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(G270), .A3(new_n295), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n465), .ZN(new_n604));
  OAI21_X1  g0404(.A(G169), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  OAI22_X1  g0406(.A1(new_n489), .A2(new_n606), .B1(new_n255), .B2(new_n532), .ZN(new_n607));
  AOI21_X1  g0407(.A(G20), .B1(G33), .B2(G283), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n278), .A2(G97), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n608), .A2(new_n609), .B1(new_n257), .B2(new_n208), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n530), .A2(G20), .A3(new_n531), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n610), .A2(KEYINPUT20), .A3(new_n611), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n607), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n595), .B1(new_n605), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT82), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT82), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n619), .B(new_n595), .C1(new_n605), .C2(new_n616), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n616), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n597), .A2(new_n598), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n289), .ZN(new_n624));
  INV_X1    g0424(.A(new_n604), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n622), .B1(new_n626), .B2(G200), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n308), .B2(new_n626), .ZN(new_n628));
  OAI22_X1  g0428(.A1(new_n334), .A2(new_n626), .B1(new_n605), .B2(new_n595), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n622), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n594), .A2(new_n621), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  NOR4_X1   g0431(.A1(new_n452), .A2(new_n550), .A3(new_n591), .A4(new_n631), .ZN(G372));
  NAND2_X1  g0432(.A1(new_n493), .A2(new_n430), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n633), .A2(new_n495), .A3(new_n492), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n589), .A2(new_n588), .ZN(new_n635));
  AND3_X1   g0435(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n564), .B1(new_n563), .B2(new_n565), .ZN(new_n637));
  OAI21_X1  g0437(.A(G190), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT81), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n635), .A2(new_n585), .A3(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n634), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n582), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT87), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n334), .B1(new_n636), .B2(new_n637), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n577), .A2(new_n579), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n558), .A2(KEYINPUT86), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT86), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n556), .A2(new_n647), .A3(new_n557), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n563), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n430), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n644), .A2(new_n645), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n650), .A2(G200), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n638), .A2(new_n588), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n633), .A2(new_n495), .A3(new_n492), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n643), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n641), .A2(new_n642), .A3(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n652), .B1(new_n641), .B2(new_n642), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT88), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n641), .A2(new_n642), .A3(new_n657), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT88), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n644), .A2(new_n581), .A3(new_n645), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n584), .B1(new_n567), .B2(G190), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n589), .A2(new_n588), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n663), .B1(new_n666), .B2(new_n585), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(KEYINPUT87), .A3(KEYINPUT26), .A4(new_n634), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n661), .A2(new_n662), .A3(new_n668), .A4(new_n652), .ZN(new_n669));
  INV_X1    g0469(.A(new_n655), .ZN(new_n670));
  INV_X1    g0470(.A(new_n594), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n626), .A2(new_n622), .A3(G169), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n619), .B1(new_n672), .B2(new_n595), .ZN(new_n673));
  INV_X1    g0473(.A(new_n620), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n630), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n670), .B1(new_n671), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n550), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n660), .A2(new_n669), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n451), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n310), .A2(new_n311), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n444), .A2(new_n448), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n336), .A2(new_n335), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n391), .A2(new_n333), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n385), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT89), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n416), .A2(new_n434), .A3(new_n437), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n437), .B1(new_n416), .B2(new_n434), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n436), .A2(KEYINPUT89), .A3(new_n438), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n681), .B1(new_n687), .B2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n304), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n680), .A2(new_n697), .ZN(G369));
  NAND3_X1  g0498(.A1(new_n212), .A2(new_n209), .A3(G13), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT27), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G213), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT90), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT91), .B(G343), .Z(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(new_n616), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n675), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n628), .ZN(new_n712));
  INV_X1    g0512(.A(G330), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n535), .A2(new_n542), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n258), .ZN(new_n716));
  INV_X1    g0516(.A(new_n547), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n511), .A2(KEYINPUT85), .B1(new_n515), .B2(new_n308), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n514), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n709), .B1(new_n716), .B2(new_n717), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n594), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n594), .A2(new_n708), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n714), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n675), .A2(new_n709), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n723), .B1(new_n722), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n726), .A2(new_n729), .ZN(G399));
  INV_X1    g0530(.A(new_n215), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G41), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n479), .A2(new_n220), .A3(new_n606), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n206), .B2(new_n733), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n667), .A2(new_n643), .A3(new_n634), .ZN(new_n739));
  INV_X1    g0539(.A(new_n652), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n496), .A2(new_n652), .A3(new_n654), .A4(new_n495), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n740), .B1(new_n741), .B2(KEYINPUT26), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n739), .B(new_n742), .C1(new_n550), .C2(new_n676), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(new_n709), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT29), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n661), .A2(new_n652), .A3(new_n668), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n677), .B1(new_n747), .B2(KEYINPUT88), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n708), .B1(new_n748), .B2(new_n669), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n746), .B1(new_n749), .B2(new_n745), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n631), .A2(new_n591), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n751), .A2(new_n549), .A3(new_n497), .A4(new_n709), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT92), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT30), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n462), .B(new_n467), .C1(new_n636), .C2(new_n637), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n604), .B1(new_n623), .B2(new_n289), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n508), .A2(new_n756), .A3(G179), .A4(new_n509), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n754), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  AND4_X1   g0558(.A1(G179), .A2(new_n508), .A3(new_n756), .A4(new_n509), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(KEYINPUT30), .A3(new_n472), .A4(new_n567), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n756), .A2(G179), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n493), .A2(new_n510), .A3(new_n650), .A4(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n758), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(new_n708), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n753), .B1(new_n764), .B2(KEYINPUT31), .ZN(new_n765));
  AOI21_X1  g0565(.A(KEYINPUT31), .B1(new_n763), .B2(new_n708), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(KEYINPUT92), .ZN(new_n767));
  AND3_X1   g0567(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n708), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n752), .A2(new_n765), .A3(new_n767), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n770), .A2(G330), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n750), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n738), .B1(new_n774), .B2(G1), .ZN(G364));
  AND2_X1   g0575(.A1(new_n209), .A2(G13), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n212), .B1(new_n776), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n732), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(G330), .B1(new_n711), .B2(new_n628), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n714), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n208), .B1(G20), .B2(new_n430), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n209), .A2(new_n334), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G190), .A2(G200), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n209), .A2(G179), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n784), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G311), .A2(new_n786), .B1(new_n789), .B2(G329), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n306), .A2(G190), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n787), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(G322), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n783), .A2(G190), .A3(new_n306), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n790), .B1(new_n791), .B2(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n308), .A2(new_n306), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n783), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(G326), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n797), .A2(new_n787), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n783), .A2(new_n792), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  OAI221_X1 g0604(.A(new_n800), .B1(new_n801), .B2(new_n802), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n285), .ZN(new_n806));
  NOR3_X1   g0606(.A1(new_n308), .A2(G179), .A3(G200), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n209), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n806), .B1(new_n503), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n796), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n811), .A2(new_n788), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n808), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G97), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n811), .B1(new_n788), .B2(new_n812), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n813), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n285), .B1(new_n477), .B2(new_n793), .C1(new_n201), .C2(new_n795), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n202), .A2(new_n803), .B1(new_n802), .B2(new_n220), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n798), .A2(new_n253), .B1(new_n785), .B2(new_n287), .ZN(new_n820));
  NOR4_X1   g0620(.A1(new_n817), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n782), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n782), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n731), .A2(new_n568), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(G45), .B2(new_n206), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G45), .B2(new_n249), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n285), .A2(new_n215), .ZN(new_n830));
  INV_X1    g0630(.A(G355), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n830), .A2(new_n831), .B1(G116), .B2(new_n215), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n826), .B1(new_n829), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g0633(.A(new_n779), .B(KEYINPUT93), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n822), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT95), .Z(new_n836));
  XNOR2_X1  g0636(.A(new_n825), .B(KEYINPUT96), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n712), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n781), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(G396));
  NOR2_X1   g0641(.A1(new_n782), .A2(new_n823), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT97), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n834), .B1(new_n843), .B2(G77), .ZN(new_n844));
  INV_X1    g0644(.A(new_n803), .ZN(new_n845));
  AOI22_X1  g0645(.A1(G137), .A2(new_n799), .B1(new_n845), .B2(G150), .ZN(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n795), .C1(new_n812), .C2(new_n785), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  OR2_X1    g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n849), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n802), .A2(new_n253), .B1(new_n788), .B2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n793), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n853), .B1(G68), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n399), .B1(new_n814), .B2(G58), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n850), .A2(new_n851), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n793), .A2(new_n220), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(G303), .B2(new_n799), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n791), .B2(new_n803), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n802), .A2(new_n477), .ZN(new_n861));
  INV_X1    g0661(.A(new_n532), .ZN(new_n862));
  OAI22_X1  g0662(.A1(new_n862), .A2(new_n785), .B1(new_n795), .B2(new_n503), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(G311), .C2(new_n789), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n864), .A2(new_n806), .A3(new_n815), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n857), .B1(new_n860), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n844), .B1(new_n866), .B2(new_n782), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n709), .A2(new_n329), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n331), .A2(new_n332), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n684), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n869), .B1(new_n337), .B2(new_n868), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n330), .B1(new_n685), .B2(new_n333), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n867), .B1(new_n875), .B2(new_n824), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n679), .A2(new_n709), .ZN(new_n877));
  INV_X1    g0677(.A(new_n875), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n679), .A2(new_n709), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n881), .A2(new_n772), .B1(new_n732), .B2(new_n778), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT99), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(new_n772), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n882), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n876), .B1(new_n884), .B2(new_n886), .ZN(G384));
  OR2_X1    g0687(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(G116), .A3(new_n210), .A4(new_n889), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT36), .Z(new_n891));
  OAI211_X1 g0691(.A(new_n207), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n253), .A2(G68), .ZN(new_n893));
  AOI211_X1 g0693(.A(new_n212), .B(G13), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT38), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT7), .B1(new_n568), .B2(G20), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(G68), .A3(new_n404), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n409), .B1(new_n898), .B2(new_n396), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n394), .B1(new_n407), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n434), .ZN(new_n901));
  INV_X1    g0701(.A(new_n706), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n446), .A2(new_n394), .A3(new_n447), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n706), .B(KEYINPUT101), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n416), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n435), .A4(new_n904), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n689), .A2(new_n690), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n903), .B1(new_n682), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n896), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT102), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n906), .A2(new_n910), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n916), .B(KEYINPUT38), .C1(new_n450), .C2(new_n903), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n914), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(KEYINPUT102), .B(new_n896), .C1(new_n911), .C2(new_n913), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT39), .ZN(new_n921));
  INV_X1    g0721(.A(new_n385), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n709), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n691), .A2(new_n692), .A3(new_n682), .ZN(new_n925));
  INV_X1    g0725(.A(new_n908), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n908), .A2(new_n435), .A3(new_n904), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n925), .A2(new_n926), .B1(new_n910), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n917), .B1(new_n929), .B2(KEYINPUT38), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n921), .A2(new_n924), .A3(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n693), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n934), .A2(new_n907), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT100), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n938), .B(new_n708), .C1(new_n387), .C2(new_n388), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n938), .B1(new_n353), .B2(new_n708), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n385), .A2(new_n391), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(G169), .B1(new_n371), .B2(new_n373), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT14), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n391), .A2(new_n945), .A3(new_n379), .A4(new_n374), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n389), .A2(new_n709), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n337), .A2(new_n708), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n950), .B(new_n920), .C1(new_n880), .C2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n937), .A2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n746), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n877), .B2(KEYINPUT29), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n696), .B1(new_n956), .B2(new_n451), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n954), .B(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT40), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n918), .A2(new_n959), .A3(new_n919), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n768), .A2(new_n766), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n752), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n949), .A2(new_n962), .A3(new_n875), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g0764(.A1(new_n949), .A2(new_n962), .A3(new_n875), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n959), .B1(new_n965), .B2(new_n930), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n451), .A2(new_n962), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(G330), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n958), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n212), .B2(new_n776), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n958), .A2(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n895), .B1(new_n973), .B2(new_n974), .ZN(G367));
  AND2_X1   g0775(.A1(new_n238), .A2(new_n827), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n826), .B1(new_n215), .B2(new_n325), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n834), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n793), .A2(new_n287), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n979), .B1(G50), .B2(new_n786), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n201), .B2(new_n802), .C1(new_n847), .C2(new_n798), .ZN(new_n981));
  INV_X1    g0781(.A(new_n795), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n982), .A2(G150), .B1(new_n845), .B2(G159), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT107), .B(G137), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n983), .B1(new_n788), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n808), .A2(new_n202), .ZN(new_n986));
  NOR4_X1   g0786(.A1(new_n981), .A2(new_n806), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n802), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT46), .B1(new_n988), .B2(new_n532), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n568), .B(new_n989), .C1(G107), .C2(new_n814), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n793), .A2(new_n222), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G303), .B2(new_n982), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n988), .A2(KEYINPUT46), .A3(G116), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n791), .C2(new_n785), .ZN(new_n994));
  XNOR2_X1  g0794(.A(KEYINPUT105), .B(G311), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n799), .A2(new_n996), .B1(new_n845), .B2(G294), .ZN(new_n997));
  XOR2_X1   g0797(.A(KEYINPUT106), .B(G317), .Z(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n788), .B2(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n987), .B1(new_n990), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT47), .Z(new_n1002));
  AOI21_X1  g0802(.A(new_n978), .B1(new_n1002), .B2(new_n782), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n709), .A2(new_n588), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n740), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n655), .B2(new_n1004), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1003), .B1(new_n837), .B2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT108), .Z(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT104), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT103), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n475), .A2(new_n494), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n492), .A2(new_n708), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1012), .A2(new_n656), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n634), .A2(new_n708), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n729), .A2(new_n1011), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n721), .B1(new_n517), .B2(new_n548), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1018), .A2(new_n675), .A3(new_n594), .A4(new_n709), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n1016), .A3(new_n724), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT103), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT45), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT44), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n729), .B2(new_n1016), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1016), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1019), .ZN(new_n1027));
  OAI211_X1 g0827(.A(KEYINPUT44), .B(new_n1026), .C1(new_n1027), .C2(new_n723), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n1022), .A2(new_n1023), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1017), .A2(new_n1021), .A3(KEYINPUT45), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n726), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1011), .B1(new_n729), .B2(new_n1016), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1020), .A2(KEYINPUT103), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1023), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1035));
  AND4_X1   g0835(.A1(new_n726), .A2(new_n1034), .A3(new_n1030), .A4(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n725), .A2(new_n728), .ZN(new_n1038));
  OR3_X1    g0838(.A1(new_n1038), .A2(new_n714), .A3(new_n1027), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n714), .B1(new_n1038), .B2(new_n1027), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n773), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n732), .B(KEYINPUT41), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1010), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1043), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n750), .A2(new_n1041), .A3(new_n772), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1046), .A2(new_n1031), .A3(new_n1036), .ZN(new_n1047));
  OAI211_X1 g0847(.A(KEYINPUT104), .B(new_n1045), .C1(new_n1047), .C2(new_n773), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n778), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1027), .A2(new_n1016), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT42), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n656), .B1(new_n1014), .B2(new_n594), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n709), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1051), .A2(KEYINPUT42), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1050), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1057), .B(new_n1058), .Z(new_n1059));
  NOR2_X1   g0859(.A1(new_n726), .A2(new_n1026), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1059), .B(new_n1060), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1009), .B1(new_n1049), .B2(new_n1061), .ZN(G387));
  NOR2_X1   g0862(.A1(new_n725), .A2(new_n837), .ZN(new_n1063));
  AOI211_X1 g0863(.A(G45), .B(new_n734), .C1(G68), .C2(G77), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n264), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n1065), .A2(KEYINPUT50), .A3(new_n253), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT50), .B1(new_n1065), .B2(new_n253), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(KEYINPUT109), .B1(new_n1068), .B2(new_n827), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(G45), .B2(new_n242), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1068), .A2(KEYINPUT109), .A3(new_n827), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(G107), .B2(new_n215), .C1(new_n735), .C2(new_n830), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n826), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n834), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n798), .A2(new_n812), .B1(new_n802), .B2(new_n287), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n991), .B(new_n1076), .C1(G150), .C2(new_n789), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n795), .A2(new_n253), .B1(new_n785), .B2(new_n202), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n1065), .B2(new_n845), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n814), .A2(new_n575), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n568), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(G322), .A2(new_n799), .B1(new_n845), .B2(new_n996), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n801), .B2(new_n785), .C1(new_n795), .C2(new_n998), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT48), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT110), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n808), .A2(new_n791), .B1(new_n802), .B2(new_n503), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1083), .A2(new_n1084), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1086), .A2(new_n1085), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1087), .B(new_n1088), .C1(new_n1084), .C2(new_n1083), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT111), .Z(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT49), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n532), .A2(new_n854), .B1(new_n789), .B2(G326), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1091), .A2(new_n399), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1090), .A2(KEYINPUT49), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1081), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1063), .B(new_n1075), .C1(new_n1095), .C2(new_n782), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n778), .B2(new_n1041), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n774), .A2(new_n1041), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1046), .A2(new_n732), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  NOR2_X1   g0900(.A1(new_n1047), .A2(new_n733), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1046), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1037), .A2(new_n778), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1026), .A2(new_n825), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT112), .Z(new_n1106));
  AOI22_X1  g0906(.A1(new_n982), .A2(G311), .B1(new_n799), .B2(G317), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT52), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n785), .A2(new_n503), .B1(new_n788), .B2(new_n794), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(G303), .B2(new_n845), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n814), .A2(new_n532), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n802), .A2(new_n791), .B1(new_n793), .B2(new_n477), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1112), .A2(new_n285), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n399), .B(new_n858), .C1(G68), .C2(new_n988), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n803), .A2(new_n253), .B1(new_n788), .B2(new_n847), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n1065), .B2(new_n786), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n814), .A2(G77), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n795), .A2(new_n812), .B1(new_n798), .B2(new_n267), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT51), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n1108), .A2(new_n1114), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n782), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n827), .A2(new_n246), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n1124), .B(new_n826), .C1(new_n222), .C2(new_n215), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n834), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT113), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1106), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1103), .A2(new_n1104), .A3(new_n1128), .ZN(G390));
  AOI21_X1  g0929(.A(new_n713), .B1(new_n752), .B2(new_n961), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n451), .A2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n697), .B(new_n1131), .C1(new_n750), .C2(new_n452), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n770), .A2(G330), .A3(new_n875), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1133), .A2(new_n950), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n875), .A3(new_n949), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n880), .A2(new_n952), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n771), .A2(new_n875), .A3(new_n949), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n949), .B1(new_n1130), .B2(new_n875), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n743), .A2(new_n709), .A3(new_n875), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n952), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1132), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n921), .A2(new_n932), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n950), .B1(new_n880), .B2(new_n952), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n924), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1141), .A2(new_n949), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1149), .A2(new_n923), .A3(new_n930), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n1148), .A2(new_n1151), .A3(new_n1138), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1135), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1145), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1148), .A2(new_n1151), .A3(new_n1138), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n951), .B1(new_n749), .B2(new_n875), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n923), .B1(new_n1156), .B2(new_n950), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1150), .B1(new_n1157), .B2(new_n1146), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1155), .B(new_n1144), .C1(new_n1158), .C2(new_n1135), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1154), .A2(new_n732), .A3(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1155), .B(new_n778), .C1(new_n1158), .C2(new_n1135), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n834), .B1(new_n843), .B2(new_n1065), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n802), .A2(new_n267), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n806), .B1(G159), .B2(new_n814), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(G50), .A2(new_n854), .B1(new_n789), .B2(G125), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n984), .ZN(new_n1167));
  XOR2_X1   g0967(.A(KEYINPUT54), .B(G143), .Z(new_n1168));
  AOI22_X1  g0968(.A1(new_n845), .A2(new_n1167), .B1(new_n786), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(G128), .ZN(new_n1171));
  OAI22_X1  g0971(.A1(new_n795), .A2(new_n852), .B1(new_n798), .B2(new_n1171), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT114), .Z(new_n1173));
  OAI22_X1  g0973(.A1(new_n798), .A2(new_n791), .B1(new_n785), .B2(new_n222), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G116), .B2(new_n982), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G87), .A2(new_n988), .B1(new_n845), .B2(G107), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1175), .A2(new_n806), .A3(new_n1118), .A4(new_n1176), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n793), .A2(new_n202), .B1(new_n788), .B2(new_n503), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT115), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1170), .A2(new_n1173), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1162), .B1(new_n1180), .B2(new_n782), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n931), .B1(new_n918), .B2(new_n919), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n925), .A2(new_n926), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n928), .A2(new_n910), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n896), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT39), .B1(new_n1186), .B2(new_n917), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1181), .B1(new_n1188), .B2(new_n824), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1161), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1160), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT116), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1160), .A2(new_n1190), .A3(KEYINPUT116), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(G378));
  NAND2_X1  g0996(.A1(new_n902), .A2(new_n272), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n312), .B(new_n1197), .Z(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1198), .B(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n823), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n779), .B1(new_n843), .B2(G50), .ZN(new_n1203));
  INV_X1    g1003(.A(G125), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n795), .A2(new_n1171), .B1(new_n798), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G132), .A2(new_n845), .B1(new_n988), .B2(new_n1168), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1206), .B1(new_n267), .B2(new_n808), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1205), .B(new_n1207), .C1(G137), .C2(new_n786), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OR2_X1    g1009(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(KEYINPUT59), .ZN(new_n1211));
  AOI211_X1 g1011(.A(G33), .B(G41), .C1(new_n854), .C2(G159), .ZN(new_n1212));
  INV_X1    g1012(.A(G124), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1212), .B1(new_n1213), .B2(new_n788), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT117), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1210), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(G77), .A2(new_n988), .B1(new_n789), .B2(G283), .ZN(new_n1217));
  OAI221_X1 g1017(.A(new_n1217), .B1(new_n201), .B2(new_n793), .C1(new_n477), .C2(new_n795), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G116), .A2(new_n799), .B1(new_n845), .B2(G97), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n325), .B2(new_n785), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n399), .A2(new_n291), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n986), .A4(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1221), .B(new_n253), .C1(G33), .C2(G41), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1222), .A2(KEYINPUT58), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1216), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1203), .B1(new_n1226), .B2(new_n782), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1202), .A2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(G330), .B1(new_n964), .B2(new_n966), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT118), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1201), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n935), .B1(new_n1188), .B2(new_n924), .ZN(new_n1233));
  OAI211_X1 g1033(.A(KEYINPUT118), .B(G330), .C1(new_n964), .C2(new_n966), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1147), .A2(new_n919), .A3(new_n918), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1235), .B2(new_n1233), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1232), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n960), .A2(new_n963), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n930), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT40), .B1(new_n1240), .B2(new_n963), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n713), .B1(new_n1239), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(KEYINPUT118), .C1(new_n937), .C2(new_n953), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1231), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1238), .A2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1228), .B1(new_n1246), .B2(new_n777), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1132), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1159), .A2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1250), .A2(KEYINPUT57), .A3(new_n1245), .A4(new_n1238), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n732), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1243), .A2(new_n1231), .A3(new_n1244), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1231), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT57), .B1(new_n1255), .B2(new_n1250), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1248), .B1(new_n1252), .B2(new_n1256), .ZN(G375));
  INV_X1    g1057(.A(new_n1143), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n950), .A2(new_n823), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n834), .B1(new_n843), .B2(G68), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n862), .A2(new_n803), .B1(new_n788), .B2(new_n801), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n979), .B(new_n1261), .C1(G283), .C2(new_n982), .ZN(new_n1262));
  OAI22_X1  g1062(.A1(new_n222), .A2(new_n802), .B1(new_n785), .B2(new_n477), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1263), .B1(G294), .B2(new_n799), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n806), .A3(new_n1080), .A4(new_n1264), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n845), .A2(new_n1168), .B1(new_n854), .B2(G58), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n568), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G50), .B2(new_n814), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n982), .A2(new_n1167), .B1(new_n799), .B2(G132), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n267), .C2(new_n785), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n802), .A2(new_n812), .B1(new_n788), .B2(new_n1171), .ZN(new_n1271));
  XOR2_X1   g1071(.A(new_n1271), .B(KEYINPUT119), .Z(new_n1272));
  OAI21_X1  g1072(.A(new_n1265), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1260), .B1(new_n1273), .B2(new_n782), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1258), .A2(new_n778), .B1(new_n1259), .B2(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1249), .A2(new_n1258), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1145), .A2(new_n1045), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(G381));
  OR2_X1    g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NOR4_X1   g1079(.A1(G381), .A2(G390), .A3(new_n1279), .A4(G384), .ZN(new_n1280));
  INV_X1    g1080(.A(G387), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(KEYINPUT120), .ZN(new_n1283));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1191), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  OR2_X1    g1086(.A1(new_n1283), .A2(new_n1286), .ZN(G407));
  INV_X1    g1087(.A(new_n707), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(new_n1288), .C2(new_n1286), .ZN(G409));
  XNOR2_X1  g1089(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1159), .A2(new_n1249), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1291), .A2(new_n1246), .A3(new_n1043), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1285), .B1(new_n1292), .B2(new_n1247), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1293), .B1(G375), .B2(new_n1195), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n707), .A2(G213), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1295), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1132), .A2(new_n1143), .A3(KEYINPUT60), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1298), .A2(new_n732), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT60), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1144), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1301), .B2(new_n1276), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(G384), .A3(new_n1275), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(G384), .B1(new_n1302), .B2(new_n1275), .ZN(new_n1305));
  OAI211_X1 g1105(.A(G2897), .B(new_n1297), .C1(new_n1304), .C2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1305), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1297), .A2(G2897), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1303), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1290), .B1(new_n1296), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT57), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n1291), .B2(new_n1246), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1314), .A2(new_n732), .A3(new_n1251), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(new_n1193), .A3(new_n1194), .A4(new_n1248), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1297), .B1(new_n1316), .B2(new_n1293), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT62), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1319));
  AND4_X1   g1119(.A1(KEYINPUT62), .A2(new_n1294), .A3(new_n1295), .A4(new_n1318), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1312), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  OAI211_X1 g1121(.A(G390), .B(new_n1009), .C1(new_n1049), .C2(new_n1061), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1322), .A2(KEYINPUT123), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(G393), .B(G396), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(G390), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G387), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1322), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1325), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT123), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1327), .A2(new_n1324), .A3(new_n1330), .A4(new_n1322), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  XNOR2_X1  g1132(.A(new_n1332), .B(KEYINPUT126), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1321), .A2(new_n1333), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1318), .A2(KEYINPUT63), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1294), .A2(new_n1335), .A3(new_n1295), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(KEYINPUT124), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT124), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1317), .A2(new_n1338), .A3(new_n1335), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1307), .A2(new_n1303), .ZN(new_n1341));
  AOI211_X1 g1141(.A(new_n1297), .B(new_n1341), .C1(new_n1316), .C2(new_n1293), .ZN(new_n1342));
  XNOR2_X1  g1142(.A(KEYINPUT121), .B(KEYINPUT63), .ZN(new_n1343));
  OAI21_X1  g1143(.A(KEYINPUT122), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1331), .ZN(new_n1346));
  AOI22_X1  g1146(.A1(new_n1323), .A2(new_n1324), .B1(new_n1327), .B2(new_n1322), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1345), .B1(new_n1346), .B2(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1310), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT122), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1343), .ZN(new_n1352));
  OAI211_X1 g1152(.A(new_n1351), .B(new_n1352), .C1(new_n1296), .C2(new_n1341), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1340), .A2(new_n1344), .A3(new_n1350), .A4(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1334), .A2(new_n1354), .ZN(G405));
  OR2_X1    g1155(.A1(new_n1332), .A2(KEYINPUT127), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1316), .B(new_n1318), .C1(new_n1284), .C2(new_n1191), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1284), .A2(new_n1191), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1316), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1341), .B1(new_n1358), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1332), .A2(KEYINPUT127), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1356), .A2(new_n1357), .A3(new_n1360), .A4(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1360), .A2(new_n1357), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1363), .A2(KEYINPUT127), .A3(new_n1332), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1362), .A2(new_n1364), .ZN(G402));
endmodule


