//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G228gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G155gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT80), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT80), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(G155gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n209), .A3(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT2), .ZN(new_n211));
  XNOR2_X1  g010(.A(G141gat), .B(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n206), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT79), .ZN(new_n219));
  AND3_X1   g018(.A1(new_n215), .A2(new_n219), .A3(new_n216), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n219), .B1(new_n215), .B2(new_n216), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n216), .A2(KEYINPUT2), .ZN(new_n222));
  OAI22_X1  g021(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n212), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT81), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n218), .A2(new_n223), .A3(KEYINPUT81), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT77), .B(KEYINPUT29), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G197gat), .B(G204gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232));
  INV_X1    g031(.A(G211gat), .ZN(new_n233));
  INV_X1    g032(.A(G218gat), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G211gat), .B(G218gat), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n230), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n236), .A2(new_n238), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n228), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n218), .A2(new_n223), .A3(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n246), .A2(new_n229), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n238), .A2(KEYINPUT75), .ZN(new_n248));
  OR2_X1    g047(.A1(new_n248), .A2(new_n236), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n236), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n205), .B1(new_n244), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n251), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(KEYINPUT76), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT76), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n251), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n247), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT3), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n224), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n205), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n254), .A2(new_n264), .A3(KEYINPUT87), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT87), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n259), .A2(new_n263), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n204), .B1(new_n243), .B2(new_n252), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G78gat), .B(G106gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(G22gat), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n265), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT87), .B1(new_n254), .B2(new_n264), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n266), .A3(new_n268), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n203), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n271), .B1(new_n265), .B2(new_n269), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n274), .A2(new_n275), .A3(new_n273), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(new_n202), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT32), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT26), .ZN(new_n285));
  AND2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n286), .A2(KEYINPUT26), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n283), .B(new_n285), .C1(new_n287), .C2(new_n284), .ZN(new_n288));
  INV_X1    g087(.A(G190gat), .ZN(new_n289));
  AND2_X1   g088(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n294));
  INV_X1    g093(.A(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT67), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(KEYINPUT28), .B(new_n289), .C1(new_n293), .C2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n297), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT28), .B1(new_n300), .B2(new_n289), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n288), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n292), .B1(new_n290), .B2(new_n291), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n296), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n307));
  AOI21_X1  g106(.A(G190gat), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n301), .B1(new_n308), .B2(KEYINPUT28), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT68), .B1(new_n309), .B2(new_n288), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G113gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(G120gat), .ZN(new_n313));
  INV_X1    g112(.A(G120gat), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n314), .A2(G113gat), .ZN(new_n315));
  OAI21_X1  g114(.A(KEYINPUT70), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G134gat), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G127gat), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XOR2_X1   g120(.A(KEYINPUT71), .B(KEYINPUT1), .Z(new_n322));
  NAND2_X1  g121(.A1(new_n314), .A2(G113gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n312), .A2(G120gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n316), .A2(new_n321), .A3(new_n322), .A4(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT69), .ZN(new_n328));
  OR3_X1    g127(.A1(new_n319), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(G113gat), .B(G120gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n329), .C1(KEYINPUT1), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT25), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT66), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n295), .A2(new_n289), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT24), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n337), .B1(new_n338), .B2(new_n283), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n334), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n286), .B1(KEYINPUT23), .B2(new_n284), .ZN(new_n342));
  INV_X1    g141(.A(G169gat), .ZN(new_n343));
  INV_X1    g142(.A(G176gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT64), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT64), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT23), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT65), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n342), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n354), .B1(new_n342), .B2(new_n350), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n339), .A2(new_n335), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n353), .B1(new_n358), .B2(KEYINPUT25), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n311), .A2(new_n333), .A3(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n311), .A2(new_n359), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n332), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n311), .A2(KEYINPUT72), .A3(new_n333), .A4(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n282), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n368), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT33), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g172(.A(G71gat), .B(G99gat), .Z(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT73), .ZN(new_n375));
  XOR2_X1   g174(.A(G15gat), .B(G43gat), .Z(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  NAND3_X1  g176(.A1(new_n370), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  AOI221_X4 g177(.A(new_n282), .B1(KEYINPUT33), .B2(new_n377), .C1(new_n366), .C2(new_n368), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n362), .A2(new_n364), .A3(new_n367), .A4(new_n365), .ZN(new_n381));
  NAND2_X1  g180(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(KEYINPUT74), .A2(KEYINPUT34), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n381), .B2(new_n383), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n388), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT33), .B1(new_n366), .B2(new_n368), .ZN(new_n391));
  INV_X1    g190(.A(new_n377), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n369), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n390), .B1(new_n393), .B2(new_n379), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n281), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT35), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n218), .A2(new_n223), .A3(KEYINPUT81), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT81), .B1(new_n218), .B2(new_n223), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n397), .B(new_n333), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT85), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT85), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n228), .A2(new_n402), .A3(new_n397), .A4(new_n333), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n218), .A2(new_n223), .A3(new_n327), .A4(new_n331), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n224), .A2(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n332), .A3(new_n246), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n406), .A2(new_n407), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n224), .A2(new_n332), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT82), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(new_n404), .ZN(new_n415));
  INV_X1    g214(.A(new_n408), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n224), .A2(new_n332), .A3(KEYINPUT82), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT4), .B(new_n333), .C1(new_n398), .C2(new_n399), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n397), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n408), .A3(new_n410), .A4(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n412), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  AND4_X1   g222(.A1(new_n412), .A2(new_n422), .A3(KEYINPUT5), .A4(new_n418), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n411), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(G1gat), .B(G29gat), .Z(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT84), .B(KEYINPUT0), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G57gat), .B(G85gat), .ZN(new_n429));
  XOR2_X1   g228(.A(new_n428), .B(new_n429), .Z(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  INV_X1    g231(.A(new_n430), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n411), .B(new_n433), .C1(new_n423), .C2(new_n424), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n432), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n412), .A3(new_n422), .ZN(new_n437));
  INV_X1    g236(.A(new_n422), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n439));
  OAI21_X1  g238(.A(KEYINPUT83), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n433), .B1(new_n441), .B2(new_n411), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n436), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n435), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n303), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT29), .B1(new_n359), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G226gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT78), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n363), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n351), .A2(KEYINPUT65), .ZN(new_n451));
  INV_X1    g250(.A(new_n357), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n342), .A2(new_n350), .A3(new_n354), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n454), .A2(new_n334), .B1(new_n352), .B2(new_n341), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n260), .B1(new_n455), .B2(new_n303), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT78), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n447), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(new_n251), .A3(new_n450), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n363), .A2(new_n447), .A3(new_n229), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n256), .A2(new_n258), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n359), .A2(new_n448), .A3(new_n445), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g263(.A(G8gat), .B(G36gat), .Z(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(G64gat), .ZN(new_n466));
  INV_X1    g265(.A(G92gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n459), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(KEYINPUT30), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT30), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n459), .A2(new_n473), .A3(new_n463), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n395), .A2(new_n396), .A3(new_n444), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n394), .A2(new_n389), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n272), .A2(new_n276), .A3(new_n203), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n202), .B1(new_n278), .B2(new_n279), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n436), .A2(new_n442), .ZN(new_n482));
  AOI211_X1 g281(.A(new_n432), .B(new_n433), .C1(new_n441), .C2(new_n411), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n475), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n444), .A2(KEYINPUT86), .A3(new_n475), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n476), .B1(new_n488), .B2(new_n396), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n281), .A3(new_n487), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n394), .A2(new_n389), .A3(KEYINPUT36), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT36), .B1(new_n394), .B2(new_n389), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g292(.A1(new_n449), .A2(new_n450), .A3(new_n458), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n460), .A2(new_n462), .ZN(new_n495));
  OAI22_X1  g294(.A1(new_n494), .A2(new_n251), .B1(new_n495), .B2(new_n461), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n470), .B1(new_n496), .B2(KEYINPUT37), .ZN(new_n497));
  XOR2_X1   g296(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n498));
  NAND3_X1  g297(.A1(new_n459), .A2(new_n463), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT89), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n459), .A2(new_n463), .A3(new_n501), .A4(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT38), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n497), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n505), .A2(new_n443), .A3(new_n435), .A4(new_n471), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT90), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n470), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n507), .B1(new_n509), .B2(KEYINPUT38), .ZN(new_n510));
  AOI211_X1 g309(.A(KEYINPUT90), .B(new_n504), .C1(new_n503), .C2(new_n508), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n408), .B1(new_n406), .B2(new_n410), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT39), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n430), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(KEYINPUT40), .A3(new_n517), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n518), .A2(new_n472), .A3(new_n431), .A4(new_n474), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT40), .B1(new_n516), .B2(new_n517), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n480), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n490), .B(new_n493), .C1(new_n512), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n489), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT16), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(G1gat), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n526), .B1(G1gat), .B2(new_n524), .ZN(new_n527));
  XOR2_X1   g326(.A(new_n527), .B(G8gat), .Z(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n529), .A2(KEYINPUT91), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(KEYINPUT91), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT15), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G29gat), .A2(G36gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(KEYINPUT92), .ZN(new_n534));
  OR3_X1    g333(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n532), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g338(.A1(new_n535), .A2(KEYINPUT93), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n535), .A2(KEYINPUT93), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n532), .A2(new_n542), .A3(new_n543), .A4(new_n534), .ZN(new_n544));
  OR2_X1    g343(.A1(new_n544), .A2(KEYINPUT94), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(KEYINPUT94), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n528), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552));
  INV_X1    g351(.A(new_n547), .ZN(new_n553));
  INV_X1    g352(.A(new_n528), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n551), .A2(new_n552), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n553), .B2(new_n554), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n547), .A2(KEYINPUT95), .A3(new_n528), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n555), .A3(new_n561), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n552), .B(KEYINPUT13), .Z(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n551), .A2(KEYINPUT18), .A3(new_n552), .A4(new_n555), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n558), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT11), .B(G169gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G197gat), .ZN(new_n568));
  XOR2_X1   g367(.A(G113gat), .B(G141gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT12), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n558), .A2(new_n571), .A3(new_n564), .A4(new_n565), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n523), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT96), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT96), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n523), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT21), .ZN(new_n581));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G71gat), .B(G78gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n584), .B(new_n585), .Z(new_n586));
  OAI21_X1  g385(.A(new_n528), .B1(new_n581), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n587), .B(G183gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(G231gat), .A2(G233gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(G127gat), .B(G155gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n591), .B(new_n233), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n586), .A2(new_n581), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n604));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT97), .B(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n608), .A2(new_n609), .B1(KEYINPUT8), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT7), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614));
  XNOR2_X1  g413(.A(G99gat), .B(G106gat), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n611), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n615), .A2(new_n614), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT99), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n549), .B2(new_n550), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n623));
  INV_X1    g422(.A(new_n620), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n623), .B1(new_n547), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n627), .A2(new_n628), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n607), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n630), .A2(new_n607), .A3(new_n631), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n584), .B(new_n585), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n616), .A2(new_n617), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n616), .A2(new_n617), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n618), .A2(new_n586), .A3(new_n619), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  NAND2_X1  g441(.A1(G230gat), .A2(G233gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n641), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n642), .B1(new_n641), .B2(new_n644), .ZN(new_n647));
  OAI21_X1  g446(.A(KEYINPUT100), .B1(new_n641), .B2(KEYINPUT10), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n620), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n639), .A2(new_n640), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n643), .B(KEYINPUT104), .Z(new_n654));
  AOI211_X1 g453(.A(new_n646), .B(new_n647), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT103), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n314), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n647), .ZN(new_n661));
  OAI21_X1  g460(.A(KEYINPUT102), .B1(new_n646), .B2(new_n647), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n643), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n659), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n602), .A2(new_n635), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n602), .A2(new_n635), .A3(KEYINPUT105), .A4(new_n666), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n580), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n444), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  INV_X1    g474(.A(new_n475), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n580), .A2(new_n676), .A3(new_n671), .ZN(new_n677));
  XNOR2_X1  g476(.A(KEYINPUT16), .B(G8gat), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n677), .B2(G8gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(KEYINPUT106), .B2(new_n680), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n678), .A2(KEYINPUT106), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n679), .A2(new_n681), .B1(new_n683), .B2(new_n684), .ZN(G1325gat));
  AOI21_X1  g484(.A(G15gat), .B1(new_n672), .B2(new_n477), .ZN(new_n686));
  INV_X1    g485(.A(new_n493), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(G15gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT107), .Z(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n672), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n672), .A2(new_n281), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  OR2_X1    g492(.A1(new_n633), .A2(new_n634), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n490), .A2(new_n493), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n510), .A2(new_n511), .ZN(new_n696));
  INV_X1    g495(.A(new_n506), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n521), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n477), .A2(new_n396), .A3(new_n480), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n484), .ZN(new_n701));
  NOR2_X1   g500(.A1(new_n484), .A2(new_n485), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT86), .B1(new_n444), .B2(new_n475), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n395), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n701), .B1(new_n704), .B2(KEYINPUT35), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n694), .B1(new_n699), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n602), .A2(new_n665), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n523), .A2(KEYINPUT44), .A3(new_n694), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n708), .A2(new_n575), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n711), .A2(KEYINPUT108), .A3(new_n444), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT108), .B1(new_n711), .B2(new_n444), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(G29gat), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n578), .B1(new_n523), .B2(new_n575), .ZN(new_n715));
  INV_X1    g514(.A(new_n575), .ZN(new_n716));
  AOI211_X1 g515(.A(KEYINPUT96), .B(new_n716), .C1(new_n489), .C2(new_n522), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n694), .B(new_n709), .C1(new_n715), .C2(new_n717), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(G29gat), .A3(new_n444), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR4_X1   g520(.A1(new_n718), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n444), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n714), .B1(new_n721), .B2(new_n722), .ZN(G1328gat));
  NOR3_X1   g522(.A1(new_n718), .A2(G36gat), .A3(new_n475), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(G36gat), .B1(new_n711), .B2(new_n475), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n724), .A2(new_n725), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(G1329gat));
  INV_X1    g528(.A(new_n709), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n577), .B2(new_n579), .ZN(new_n731));
  INV_X1    g530(.A(G43gat), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n731), .A2(new_n732), .A3(new_n477), .A4(new_n694), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT47), .ZN(new_n734));
  OAI21_X1  g533(.A(G43gat), .B1(new_n711), .B2(new_n493), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n734), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  INV_X1    g537(.A(G50gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n731), .A2(new_n739), .A3(new_n281), .A4(new_n694), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  OAI21_X1  g540(.A(G50gat), .B1(new_n711), .B2(new_n480), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(G1331gat));
  NAND2_X1  g544(.A1(new_n602), .A2(new_n635), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n489), .B2(new_n522), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n575), .A2(new_n666), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n673), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n475), .ZN(new_n753));
  NOR2_X1   g552(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n754));
  AND2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n753), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n753), .B2(new_n754), .ZN(G1333gat));
  OAI21_X1  g556(.A(G71gat), .B1(new_n749), .B2(new_n493), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n750), .A2(new_n477), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n758), .B1(new_n759), .B2(G71gat), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g560(.A1(new_n750), .A2(new_n281), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g562(.A(new_n635), .B1(new_n489), .B2(new_n522), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n602), .A2(new_n575), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n765), .B1(new_n764), .B2(new_n766), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(new_n666), .ZN(new_n769));
  AOI21_X1  g568(.A(G85gat), .B1(new_n769), .B2(new_n673), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT44), .B1(new_n523), .B2(new_n694), .ZN(new_n771));
  AOI211_X1 g570(.A(new_n707), .B(new_n635), .C1(new_n489), .C2(new_n522), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n665), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n444), .A2(new_n609), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n770), .B1(new_n774), .B2(new_n775), .ZN(G1336gat));
  NOR2_X1   g575(.A1(new_n771), .A2(new_n772), .ZN(new_n777));
  INV_X1    g576(.A(new_n773), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n777), .A2(KEYINPUT110), .A3(new_n676), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n708), .A2(new_n676), .A3(new_n710), .A4(new_n778), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n608), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n523), .A2(new_n694), .A3(new_n766), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT51), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n475), .A2(G92gat), .ZN(new_n789));
  AND4_X1   g588(.A1(new_n665), .A2(new_n787), .A3(new_n788), .A4(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n784), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n780), .A2(new_n793), .A3(new_n783), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n780), .B2(new_n783), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n790), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n792), .B1(new_n796), .B2(new_n785), .ZN(G1337gat));
  INV_X1    g596(.A(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n769), .A2(new_n798), .A3(new_n477), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n774), .A2(new_n687), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n800), .B2(new_n798), .ZN(G1338gat));
  NOR2_X1   g600(.A1(new_n767), .A2(new_n768), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT111), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n480), .A2(G106gat), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n665), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n787), .A2(new_n665), .A3(new_n788), .A4(new_n804), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n708), .A2(new_n281), .A3(new_n710), .A4(new_n778), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(G106gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G106gat), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n808), .A2(KEYINPUT112), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n812), .B(new_n806), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(G1339gat));
  INV_X1    g616(.A(new_n602), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  INV_X1    g618(.A(new_n654), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n648), .A2(new_n820), .A3(new_n649), .A4(new_n652), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n653), .A2(new_n824), .A3(new_n654), .ZN(new_n825));
  INV_X1    g624(.A(new_n659), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n819), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n822), .A2(KEYINPUT55), .A3(new_n826), .A4(new_n825), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n829), .A2(new_n830), .A3(new_n664), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n664), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n575), .A2(new_n828), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n562), .A2(new_n563), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n552), .B1(new_n551), .B2(new_n555), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n570), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n574), .A2(new_n665), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n694), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n828), .A3(new_n831), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n574), .A2(new_n837), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n840), .A2(new_n635), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n818), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n667), .A2(new_n575), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n481), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n676), .A2(new_n444), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n575), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n665), .ZN(new_n851));
  XOR2_X1   g650(.A(KEYINPUT114), .B(G120gat), .Z(new_n852));
  XNOR2_X1  g651(.A(new_n851), .B(new_n852), .ZN(G1341gat));
  NAND2_X1  g652(.A1(new_n848), .A2(new_n602), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n319), .A3(new_n694), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n848), .A2(new_n694), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n857), .B(new_n858), .C1(new_n319), .C2(new_n859), .ZN(G1343gat));
  NOR2_X1   g659(.A1(new_n687), .A2(new_n444), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n834), .A2(new_n838), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n635), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n840), .A2(new_n635), .A3(new_n841), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n602), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n861), .B(new_n281), .C1(new_n865), .C2(new_n844), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n480), .B1(new_n843), .B2(new_n845), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n861), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n716), .A2(G141gat), .ZN(new_n871));
  XOR2_X1   g670(.A(new_n871), .B(KEYINPUT117), .Z(new_n872));
  NAND4_X1  g671(.A1(new_n868), .A2(new_n475), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT119), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n493), .A2(new_n847), .ZN(new_n875));
  XOR2_X1   g674(.A(KEYINPUT115), .B(KEYINPUT57), .Z(new_n876));
  NOR2_X1   g675(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT116), .B1(new_n823), .B2(new_n827), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT116), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n822), .A2(new_n880), .A3(new_n826), .A4(new_n825), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n879), .A2(new_n819), .A3(new_n881), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n575), .A2(new_n664), .A3(new_n829), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n694), .B1(new_n883), .B2(new_n838), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n818), .B1(new_n884), .B2(new_n842), .ZN(new_n885));
  AOI211_X1 g684(.A(new_n878), .B(new_n480), .C1(new_n885), .C2(new_n845), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n575), .B(new_n875), .C1(new_n877), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(G141gat), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n874), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT58), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n890), .B1(new_n873), .B2(KEYINPUT119), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n866), .A2(new_n676), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n887), .A2(G141gat), .B1(new_n872), .B2(new_n892), .ZN(new_n893));
  OAI22_X1  g692(.A1(new_n889), .A2(new_n891), .B1(new_n890), .B2(new_n893), .ZN(G1344gat));
  OAI211_X1 g693(.A(new_n665), .B(new_n875), .C1(new_n877), .C2(new_n886), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(G148gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n843), .A2(new_n845), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n898), .A2(new_n281), .A3(new_n876), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n669), .A2(new_n716), .A3(new_n670), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n901), .B2(new_n281), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n665), .B(new_n875), .C1(new_n899), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n896), .B1(new_n903), .B2(G148gat), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n666), .A2(G148gat), .ZN(new_n905));
  NAND4_X1  g704(.A1(new_n868), .A2(new_n475), .A3(new_n870), .A4(new_n905), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(KEYINPUT120), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n897), .A2(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G1345gat));
  AND2_X1   g708(.A1(new_n207), .A2(new_n209), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n875), .B1(new_n877), .B2(new_n886), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n818), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n868), .A2(new_n475), .A3(new_n870), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n818), .A2(new_n910), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(G1346gat));
  OAI21_X1  g714(.A(G162gat), .B1(new_n911), .B2(new_n635), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n694), .A2(new_n214), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n913), .B2(new_n917), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n673), .A2(new_n475), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  AOI211_X1 g719(.A(new_n481), .B(new_n920), .C1(new_n843), .C2(new_n845), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n575), .C1(KEYINPUT121), .C2(new_n343), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n343), .A2(KEYINPUT121), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(G1348gat));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n665), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g725(.A1(new_n306), .A2(new_n307), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n846), .A2(new_n927), .A3(new_n602), .A4(new_n919), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n921), .A2(new_n930), .A3(new_n927), .A4(new_n602), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n921), .A2(new_n602), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT123), .B1(new_n933), .B2(G183gat), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n934), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n289), .A3(new_n694), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT124), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n921), .A2(new_n694), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(G190gat), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n945), .A2(KEYINPUT61), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT61), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n943), .A2(new_n944), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n941), .A2(new_n947), .A3(new_n949), .ZN(G1351gat));
  OR2_X1    g749(.A1(new_n899), .A2(new_n902), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n687), .A2(new_n920), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n716), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n869), .A2(new_n952), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n955), .B(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n958), .A3(new_n575), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n954), .A2(new_n959), .ZN(G1352gat));
  XNOR2_X1  g759(.A(KEYINPUT127), .B(G204gat), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n955), .A2(new_n665), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  OR2_X1    g763(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n951), .A2(new_n665), .A3(new_n952), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n964), .B(new_n965), .C1(new_n966), .C2(new_n962), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n957), .A2(new_n233), .A3(new_n602), .ZN(new_n968));
  OAI211_X1 g767(.A(new_n602), .B(new_n952), .C1(new_n899), .C2(new_n902), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  INV_X1    g771(.A(new_n953), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n635), .A2(new_n234), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n955), .A2(KEYINPUT126), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n955), .A2(KEYINPUT126), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(new_n694), .A3(new_n976), .ZN(new_n977));
  AOI22_X1  g776(.A1(new_n973), .A2(new_n974), .B1(new_n977), .B2(new_n234), .ZN(G1355gat));
endmodule


