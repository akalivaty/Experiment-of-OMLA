//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948;
  XOR2_X1   g000(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G227gat), .A2(G233gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n209), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n208), .A2(KEYINPUT25), .A3(new_n210), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT24), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G183gat), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n212), .B1(new_n222), .B2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n217), .A2(new_n224), .A3(new_n220), .A4(new_n221), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n220), .A2(new_n221), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT25), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n223), .A2(new_n225), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n206), .A2(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n213), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n211), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n235), .A2(new_n206), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n218), .A2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G183gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n219), .B1(new_n242), .B2(KEYINPUT28), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT68), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(KEYINPUT28), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  AOI21_X1  g047(.A(G190gat), .B1(new_n248), .B2(KEYINPUT67), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n246), .A2(new_n247), .A3(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n245), .B1(new_n244), .B2(new_n250), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n237), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n245), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n241), .A2(KEYINPUT68), .A3(new_n243), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n247), .B1(new_n246), .B2(new_n249), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n244), .A2(new_n245), .A3(new_n250), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n261), .A2(KEYINPUT69), .A3(new_n237), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n231), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  XOR2_X1   g062(.A(G113gat), .B(G120gat), .Z(new_n264));
  INV_X1    g063(.A(KEYINPUT1), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G127gat), .B(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n264), .A2(new_n265), .A3(new_n267), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n263), .A2(new_n272), .ZN(new_n273));
  AOI211_X1 g072(.A(new_n271), .B(new_n231), .C1(new_n255), .C2(new_n262), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n205), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT32), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(G15gat), .B(G43gat), .Z(new_n279));
  XNOR2_X1  g078(.A(G71gat), .B(G99gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n276), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n275), .B(KEYINPUT32), .C1(new_n277), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n223), .A2(new_n225), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n229), .A2(new_n230), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(new_n261), .B2(new_n237), .ZN(new_n288));
  INV_X1    g087(.A(new_n237), .ZN(new_n289));
  AOI211_X1 g088(.A(new_n254), .B(new_n289), .C1(new_n259), .C2(new_n260), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(new_n271), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n263), .A2(new_n272), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n292), .A2(new_n293), .A3(new_n204), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n282), .A2(new_n284), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n282), .B2(new_n284), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n203), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n294), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n204), .B1(new_n292), .B2(new_n293), .ZN(new_n299));
  INV_X1    g098(.A(new_n277), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n281), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n284), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n298), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n282), .A2(new_n284), .A3(new_n294), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n202), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n297), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT74), .B(G197gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(G211gat), .ZN(new_n312));
  INV_X1    g111(.A(G218gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n311), .B1(KEYINPUT22), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(G211gat), .B(G218gat), .Z(new_n316));
  XNOR2_X1  g115(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G155gat), .ZN(new_n319));
  INV_X1    g118(.A(G162gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n324), .B2(KEYINPUT2), .ZN(new_n325));
  XNOR2_X1  g124(.A(KEYINPUT78), .B(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(G141gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G148gat), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n329), .A2(G141gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n325), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  XNOR2_X1  g131(.A(G141gat), .B(G148gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n322), .B(new_n324), .C1(new_n333), .C2(KEYINPUT2), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n318), .B1(KEYINPUT29), .B2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT3), .B1(new_n317), .B2(new_n338), .ZN(new_n339));
  XOR2_X1   g138(.A(KEYINPUT78), .B(G148gat), .Z(new_n340));
  AOI21_X1  g139(.A(new_n330), .B1(new_n340), .B2(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n321), .B1(new_n342), .B2(new_n323), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n334), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n337), .B1(new_n339), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT83), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n350), .B(G50gat), .ZN(new_n351));
  NAND2_X1  g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n352), .B(G22gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n351), .B(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n348), .B(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n309), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT29), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n263), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n287), .A2(new_n253), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n362), .A2(new_n357), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n361), .A2(new_n317), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n358), .B1(new_n362), .B2(new_n338), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n366), .B1(new_n263), .B2(new_n357), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n291), .A2(KEYINPUT75), .A3(new_n358), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n364), .B1(new_n369), .B2(new_n317), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI211_X1 g171(.A(new_n318), .B(new_n365), .C1(new_n367), .C2(new_n368), .ZN(new_n373));
  OAI21_X1  g172(.A(KEYINPUT76), .B1(new_n373), .B2(new_n364), .ZN(new_n374));
  XNOR2_X1  g173(.A(G8gat), .B(G36gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(G64gat), .B(G92gat), .ZN(new_n376));
  XOR2_X1   g175(.A(new_n375), .B(new_n376), .Z(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n372), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n372), .A2(new_n374), .A3(new_n381), .A4(new_n378), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n271), .A2(new_n344), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n331), .A2(new_n334), .B1(new_n269), .B2(new_n270), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(KEYINPUT4), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n335), .A3(new_n271), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n271), .B2(new_n344), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n390), .A2(new_n392), .A3(new_n388), .A4(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n388), .ZN(new_n396));
  OAI211_X1 g195(.A(KEYINPUT80), .B(new_n396), .C1(new_n385), .C2(new_n386), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n389), .A2(new_n395), .A3(KEYINPUT5), .A4(new_n397), .ZN(new_n398));
  XOR2_X1   g197(.A(G1gat), .B(G29gat), .Z(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G57gat), .B(G85gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n392), .A2(new_n388), .ZN(new_n404));
  INV_X1    g203(.A(new_n393), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n385), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT5), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n385), .A2(KEYINPUT4), .ZN(new_n408));
  NAND4_X1  g207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n398), .A2(new_n403), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n403), .B1(new_n398), .B2(new_n409), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n411), .A2(new_n412), .A3(KEYINPUT6), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(KEYINPUT6), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n370), .A2(new_n377), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n418), .B(KEYINPUT30), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n383), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT35), .B1(new_n356), .B2(new_n420), .ZN(new_n421));
  AND2_X1   g220(.A1(new_n383), .A2(new_n419), .ZN(new_n422));
  INV_X1    g221(.A(new_n355), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n297), .B2(new_n308), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT84), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n413), .B2(new_n415), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n414), .A2(KEYINPUT84), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT35), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n422), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n295), .A2(new_n296), .A3(new_n203), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n202), .B1(new_n306), .B2(new_n307), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT36), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT72), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n309), .A2(new_n435), .A3(KEYINPUT36), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT36), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n297), .A2(new_n437), .A3(new_n308), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT73), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n297), .A2(new_n440), .A3(new_n308), .A4(new_n437), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n434), .A2(new_n436), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n420), .A2(new_n423), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n408), .A2(new_n392), .A3(new_n406), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n396), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n387), .A2(new_n388), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n445), .A2(KEYINPUT39), .A3(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(new_n403), .C1(KEYINPUT39), .C2(new_n445), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT40), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n412), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n449), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n383), .B2(new_n419), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n377), .B1(new_n370), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n369), .A2(new_n318), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n361), .A2(new_n363), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n458), .B2(new_n317), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT38), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n461), .A2(new_n426), .A3(new_n418), .A4(new_n427), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT38), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n372), .A2(new_n374), .A3(KEYINPUT37), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(new_n464), .B2(new_n456), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n355), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n443), .B1(new_n454), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n430), .B1(new_n442), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT85), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n430), .B(new_n470), .C1(new_n442), .C2(new_n467), .ZN(new_n471));
  XNOR2_X1  g270(.A(G113gat), .B(G141gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G197gat), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT11), .B(G169gat), .Z(new_n474));
  XNOR2_X1  g273(.A(new_n473), .B(new_n474), .ZN(new_n475));
  XOR2_X1   g274(.A(new_n475), .B(KEYINPUT12), .Z(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G29gat), .ZN(new_n478));
  INV_X1    g277(.A(G36gat), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT14), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n481), .A2(G29gat), .A3(G36gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT86), .B(G36gat), .ZN(new_n483));
  AOI211_X1 g282(.A(new_n480), .B(new_n482), .C1(G29gat), .C2(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n486));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n486), .B2(new_n487), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT17), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT16), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n491), .B1(new_n492), .B2(G1gat), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(G1gat), .B2(new_n491), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n496), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n489), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n497), .A2(KEYINPUT18), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n489), .B(new_n498), .ZN(new_n502));
  XOR2_X1   g301(.A(new_n500), .B(KEYINPUT13), .Z(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n477), .B1(new_n505), .B2(KEYINPUT87), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n501), .A2(new_n504), .ZN(new_n507));
  INV_X1    g306(.A(new_n499), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n508), .B1(new_n490), .B2(new_n496), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT18), .B1(new_n509), .B2(new_n500), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n506), .B(new_n511), .Z(new_n512));
  INV_X1    g311(.A(G230gat), .ZN(new_n513));
  INV_X1    g312(.A(G233gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n518));
  OR2_X1    g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G71gat), .B(G78gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT93), .ZN(new_n525));
  NAND2_X1  g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT93), .B1(new_n528), .B2(new_n523), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT7), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT91), .ZN(new_n534));
  AND2_X1   g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G85gat), .ZN(new_n537));
  INV_X1    g336(.A(G92gat), .ZN(new_n538));
  OAI211_X1 g337(.A(KEYINPUT91), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT92), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(KEYINPUT8), .A2(new_n526), .B1(new_n537), .B2(new_n538), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n530), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n536), .A2(KEYINPUT92), .A3(new_n539), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT92), .B1(new_n536), .B2(new_n539), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n530), .B(new_n545), .C1(new_n547), .C2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n522), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT96), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n553));
  INV_X1    g352(.A(new_n530), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n555), .A2(new_n521), .A3(new_n549), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n552), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n555), .A2(new_n549), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n522), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT10), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT10), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n516), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n557), .A2(new_n515), .A3(new_n559), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(G120gat), .B(G148gat), .Z(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT97), .ZN(new_n568));
  XOR2_X1   g367(.A(G176gat), .B(G204gat), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NOR3_X1   g369(.A1(new_n564), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT98), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n570), .B1(new_n564), .B2(new_n566), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n574), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n521), .A2(KEYINPUT21), .ZN(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n498), .B1(KEYINPUT21), .B2(new_n521), .ZN(new_n581));
  XOR2_X1   g380(.A(new_n580), .B(new_n581), .Z(new_n582));
  XNOR2_X1  g381(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT89), .ZN(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT88), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n582), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n490), .A2(new_n558), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n546), .A2(new_n550), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n489), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n591), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT41), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n598), .B(KEYINPUT90), .Z(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G134gat), .B(G162gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n605));
  INV_X1    g404(.A(new_n603), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n591), .A2(new_n606), .A3(new_n593), .A4(new_n594), .ZN(new_n607));
  AND3_X1   g406(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n605), .B1(new_n604), .B2(new_n607), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n577), .A2(new_n590), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT99), .Z(new_n612));
  NAND4_X1  g411(.A1(new_n469), .A2(new_n471), .A3(new_n512), .A4(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT100), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(new_n417), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g415(.A1(new_n614), .A2(new_n422), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT101), .B1(new_n617), .B2(new_n495), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  OAI211_X1 g418(.A(new_n619), .B(G8gat), .C1(new_n614), .C2(new_n422), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT42), .ZN(new_n621));
  XOR2_X1   g420(.A(KEYINPUT16), .B(G8gat), .Z(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n617), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NOR4_X1   g423(.A1(new_n614), .A2(KEYINPUT42), .A3(new_n422), .A4(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n618), .B(new_n620), .C1(new_n623), .C2(new_n625), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n438), .A2(KEYINPUT73), .ZN(new_n628));
  INV_X1    g427(.A(new_n441), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n435), .B1(new_n309), .B2(KEYINPUT36), .ZN(new_n630));
  AOI211_X1 g429(.A(KEYINPUT72), .B(new_n437), .C1(new_n297), .C2(new_n308), .ZN(new_n631));
  OAI22_X1  g430(.A1(new_n628), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT103), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n614), .A2(new_n627), .A3(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n309), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n627), .B1(new_n614), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(KEYINPUT102), .B(new_n627), .C1(new_n614), .C2(new_n636), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(G1326gat));
  NOR2_X1   g440(.A1(new_n614), .A2(new_n355), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  INV_X1    g443(.A(KEYINPUT44), .ZN(new_n645));
  INV_X1    g444(.A(new_n430), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n647), .B1(new_n442), .B2(new_n467), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n383), .A2(new_n419), .ZN(new_n649));
  INV_X1    g448(.A(new_n453), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n466), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n651), .A2(new_n652), .B1(new_n420), .B2(new_n423), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n632), .A2(KEYINPUT105), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n646), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n645), .B1(new_n655), .B2(new_n610), .ZN(new_n656));
  INV_X1    g455(.A(new_n610), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n469), .A2(KEYINPUT44), .A3(new_n471), .A4(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n577), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n506), .B(new_n511), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n660), .A2(new_n661), .A3(new_n590), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(G29gat), .B1(new_n663), .B2(new_n417), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n660), .A2(new_n590), .A3(new_n610), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n469), .A2(new_n471), .A3(new_n512), .A4(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n416), .A2(new_n478), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OR3_X1    g468(.A1(new_n667), .A2(new_n665), .A3(new_n668), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(G1328gat));
  OAI21_X1  g470(.A(new_n483), .B1(new_n663), .B2(new_n422), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n422), .A2(new_n483), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT46), .B1(new_n667), .B2(new_n673), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n667), .A2(KEYINPUT46), .A3(new_n673), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(G1329gat));
  OAI21_X1  g475(.A(G43gat), .B1(new_n663), .B2(new_n632), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n636), .A2(G43gat), .ZN(new_n679));
  OR3_X1    g478(.A1(new_n667), .A2(KEYINPUT106), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(KEYINPUT106), .B1(new_n667), .B2(new_n679), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n678), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n659), .A2(new_n633), .A3(new_n662), .ZN(new_n684));
  AOI22_X1  g483(.A1(new_n684), .A2(G43gat), .B1(new_n681), .B2(new_n680), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n685), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g485(.A1(new_n667), .A2(G50gat), .A3(new_n355), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n656), .A2(new_n658), .A3(new_n423), .A4(new_n662), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n688), .B2(G50gat), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT48), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n689), .A2(KEYINPUT107), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(KEYINPUT107), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n690), .A2(KEYINPUT107), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n689), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n691), .A2(new_n694), .ZN(G1331gat));
  INV_X1    g494(.A(new_n590), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n512), .A2(new_n696), .A3(new_n657), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n660), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT108), .Z(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n655), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n416), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G57gat), .ZN(G1332gat));
  INV_X1    g501(.A(KEYINPUT49), .ZN(new_n703));
  INV_X1    g502(.A(G64gat), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n700), .B(new_n649), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1333gat));
  NAND2_X1  g506(.A1(new_n700), .A2(new_n633), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n636), .A2(G71gat), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n708), .A2(G71gat), .B1(new_n700), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g510(.A1(new_n700), .A2(new_n423), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT109), .B(G78gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1335gat));
  NOR3_X1   g513(.A1(new_n512), .A2(new_n590), .A3(new_n577), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n659), .A2(new_n416), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(G85gat), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n512), .A2(new_n590), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n648), .A2(new_n654), .ZN(new_n719));
  OAI211_X1 g518(.A(new_n657), .B(new_n718), .C1(new_n719), .C2(new_n646), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT51), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n655), .A2(new_n610), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(KEYINPUT51), .A3(new_n718), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n660), .A2(new_n537), .A3(new_n416), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT110), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n717), .B1(new_n726), .B2(new_n728), .ZN(G1336gat));
  NOR2_X1   g528(.A1(new_n422), .A2(new_n577), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n725), .A2(new_n538), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n656), .A2(new_n658), .A3(new_n649), .A4(new_n715), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G92gat), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n733), .B2(KEYINPUT111), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n731), .B(new_n733), .C1(KEYINPUT111), .C2(new_n735), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1337gat));
  NOR3_X1   g538(.A1(new_n636), .A2(G99gat), .A3(new_n577), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n656), .A2(new_n658), .A3(new_n633), .A4(new_n715), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G99gat), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT112), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n741), .A2(new_n746), .A3(new_n743), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1338gat));
  NOR3_X1   g547(.A1(new_n577), .A2(G106gat), .A3(new_n355), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT53), .B1(new_n725), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n656), .A2(new_n658), .A3(new_n423), .A4(new_n715), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT116), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT113), .B(G106gat), .Z(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(KEYINPUT116), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n751), .A2(KEYINPUT114), .A3(new_n753), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT114), .B1(new_n751), .B2(new_n753), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n749), .B(KEYINPUT115), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n722), .B2(new_n724), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n756), .B1(new_n761), .B2(new_n762), .ZN(G1339gat));
  NAND2_X1  g562(.A1(new_n556), .A2(new_n552), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n521), .B1(new_n555), .B2(new_n549), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n559), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n561), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n562), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n768), .A2(new_n515), .A3(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(KEYINPUT54), .A3(new_n563), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT54), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n772), .B(new_n516), .C1(new_n560), .C2(new_n562), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n773), .A2(KEYINPUT117), .A3(new_n570), .ZN(new_n774));
  AOI21_X1  g573(.A(KEYINPUT117), .B1(new_n773), .B2(new_n570), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n571), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n770), .A2(KEYINPUT54), .A3(new_n563), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n773), .A2(new_n570), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n773), .A2(KEYINPUT117), .A3(new_n570), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n779), .B1(new_n785), .B2(KEYINPUT55), .ZN(new_n786));
  OAI211_X1 g585(.A(KEYINPUT55), .B(new_n771), .C1(new_n774), .C2(new_n775), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(KEYINPUT118), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n778), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT119), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT119), .B(new_n778), .C1(new_n786), .C2(new_n788), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n791), .A2(new_n512), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n509), .A2(new_n500), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n502), .A2(new_n503), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g595(.A1(new_n511), .A2(new_n477), .B1(new_n796), .B2(new_n475), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(new_n575), .A3(new_n576), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n657), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n657), .A2(new_n797), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n791), .A2(new_n800), .A3(new_n792), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n696), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n697), .A2(new_n577), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n423), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n422), .A2(new_n416), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n636), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(G113gat), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n807), .A2(new_n808), .A3(new_n661), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n417), .B1(new_n802), .B2(new_n803), .ZN(new_n810));
  AND3_X1   g609(.A1(new_n810), .A2(new_n422), .A3(new_n424), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n512), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n812), .B2(new_n808), .ZN(G1340gat));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n660), .ZN(new_n814));
  INV_X1    g613(.A(G120gat), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g615(.A1(new_n804), .A2(G120gat), .A3(new_n660), .A4(new_n806), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT120), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n816), .A2(new_n820), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(G1341gat));
  INV_X1    g621(.A(G127gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n811), .A2(new_n823), .A3(new_n590), .ZN(new_n824));
  OAI21_X1  g623(.A(G127gat), .B1(new_n807), .B2(new_n696), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1342gat));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n804), .A2(new_n657), .A3(new_n806), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n828), .A2(new_n829), .A3(G134gat), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(G134gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(G134gat), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n649), .A2(new_n610), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n810), .A2(new_n833), .A3(new_n424), .A4(new_n834), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT56), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n827), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n835), .B(new_n838), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(KEYINPUT122), .C1(new_n831), .C2(new_n830), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n442), .A2(new_n805), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n802), .A2(new_n803), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n843), .B2(new_n423), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n798), .B1(new_n661), .B2(new_n789), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n610), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n696), .B1(new_n848), .B2(new_n801), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n845), .B(new_n355), .C1(new_n849), .C2(new_n803), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n842), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n661), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n633), .A2(new_n355), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n810), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n854), .A2(new_n649), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n327), .A3(new_n512), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT58), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n852), .A2(new_n859), .A3(new_n856), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n842), .A2(new_n660), .ZN(new_n862));
  INV_X1    g661(.A(new_n789), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n800), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n590), .B1(new_n865), .B2(KEYINPUT124), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n846), .A2(new_n610), .B1(new_n800), .B2(new_n863), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT124), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n866), .A2(new_n869), .B1(new_n661), .B2(new_n612), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n845), .B1(new_n870), .B2(new_n355), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n355), .A2(new_n845), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n843), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n862), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT59), .B1(new_n874), .B2(new_n329), .ZN(new_n875));
  OAI211_X1 g674(.A(new_n660), .B(new_n842), .C1(new_n844), .C2(new_n850), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n340), .A2(KEYINPUT59), .ZN(new_n878));
  AND3_X1   g677(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n877), .B1(new_n876), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n855), .A2(new_n340), .A3(new_n660), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1345gat));
  OAI21_X1  g682(.A(G155gat), .B1(new_n851), .B2(new_n696), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n855), .A2(new_n319), .A3(new_n590), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1346gat));
  OAI21_X1  g685(.A(G162gat), .B1(new_n851), .B2(new_n610), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n834), .A2(new_n320), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n854), .B2(new_n888), .ZN(G1347gat));
  NAND2_X1  g688(.A1(new_n649), .A2(new_n417), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n636), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n804), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(G169gat), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n661), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n416), .B1(new_n802), .B2(new_n803), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(new_n424), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n422), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n512), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n894), .B1(new_n898), .B2(new_n893), .ZN(G1348gat));
  OAI21_X1  g698(.A(G176gat), .B1(new_n892), .B2(new_n577), .ZN(new_n900));
  INV_X1    g699(.A(new_n730), .ZN(new_n901));
  OR2_X1    g700(.A1(new_n901), .A2(G176gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n900), .B1(new_n896), .B2(new_n902), .ZN(G1349gat));
  NAND3_X1  g702(.A1(new_n897), .A2(new_n246), .A3(new_n590), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n892), .B2(new_n696), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n908), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1350gat));
  NAND3_X1  g709(.A1(new_n897), .A2(new_n219), .A3(new_n657), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n912));
  INV_X1    g711(.A(new_n892), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n657), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n914), .B2(G190gat), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT61), .B(new_n219), .C1(new_n913), .C2(new_n657), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(G1351gat));
  NAND3_X1  g716(.A1(new_n895), .A2(new_n853), .A3(new_n649), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n512), .ZN(new_n921));
  INV_X1    g720(.A(G197gat), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n871), .A2(new_n873), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n633), .A2(new_n890), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n661), .A2(new_n922), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n921), .A2(new_n922), .B1(new_n926), .B2(new_n927), .ZN(G1352gat));
  OAI21_X1  g727(.A(G204gat), .B1(new_n925), .B2(new_n577), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n895), .A2(new_n853), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(G204gat), .A3(new_n901), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(G1353gat));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n312), .A3(new_n590), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n866), .A2(new_n869), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n612), .A2(new_n661), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n939), .B2(new_n423), .ZN(new_n940));
  INV_X1    g739(.A(new_n873), .ZN(new_n941));
  OAI211_X1 g740(.A(new_n590), .B(new_n924), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n942), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT63), .B1(new_n942), .B2(G211gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n936), .B1(new_n943), .B2(new_n944), .ZN(G1354gat));
  NAND2_X1  g744(.A1(new_n920), .A2(new_n657), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n657), .A2(G218gat), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT126), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n946), .A2(new_n313), .B1(new_n926), .B2(new_n948), .ZN(G1355gat));
endmodule


